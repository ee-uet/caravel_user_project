magic
tech sky130A
magscale 1 2
timestamp 1624055108
<< obsli1 >>
rect 489 493 578835 700791
<< obsm1 >>
rect 435 428 583450 702840
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 478 703464 8030 703520
rect 8254 703464 24222 703520
rect 24446 703464 40414 703520
rect 40638 703464 56698 703520
rect 56922 703464 72890 703520
rect 73114 703464 89082 703520
rect 89306 703464 105366 703520
rect 105590 703464 121558 703520
rect 121782 703464 137750 703520
rect 137974 703464 154034 703520
rect 154258 703464 170226 703520
rect 170450 703464 186418 703520
rect 186642 703464 202702 703520
rect 202926 703464 218894 703520
rect 219118 703464 235086 703520
rect 235310 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 300038 703520
rect 300262 703464 316230 703520
rect 316454 703464 332422 703520
rect 332646 703464 348706 703520
rect 348930 703464 364898 703520
rect 365122 703464 381090 703520
rect 381314 703464 397374 703520
rect 397598 703464 413566 703520
rect 413790 703464 429758 703520
rect 429982 703464 446042 703520
rect 446266 703464 462234 703520
rect 462458 703464 478426 703520
rect 478650 703464 494710 703520
rect 494934 703464 510902 703520
rect 511126 703464 527094 703520
rect 527318 703464 543378 703520
rect 543602 703464 559570 703520
rect 559794 703464 575762 703520
rect 575986 703464 583444 703520
rect 478 536 583444 703464
rect 478 478 486 536
rect 710 478 1590 536
rect 1814 478 2786 536
rect 3010 478 3982 536
rect 4206 478 5178 536
rect 5402 478 6374 536
rect 6598 478 7570 536
rect 7794 478 8674 536
rect 8898 478 9870 536
rect 10094 478 11066 536
rect 11290 478 12262 536
rect 12486 478 13458 536
rect 13682 478 14654 536
rect 14878 478 15850 536
rect 16074 478 16954 536
rect 17178 478 18150 536
rect 18374 478 19346 536
rect 19570 478 20542 536
rect 20766 478 21738 536
rect 21962 478 22934 536
rect 23158 478 24130 536
rect 24354 478 25234 536
rect 25458 478 26430 536
rect 26654 478 27626 536
rect 27850 478 28822 536
rect 29046 478 30018 536
rect 30242 478 31214 536
rect 31438 478 32318 536
rect 32542 478 33514 536
rect 33738 478 34710 536
rect 34934 478 35906 536
rect 36130 478 37102 536
rect 37326 478 38298 536
rect 38522 478 39494 536
rect 39718 478 40598 536
rect 40822 478 41794 536
rect 42018 478 42990 536
rect 43214 478 44186 536
rect 44410 478 45382 536
rect 45606 478 46578 536
rect 46802 478 47774 536
rect 47998 478 48878 536
rect 49102 478 50074 536
rect 50298 478 51270 536
rect 51494 478 52466 536
rect 52690 478 53662 536
rect 53886 478 54858 536
rect 55082 478 55962 536
rect 56186 478 57158 536
rect 57382 478 58354 536
rect 58578 478 59550 536
rect 59774 478 60746 536
rect 60970 478 61942 536
rect 62166 478 63138 536
rect 63362 478 64242 536
rect 64466 478 65438 536
rect 65662 478 66634 536
rect 66858 478 67830 536
rect 68054 478 69026 536
rect 69250 478 70222 536
rect 70446 478 71418 536
rect 71642 478 72522 536
rect 72746 478 73718 536
rect 73942 478 74914 536
rect 75138 478 76110 536
rect 76334 478 77306 536
rect 77530 478 78502 536
rect 78726 478 79606 536
rect 79830 478 80802 536
rect 81026 478 81998 536
rect 82222 478 83194 536
rect 83418 478 84390 536
rect 84614 478 85586 536
rect 85810 478 86782 536
rect 87006 478 87886 536
rect 88110 478 89082 536
rect 89306 478 90278 536
rect 90502 478 91474 536
rect 91698 478 92670 536
rect 92894 478 93866 536
rect 94090 478 95062 536
rect 95286 478 96166 536
rect 96390 478 97362 536
rect 97586 478 98558 536
rect 98782 478 99754 536
rect 99978 478 100950 536
rect 101174 478 102146 536
rect 102370 478 103250 536
rect 103474 478 104446 536
rect 104670 478 105642 536
rect 105866 478 106838 536
rect 107062 478 108034 536
rect 108258 478 109230 536
rect 109454 478 110426 536
rect 110650 478 111530 536
rect 111754 478 112726 536
rect 112950 478 113922 536
rect 114146 478 115118 536
rect 115342 478 116314 536
rect 116538 478 117510 536
rect 117734 478 118706 536
rect 118930 478 119810 536
rect 120034 478 121006 536
rect 121230 478 122202 536
rect 122426 478 123398 536
rect 123622 478 124594 536
rect 124818 478 125790 536
rect 126014 478 126894 536
rect 127118 478 128090 536
rect 128314 478 129286 536
rect 129510 478 130482 536
rect 130706 478 131678 536
rect 131902 478 132874 536
rect 133098 478 134070 536
rect 134294 478 135174 536
rect 135398 478 136370 536
rect 136594 478 137566 536
rect 137790 478 138762 536
rect 138986 478 139958 536
rect 140182 478 141154 536
rect 141378 478 142350 536
rect 142574 478 143454 536
rect 143678 478 144650 536
rect 144874 478 145846 536
rect 146070 478 147042 536
rect 147266 478 148238 536
rect 148462 478 149434 536
rect 149658 478 150538 536
rect 150762 478 151734 536
rect 151958 478 152930 536
rect 153154 478 154126 536
rect 154350 478 155322 536
rect 155546 478 156518 536
rect 156742 478 157714 536
rect 157938 478 158818 536
rect 159042 478 160014 536
rect 160238 478 161210 536
rect 161434 478 162406 536
rect 162630 478 163602 536
rect 163826 478 164798 536
rect 165022 478 165994 536
rect 166218 478 167098 536
rect 167322 478 168294 536
rect 168518 478 169490 536
rect 169714 478 170686 536
rect 170910 478 171882 536
rect 172106 478 173078 536
rect 173302 478 174182 536
rect 174406 478 175378 536
rect 175602 478 176574 536
rect 176798 478 177770 536
rect 177994 478 178966 536
rect 179190 478 180162 536
rect 180386 478 181358 536
rect 181582 478 182462 536
rect 182686 478 183658 536
rect 183882 478 184854 536
rect 185078 478 186050 536
rect 186274 478 187246 536
rect 187470 478 188442 536
rect 188666 478 189638 536
rect 189862 478 190742 536
rect 190966 478 191938 536
rect 192162 478 193134 536
rect 193358 478 194330 536
rect 194554 478 195526 536
rect 195750 478 196722 536
rect 196946 478 197826 536
rect 198050 478 199022 536
rect 199246 478 200218 536
rect 200442 478 201414 536
rect 201638 478 202610 536
rect 202834 478 203806 536
rect 204030 478 205002 536
rect 205226 478 206106 536
rect 206330 478 207302 536
rect 207526 478 208498 536
rect 208722 478 209694 536
rect 209918 478 210890 536
rect 211114 478 212086 536
rect 212310 478 213282 536
rect 213506 478 214386 536
rect 214610 478 215582 536
rect 215806 478 216778 536
rect 217002 478 217974 536
rect 218198 478 219170 536
rect 219394 478 220366 536
rect 220590 478 221470 536
rect 221694 478 222666 536
rect 222890 478 223862 536
rect 224086 478 225058 536
rect 225282 478 226254 536
rect 226478 478 227450 536
rect 227674 478 228646 536
rect 228870 478 229750 536
rect 229974 478 230946 536
rect 231170 478 232142 536
rect 232366 478 233338 536
rect 233562 478 234534 536
rect 234758 478 235730 536
rect 235954 478 236926 536
rect 237150 478 238030 536
rect 238254 478 239226 536
rect 239450 478 240422 536
rect 240646 478 241618 536
rect 241842 478 242814 536
rect 243038 478 244010 536
rect 244234 478 245114 536
rect 245338 478 246310 536
rect 246534 478 247506 536
rect 247730 478 248702 536
rect 248926 478 249898 536
rect 250122 478 251094 536
rect 251318 478 252290 536
rect 252514 478 253394 536
rect 253618 478 254590 536
rect 254814 478 255786 536
rect 256010 478 256982 536
rect 257206 478 258178 536
rect 258402 478 259374 536
rect 259598 478 260570 536
rect 260794 478 261674 536
rect 261898 478 262870 536
rect 263094 478 264066 536
rect 264290 478 265262 536
rect 265486 478 266458 536
rect 266682 478 267654 536
rect 267878 478 268758 536
rect 268982 478 269954 536
rect 270178 478 271150 536
rect 271374 478 272346 536
rect 272570 478 273542 536
rect 273766 478 274738 536
rect 274962 478 275934 536
rect 276158 478 277038 536
rect 277262 478 278234 536
rect 278458 478 279430 536
rect 279654 478 280626 536
rect 280850 478 281822 536
rect 282046 478 283018 536
rect 283242 478 284214 536
rect 284438 478 285318 536
rect 285542 478 286514 536
rect 286738 478 287710 536
rect 287934 478 288906 536
rect 289130 478 290102 536
rect 290326 478 291298 536
rect 291522 478 292494 536
rect 292718 478 293598 536
rect 293822 478 294794 536
rect 295018 478 295990 536
rect 296214 478 297186 536
rect 297410 478 298382 536
rect 298606 478 299578 536
rect 299802 478 300682 536
rect 300906 478 301878 536
rect 302102 478 303074 536
rect 303298 478 304270 536
rect 304494 478 305466 536
rect 305690 478 306662 536
rect 306886 478 307858 536
rect 308082 478 308962 536
rect 309186 478 310158 536
rect 310382 478 311354 536
rect 311578 478 312550 536
rect 312774 478 313746 536
rect 313970 478 314942 536
rect 315166 478 316138 536
rect 316362 478 317242 536
rect 317466 478 318438 536
rect 318662 478 319634 536
rect 319858 478 320830 536
rect 321054 478 322026 536
rect 322250 478 323222 536
rect 323446 478 324326 536
rect 324550 478 325522 536
rect 325746 478 326718 536
rect 326942 478 327914 536
rect 328138 478 329110 536
rect 329334 478 330306 536
rect 330530 478 331502 536
rect 331726 478 332606 536
rect 332830 478 333802 536
rect 334026 478 334998 536
rect 335222 478 336194 536
rect 336418 478 337390 536
rect 337614 478 338586 536
rect 338810 478 339782 536
rect 340006 478 340886 536
rect 341110 478 342082 536
rect 342306 478 343278 536
rect 343502 478 344474 536
rect 344698 478 345670 536
rect 345894 478 346866 536
rect 347090 478 347970 536
rect 348194 478 349166 536
rect 349390 478 350362 536
rect 350586 478 351558 536
rect 351782 478 352754 536
rect 352978 478 353950 536
rect 354174 478 355146 536
rect 355370 478 356250 536
rect 356474 478 357446 536
rect 357670 478 358642 536
rect 358866 478 359838 536
rect 360062 478 361034 536
rect 361258 478 362230 536
rect 362454 478 363426 536
rect 363650 478 364530 536
rect 364754 478 365726 536
rect 365950 478 366922 536
rect 367146 478 368118 536
rect 368342 478 369314 536
rect 369538 478 370510 536
rect 370734 478 371614 536
rect 371838 478 372810 536
rect 373034 478 374006 536
rect 374230 478 375202 536
rect 375426 478 376398 536
rect 376622 478 377594 536
rect 377818 478 378790 536
rect 379014 478 379894 536
rect 380118 478 381090 536
rect 381314 478 382286 536
rect 382510 478 383482 536
rect 383706 478 384678 536
rect 384902 478 385874 536
rect 386098 478 387070 536
rect 387294 478 388174 536
rect 388398 478 389370 536
rect 389594 478 390566 536
rect 390790 478 391762 536
rect 391986 478 392958 536
rect 393182 478 394154 536
rect 394378 478 395258 536
rect 395482 478 396454 536
rect 396678 478 397650 536
rect 397874 478 398846 536
rect 399070 478 400042 536
rect 400266 478 401238 536
rect 401462 478 402434 536
rect 402658 478 403538 536
rect 403762 478 404734 536
rect 404958 478 405930 536
rect 406154 478 407126 536
rect 407350 478 408322 536
rect 408546 478 409518 536
rect 409742 478 410714 536
rect 410938 478 411818 536
rect 412042 478 413014 536
rect 413238 478 414210 536
rect 414434 478 415406 536
rect 415630 478 416602 536
rect 416826 478 417798 536
rect 418022 478 418902 536
rect 419126 478 420098 536
rect 420322 478 421294 536
rect 421518 478 422490 536
rect 422714 478 423686 536
rect 423910 478 424882 536
rect 425106 478 426078 536
rect 426302 478 427182 536
rect 427406 478 428378 536
rect 428602 478 429574 536
rect 429798 478 430770 536
rect 430994 478 431966 536
rect 432190 478 433162 536
rect 433386 478 434358 536
rect 434582 478 435462 536
rect 435686 478 436658 536
rect 436882 478 437854 536
rect 438078 478 439050 536
rect 439274 478 440246 536
rect 440470 478 441442 536
rect 441666 478 442546 536
rect 442770 478 443742 536
rect 443966 478 444938 536
rect 445162 478 446134 536
rect 446358 478 447330 536
rect 447554 478 448526 536
rect 448750 478 449722 536
rect 449946 478 450826 536
rect 451050 478 452022 536
rect 452246 478 453218 536
rect 453442 478 454414 536
rect 454638 478 455610 536
rect 455834 478 456806 536
rect 457030 478 458002 536
rect 458226 478 459106 536
rect 459330 478 460302 536
rect 460526 478 461498 536
rect 461722 478 462694 536
rect 462918 478 463890 536
rect 464114 478 465086 536
rect 465310 478 466190 536
rect 466414 478 467386 536
rect 467610 478 468582 536
rect 468806 478 469778 536
rect 470002 478 470974 536
rect 471198 478 472170 536
rect 472394 478 473366 536
rect 473590 478 474470 536
rect 474694 478 475666 536
rect 475890 478 476862 536
rect 477086 478 478058 536
rect 478282 478 479254 536
rect 479478 478 480450 536
rect 480674 478 481646 536
rect 481870 478 482750 536
rect 482974 478 483946 536
rect 484170 478 485142 536
rect 485366 478 486338 536
rect 486562 478 487534 536
rect 487758 478 488730 536
rect 488954 478 489834 536
rect 490058 478 491030 536
rect 491254 478 492226 536
rect 492450 478 493422 536
rect 493646 478 494618 536
rect 494842 478 495814 536
rect 496038 478 497010 536
rect 497234 478 498114 536
rect 498338 478 499310 536
rect 499534 478 500506 536
rect 500730 478 501702 536
rect 501926 478 502898 536
rect 503122 478 504094 536
rect 504318 478 505290 536
rect 505514 478 506394 536
rect 506618 478 507590 536
rect 507814 478 508786 536
rect 509010 478 509982 536
rect 510206 478 511178 536
rect 511402 478 512374 536
rect 512598 478 513478 536
rect 513702 478 514674 536
rect 514898 478 515870 536
rect 516094 478 517066 536
rect 517290 478 518262 536
rect 518486 478 519458 536
rect 519682 478 520654 536
rect 520878 478 521758 536
rect 521982 478 522954 536
rect 523178 478 524150 536
rect 524374 478 525346 536
rect 525570 478 526542 536
rect 526766 478 527738 536
rect 527962 478 528934 536
rect 529158 478 530038 536
rect 530262 478 531234 536
rect 531458 478 532430 536
rect 532654 478 533626 536
rect 533850 478 534822 536
rect 535046 478 536018 536
rect 536242 478 537122 536
rect 537346 478 538318 536
rect 538542 478 539514 536
rect 539738 478 540710 536
rect 540934 478 541906 536
rect 542130 478 543102 536
rect 543326 478 544298 536
rect 544522 478 545402 536
rect 545626 478 546598 536
rect 546822 478 547794 536
rect 548018 478 548990 536
rect 549214 478 550186 536
rect 550410 478 551382 536
rect 551606 478 552578 536
rect 552802 478 553682 536
rect 553906 478 554878 536
rect 555102 478 556074 536
rect 556298 478 557270 536
rect 557494 478 558466 536
rect 558690 478 559662 536
rect 559886 478 560766 536
rect 560990 478 561962 536
rect 562186 478 563158 536
rect 563382 478 564354 536
rect 564578 478 565550 536
rect 565774 478 566746 536
rect 566970 478 567942 536
rect 568166 478 569046 536
rect 569270 478 570242 536
rect 570466 478 571438 536
rect 571662 478 572634 536
rect 572858 478 573830 536
rect 574054 478 575026 536
rect 575250 478 576222 536
rect 576446 478 577326 536
rect 577550 478 578522 536
rect 578746 478 579718 536
rect 579942 478 580914 536
rect 581138 478 582110 536
rect 582334 478 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 473 697540 583520 701793
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 473 697004 583440 697140
rect 473 684484 583520 697004
rect 560 684084 583520 684484
rect 473 684076 583520 684084
rect 473 683676 583440 684076
rect 473 671428 583520 683676
rect 560 671028 583520 671428
rect 473 670884 583520 671028
rect 473 670484 583440 670884
rect 473 658372 583520 670484
rect 560 657972 583520 658372
rect 473 657556 583520 657972
rect 473 657156 583440 657556
rect 473 645316 583520 657156
rect 560 644916 583520 645316
rect 473 644228 583520 644916
rect 473 643828 583440 644228
rect 473 632260 583520 643828
rect 560 631860 583520 632260
rect 473 631036 583520 631860
rect 473 630636 583440 631036
rect 473 619340 583520 630636
rect 560 618940 583520 619340
rect 473 617708 583520 618940
rect 473 617308 583440 617708
rect 473 606284 583520 617308
rect 560 605884 583520 606284
rect 473 604380 583520 605884
rect 473 603980 583440 604380
rect 473 593228 583520 603980
rect 560 592828 583520 593228
rect 473 591188 583520 592828
rect 473 590788 583440 591188
rect 473 580172 583520 590788
rect 560 579772 583520 580172
rect 473 577860 583520 579772
rect 473 577460 583440 577860
rect 473 567116 583520 577460
rect 560 566716 583520 567116
rect 473 564532 583520 566716
rect 473 564132 583440 564532
rect 473 554060 583520 564132
rect 560 553660 583520 554060
rect 473 551340 583520 553660
rect 473 550940 583440 551340
rect 473 541004 583520 550940
rect 560 540604 583520 541004
rect 473 538012 583520 540604
rect 473 537612 583440 538012
rect 473 528084 583520 537612
rect 560 527684 583520 528084
rect 473 524684 583520 527684
rect 473 524284 583440 524684
rect 473 515028 583520 524284
rect 560 514628 583520 515028
rect 473 511492 583520 514628
rect 473 511092 583440 511492
rect 473 501972 583520 511092
rect 560 501572 583520 501972
rect 473 498164 583520 501572
rect 473 497764 583440 498164
rect 473 488916 583520 497764
rect 560 488516 583520 488916
rect 473 484836 583520 488516
rect 473 484436 583440 484836
rect 473 475860 583520 484436
rect 560 475460 583520 475860
rect 473 471644 583520 475460
rect 473 471244 583440 471644
rect 473 462804 583520 471244
rect 560 462404 583520 462804
rect 473 458316 583520 462404
rect 473 457916 583440 458316
rect 473 449748 583520 457916
rect 560 449348 583520 449748
rect 473 444988 583520 449348
rect 473 444588 583440 444988
rect 473 436828 583520 444588
rect 560 436428 583520 436828
rect 473 431796 583520 436428
rect 473 431396 583440 431796
rect 473 423772 583520 431396
rect 560 423372 583520 423772
rect 473 418468 583520 423372
rect 473 418068 583440 418468
rect 473 410716 583520 418068
rect 560 410316 583520 410716
rect 473 405140 583520 410316
rect 473 404740 583440 405140
rect 473 397660 583520 404740
rect 560 397260 583520 397660
rect 473 391948 583520 397260
rect 473 391548 583440 391948
rect 473 384604 583520 391548
rect 560 384204 583520 384604
rect 473 378620 583520 384204
rect 473 378220 583440 378620
rect 473 371548 583520 378220
rect 560 371148 583520 371548
rect 473 365292 583520 371148
rect 473 364892 583440 365292
rect 473 358628 583520 364892
rect 560 358228 583520 358628
rect 473 352100 583520 358228
rect 473 351700 583440 352100
rect 473 345572 583520 351700
rect 560 345172 583520 345572
rect 473 338772 583520 345172
rect 473 338372 583440 338772
rect 473 332516 583520 338372
rect 560 332116 583520 332516
rect 473 325444 583520 332116
rect 473 325044 583440 325444
rect 473 319460 583520 325044
rect 560 319060 583520 319460
rect 473 312252 583520 319060
rect 473 311852 583440 312252
rect 473 306404 583520 311852
rect 560 306004 583520 306404
rect 473 298924 583520 306004
rect 473 298524 583440 298924
rect 473 293348 583520 298524
rect 560 292948 583520 293348
rect 473 285596 583520 292948
rect 473 285196 583440 285596
rect 473 280292 583520 285196
rect 560 279892 583520 280292
rect 473 272404 583520 279892
rect 473 272004 583440 272404
rect 473 267372 583520 272004
rect 560 266972 583520 267372
rect 473 259076 583520 266972
rect 473 258676 583440 259076
rect 473 254316 583520 258676
rect 560 253916 583520 254316
rect 473 245748 583520 253916
rect 473 245348 583440 245748
rect 473 241260 583520 245348
rect 560 240860 583520 241260
rect 473 232556 583520 240860
rect 473 232156 583440 232556
rect 473 228204 583520 232156
rect 560 227804 583520 228204
rect 473 219228 583520 227804
rect 473 218828 583440 219228
rect 473 215148 583520 218828
rect 560 214748 583520 215148
rect 473 205900 583520 214748
rect 473 205500 583440 205900
rect 473 202092 583520 205500
rect 560 201692 583520 202092
rect 473 192708 583520 201692
rect 473 192308 583440 192708
rect 473 189036 583520 192308
rect 560 188636 583520 189036
rect 473 179380 583520 188636
rect 473 178980 583440 179380
rect 473 176116 583520 178980
rect 560 175716 583520 176116
rect 473 166052 583520 175716
rect 473 165652 583440 166052
rect 473 163060 583520 165652
rect 560 162660 583520 163060
rect 473 152860 583520 162660
rect 473 152460 583440 152860
rect 473 150004 583520 152460
rect 560 149604 583520 150004
rect 473 139532 583520 149604
rect 473 139132 583440 139532
rect 473 136948 583520 139132
rect 560 136548 583520 136948
rect 473 126204 583520 136548
rect 473 125804 583440 126204
rect 473 123892 583520 125804
rect 560 123492 583520 123892
rect 473 113012 583520 123492
rect 473 112612 583440 113012
rect 473 110836 583520 112612
rect 560 110436 583520 110836
rect 473 99684 583520 110436
rect 473 99284 583440 99684
rect 473 97780 583520 99284
rect 560 97380 583520 97780
rect 473 86356 583520 97380
rect 473 85956 583440 86356
rect 473 84860 583520 85956
rect 560 84460 583520 84860
rect 473 73164 583520 84460
rect 473 72764 583440 73164
rect 473 71804 583520 72764
rect 560 71404 583520 71804
rect 473 59836 583520 71404
rect 473 59436 583440 59836
rect 473 58748 583520 59436
rect 560 58348 583520 58748
rect 473 46508 583520 58348
rect 473 46108 583440 46508
rect 473 45692 583520 46108
rect 560 45292 583520 45692
rect 473 33316 583520 45292
rect 473 32916 583440 33316
rect 473 32636 583520 32916
rect 560 32236 583520 32636
rect 473 19988 583520 32236
rect 473 19588 583440 19988
rect 473 19580 583520 19588
rect 560 19180 583520 19580
rect 473 6796 583520 19180
rect 473 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 473 579 583520 6260
<< metal4 >>
rect -8576 -7504 -7976 711440
rect -7636 -6564 -7036 710500
rect -6696 -5624 -6096 709560
rect -5756 -4684 -5156 708620
rect -4816 -3744 -4216 707680
rect -3876 -2804 -3276 706740
rect -2936 -1864 -2336 705800
rect -1996 -924 -1396 704860
rect 1804 -1864 2404 705800
rect 5404 -3744 6004 707680
rect 9004 -5624 9604 709560
rect 12604 -7504 13204 711440
rect 19804 690352 20404 705800
rect 23404 690400 24004 707680
rect 27004 690400 27604 709560
rect 30604 690400 31204 711440
rect 37804 690352 38404 705800
rect 41404 690400 42004 707680
rect 45004 690400 45604 709560
rect 48604 690400 49204 711440
rect 55804 690352 56404 705800
rect 59404 690400 60004 707680
rect 63004 690400 63604 709560
rect 66604 690400 67204 711440
rect 73804 690352 74404 705800
rect 77404 690400 78004 707680
rect 19804 620992 20404 630448
rect 23404 621040 24004 630400
rect 27004 621040 27604 630400
rect 30604 621040 31204 630400
rect 37804 620992 38404 630448
rect 41404 621040 42004 630400
rect 45004 621040 45604 630400
rect 48604 621040 49204 630400
rect 55804 620992 56404 630448
rect 59404 621040 60004 630400
rect 63004 621040 63604 630400
rect 66604 621040 67204 630400
rect 73804 620992 74404 630448
rect 77404 621040 78004 630400
rect 19804 551632 20404 561088
rect 23404 551680 24004 561040
rect 27004 551680 27604 561040
rect 30604 551680 31204 561040
rect 37804 551632 38404 561088
rect 41404 551680 42004 561040
rect 45004 551680 45604 561040
rect 48604 551680 49204 561040
rect 55804 551632 56404 561088
rect 59404 551680 60004 561040
rect 63004 551680 63604 561040
rect 66604 551680 67204 561040
rect 73804 551632 74404 561088
rect 77404 551680 78004 561040
rect 19804 482272 20404 491728
rect 23404 482320 24004 491680
rect 27004 482320 27604 491680
rect 30604 482320 31204 491680
rect 37804 482272 38404 491728
rect 41404 482320 42004 491680
rect 45004 482320 45604 491680
rect 48604 482320 49204 491680
rect 55804 482272 56404 491728
rect 59404 482320 60004 491680
rect 63004 482320 63604 491680
rect 66604 482320 67204 491680
rect 73804 482272 74404 491728
rect 77404 482320 78004 491680
rect 19804 412912 20404 422368
rect 23404 412960 24004 422320
rect 27004 412960 27604 422320
rect 30604 412960 31204 422320
rect 37804 412912 38404 422368
rect 41404 412960 42004 422320
rect 45004 412960 45604 422320
rect 48604 412960 49204 422320
rect 55804 412912 56404 422368
rect 59404 412960 60004 422320
rect 63004 412960 63604 422320
rect 66604 412960 67204 422320
rect 73804 412912 74404 422368
rect 77404 412960 78004 422320
rect 19804 343552 20404 353008
rect 23404 343600 24004 352960
rect 27004 343600 27604 352960
rect 30604 343600 31204 352960
rect 37804 343552 38404 353008
rect 41404 343600 42004 352960
rect 45004 343600 45604 352960
rect 48604 343600 49204 352960
rect 55804 343552 56404 353008
rect 59404 343600 60004 352960
rect 63004 343600 63604 352960
rect 66604 343600 67204 352960
rect 73804 343552 74404 353008
rect 77404 343600 78004 352960
rect 19804 274192 20404 283648
rect 23404 274240 24004 283600
rect 27004 274240 27604 283600
rect 30604 274240 31204 283600
rect 37804 274192 38404 283648
rect 41404 274240 42004 283600
rect 45004 274240 45604 283600
rect 48604 274240 49204 283600
rect 55804 274192 56404 283648
rect 59404 274240 60004 283600
rect 63004 274240 63604 283600
rect 66604 274240 67204 283600
rect 73804 274192 74404 283648
rect 77404 274240 78004 283600
rect 19804 204832 20404 214288
rect 23404 204880 24004 214240
rect 27004 204880 27604 214240
rect 30604 204880 31204 214240
rect 37804 204832 38404 214288
rect 41404 204880 42004 214240
rect 45004 204880 45604 214240
rect 48604 204880 49204 214240
rect 55804 204832 56404 214288
rect 59404 204880 60004 214240
rect 63004 204880 63604 214240
rect 66604 204880 67204 214240
rect 73804 204832 74404 214288
rect 77404 204880 78004 214240
rect 19804 -1864 20404 144928
rect 23404 -3744 24004 144880
rect 27004 -5624 27604 144880
rect 30604 -7504 31204 144880
rect 37804 132152 38404 144928
rect 41404 132200 42004 144880
rect 45004 132200 45604 144880
rect 48604 132200 49204 144880
rect 55804 132152 56404 144928
rect 59404 132200 60004 144880
rect 63004 132200 63604 144880
rect 66604 132200 67204 144880
rect 73804 132152 74404 144928
rect 77404 132200 78004 144880
rect 37804 -1864 38404 8248
rect 41404 -3744 42004 8200
rect 45004 -5624 45604 8200
rect 48604 -7504 49204 8200
rect 55804 -1864 56404 8248
rect 59404 -3744 60004 8200
rect 63004 -5624 63604 8200
rect 66604 -7504 67204 8200
rect 73804 -1864 74404 8248
rect 77404 -3744 78004 8200
rect 81004 -5624 81604 709560
rect 84604 -7504 85204 711440
rect 91804 -1864 92404 705800
rect 95404 132200 96004 707680
rect 99004 690400 99604 709560
rect 102604 690400 103204 711440
rect 109804 690352 110404 705800
rect 113404 690400 114004 707680
rect 117004 690400 117604 709560
rect 120604 690400 121204 711440
rect 127804 690352 128404 705800
rect 131404 690400 132004 707680
rect 99004 621040 99604 630400
rect 102604 621040 103204 630400
rect 109804 620992 110404 630448
rect 113404 621040 114004 630400
rect 117004 621040 117604 630400
rect 120604 621040 121204 630400
rect 127804 620992 128404 630448
rect 131404 621040 132004 630400
rect 99004 551680 99604 561040
rect 102604 551680 103204 561040
rect 109804 551632 110404 561088
rect 113404 551680 114004 561040
rect 117004 551680 117604 561040
rect 120604 551680 121204 561040
rect 127804 551632 128404 561088
rect 131404 551680 132004 561040
rect 99004 482320 99604 491680
rect 102604 482320 103204 491680
rect 109804 482272 110404 491728
rect 113404 482320 114004 491680
rect 117004 482320 117604 491680
rect 120604 482320 121204 491680
rect 127804 482272 128404 491728
rect 131404 482320 132004 491680
rect 99004 412960 99604 422320
rect 102604 412960 103204 422320
rect 109804 412912 110404 422368
rect 113404 412960 114004 422320
rect 117004 412960 117604 422320
rect 120604 412960 121204 422320
rect 127804 412912 128404 422368
rect 131404 412960 132004 422320
rect 99004 343600 99604 352960
rect 102604 343600 103204 352960
rect 109804 343552 110404 353008
rect 113404 343600 114004 352960
rect 117004 343600 117604 352960
rect 120604 343600 121204 352960
rect 127804 343552 128404 353008
rect 131404 343600 132004 352960
rect 99004 274240 99604 283600
rect 102604 274240 103204 283600
rect 109804 274192 110404 283648
rect 113404 274240 114004 283600
rect 117004 274240 117604 283600
rect 120604 274240 121204 283600
rect 127804 274192 128404 283648
rect 131404 274240 132004 283600
rect 99004 204880 99604 214240
rect 102604 204880 103204 214240
rect 109804 204832 110404 214288
rect 113404 204880 114004 214240
rect 117004 204880 117604 214240
rect 120604 204880 121204 214240
rect 127804 204832 128404 214288
rect 131404 204880 132004 214240
rect 99004 132200 99604 144880
rect 102604 132200 103204 144880
rect 109804 132152 110404 144928
rect 113404 132200 114004 144880
rect 117004 132200 117604 144880
rect 120604 132200 121204 144880
rect 127804 132152 128404 144928
rect 131404 132200 132004 144880
rect 135004 132200 135604 709560
rect 138604 132200 139204 711440
rect 145804 690352 146404 705800
rect 149404 690400 150004 707680
rect 153004 690400 153604 709560
rect 156604 690400 157204 711440
rect 163804 690352 164404 705800
rect 167404 690400 168004 707680
rect 171004 690400 171604 709560
rect 174604 690400 175204 711440
rect 145804 620992 146404 630448
rect 149404 621040 150004 630400
rect 153004 621040 153604 630400
rect 156604 621040 157204 630400
rect 163804 620992 164404 630448
rect 167404 621040 168004 630400
rect 171004 621040 171604 630400
rect 174604 621040 175204 630400
rect 145804 551632 146404 561088
rect 149404 551680 150004 561040
rect 153004 551680 153604 561040
rect 156604 551680 157204 561040
rect 163804 551632 164404 561088
rect 167404 551680 168004 561040
rect 171004 551680 171604 561040
rect 174604 551680 175204 561040
rect 145804 482272 146404 491728
rect 149404 482320 150004 491680
rect 153004 482320 153604 491680
rect 156604 482320 157204 491680
rect 163804 482272 164404 491728
rect 167404 482320 168004 491680
rect 171004 482320 171604 491680
rect 174604 482320 175204 491680
rect 145804 412912 146404 422368
rect 149404 412960 150004 422320
rect 153004 412960 153604 422320
rect 156604 412960 157204 422320
rect 163804 412912 164404 422368
rect 167404 412960 168004 422320
rect 171004 412960 171604 422320
rect 174604 412960 175204 422320
rect 145804 343552 146404 353008
rect 149404 343600 150004 352960
rect 153004 343600 153604 352960
rect 156604 343600 157204 352960
rect 163804 343552 164404 353008
rect 167404 343600 168004 352960
rect 171004 343600 171604 352960
rect 174604 343600 175204 352960
rect 145804 274192 146404 283648
rect 149404 274240 150004 283600
rect 153004 274240 153604 283600
rect 156604 274240 157204 283600
rect 163804 274192 164404 283648
rect 167404 274240 168004 283600
rect 171004 274240 171604 283600
rect 174604 274240 175204 283600
rect 145804 204832 146404 214288
rect 149404 204880 150004 214240
rect 153004 204880 153604 214240
rect 156604 204880 157204 214240
rect 163804 204832 164404 214288
rect 167404 204880 168004 214240
rect 171004 204880 171604 214240
rect 174604 204880 175204 214240
rect 145804 132152 146404 144928
rect 149404 132200 150004 144880
rect 153004 132200 153604 144880
rect 156604 132200 157204 144880
rect 95404 -3744 96004 8200
rect 99004 -5624 99604 8200
rect 102604 -7504 103204 8200
rect 109804 -1864 110404 8248
rect 113404 -3744 114004 8200
rect 117004 -5624 117604 8200
rect 120604 -7504 121204 8200
rect 127804 -1864 128404 8248
rect 131404 -3744 132004 8200
rect 135004 -5624 135604 8200
rect 138604 -7504 139204 8200
rect 145804 -1864 146404 8248
rect 149404 -3744 150004 8200
rect 153004 -5624 153604 8200
rect 156604 -7504 157204 8200
rect 163804 -1864 164404 144928
rect 167404 132200 168004 144880
rect 171004 132200 171604 144880
rect 174604 132200 175204 144880
rect 181804 132152 182404 705800
rect 185404 690400 186004 707680
rect 189004 690400 189604 709560
rect 192604 690400 193204 711440
rect 199804 690352 200404 705800
rect 203404 690400 204004 707680
rect 207004 690400 207604 709560
rect 210604 690400 211204 711440
rect 217804 690352 218404 705800
rect 221404 690400 222004 707680
rect 185404 621040 186004 630400
rect 189004 621040 189604 630400
rect 192604 621040 193204 630400
rect 199804 620992 200404 630448
rect 203404 621040 204004 630400
rect 207004 621040 207604 630400
rect 210604 621040 211204 630400
rect 217804 620992 218404 630448
rect 221404 621040 222004 630400
rect 185404 551680 186004 561040
rect 189004 551680 189604 561040
rect 192604 551680 193204 561040
rect 199804 551632 200404 561088
rect 203404 551680 204004 561040
rect 207004 551680 207604 561040
rect 210604 551680 211204 561040
rect 217804 551632 218404 561088
rect 221404 551680 222004 561040
rect 185404 482320 186004 491680
rect 189004 482320 189604 491680
rect 192604 482320 193204 491680
rect 199804 482272 200404 491728
rect 203404 482320 204004 491680
rect 207004 482320 207604 491680
rect 210604 482320 211204 491680
rect 217804 482272 218404 491728
rect 221404 482320 222004 491680
rect 185404 412960 186004 422320
rect 189004 412960 189604 422320
rect 192604 412960 193204 422320
rect 199804 412912 200404 422368
rect 203404 412960 204004 422320
rect 207004 412960 207604 422320
rect 210604 412960 211204 422320
rect 217804 412912 218404 422368
rect 221404 412960 222004 422320
rect 185404 343600 186004 352960
rect 189004 343600 189604 352960
rect 192604 343600 193204 352960
rect 199804 343552 200404 353008
rect 203404 343600 204004 352960
rect 207004 343600 207604 352960
rect 210604 343600 211204 352960
rect 217804 343552 218404 353008
rect 221404 343600 222004 352960
rect 185404 274240 186004 283600
rect 189004 274240 189604 283600
rect 192604 274240 193204 283600
rect 199804 274192 200404 283648
rect 203404 274240 204004 283600
rect 207004 274240 207604 283600
rect 210604 274240 211204 283600
rect 217804 274192 218404 283648
rect 221404 274240 222004 283600
rect 185404 204880 186004 214240
rect 189004 204880 189604 214240
rect 192604 204880 193204 214240
rect 199804 204832 200404 214288
rect 203404 204880 204004 214240
rect 207004 204880 207604 214240
rect 210604 204880 211204 214240
rect 217804 204832 218404 214288
rect 221404 204880 222004 214240
rect 185404 132200 186004 144880
rect 189004 132200 189604 144880
rect 192604 132200 193204 144880
rect 199804 132152 200404 144928
rect 203404 132200 204004 144880
rect 207004 132200 207604 144880
rect 210604 132200 211204 144880
rect 217804 132152 218404 144928
rect 221404 132200 222004 144880
rect 225004 132200 225604 709560
rect 228604 690400 229204 711440
rect 235804 690352 236404 705800
rect 239404 690400 240004 707680
rect 243004 690400 243604 709560
rect 246604 690400 247204 711440
rect 253804 690352 254404 705800
rect 257404 690400 258004 707680
rect 261004 690400 261604 709560
rect 264604 690400 265204 711440
rect 228604 621040 229204 630400
rect 235804 620992 236404 630448
rect 239404 621040 240004 630400
rect 243004 621040 243604 630400
rect 246604 621040 247204 630400
rect 253804 620992 254404 630448
rect 257404 621040 258004 630400
rect 261004 621040 261604 630400
rect 264604 621040 265204 630400
rect 228604 551680 229204 561040
rect 235804 551632 236404 561088
rect 239404 551680 240004 561040
rect 243004 551680 243604 561040
rect 246604 551680 247204 561040
rect 253804 551632 254404 561088
rect 257404 551680 258004 561040
rect 261004 551680 261604 561040
rect 264604 551680 265204 561040
rect 228604 482320 229204 491680
rect 235804 482272 236404 491728
rect 239404 482320 240004 491680
rect 243004 482320 243604 491680
rect 246604 482320 247204 491680
rect 253804 482272 254404 491728
rect 257404 482320 258004 491680
rect 261004 482320 261604 491680
rect 264604 482320 265204 491680
rect 228604 412960 229204 422320
rect 235804 412912 236404 422368
rect 239404 412960 240004 422320
rect 243004 412960 243604 422320
rect 246604 412960 247204 422320
rect 253804 412912 254404 422368
rect 257404 412960 258004 422320
rect 261004 412960 261604 422320
rect 264604 412960 265204 422320
rect 228604 343600 229204 352960
rect 235804 343552 236404 353008
rect 239404 343600 240004 352960
rect 243004 343600 243604 352960
rect 246604 343600 247204 352960
rect 253804 343552 254404 353008
rect 257404 343600 258004 352960
rect 261004 343600 261604 352960
rect 264604 343600 265204 352960
rect 228604 274240 229204 283600
rect 235804 274192 236404 283648
rect 239404 274240 240004 283600
rect 243004 274240 243604 283600
rect 246604 274240 247204 283600
rect 253804 274192 254404 283648
rect 257404 274240 258004 283600
rect 261004 274240 261604 283600
rect 264604 274240 265204 283600
rect 228604 204880 229204 214240
rect 235804 204832 236404 214288
rect 239404 204880 240004 214240
rect 243004 204880 243604 214240
rect 246604 204880 247204 214240
rect 253804 204832 254404 214288
rect 257404 204880 258004 214240
rect 261004 204880 261604 214240
rect 264604 204880 265204 214240
rect 228604 132200 229204 144880
rect 167404 -3744 168004 8200
rect 171004 -5624 171604 8200
rect 174604 -7504 175204 8200
rect 181804 -1864 182404 8248
rect 185404 -3744 186004 8200
rect 189004 -5624 189604 8200
rect 192604 -7504 193204 8200
rect 199804 -1864 200404 8248
rect 203404 -3744 204004 8200
rect 207004 -5624 207604 8200
rect 210604 -7504 211204 8200
rect 217804 -1864 218404 8248
rect 221404 -3744 222004 8200
rect 225004 -5624 225604 8200
rect 228604 -7504 229204 8200
rect 235804 -1864 236404 144928
rect 239404 132200 240004 144880
rect 243004 132200 243604 144880
rect 246604 132200 247204 144880
rect 253804 132152 254404 144928
rect 257404 132200 258004 144880
rect 261004 132200 261604 144880
rect 264604 132200 265204 144880
rect 271804 132152 272404 705800
rect 275404 690400 276004 707680
rect 279004 690400 279604 709560
rect 282604 690400 283204 711440
rect 289804 690352 290404 705800
rect 293404 690400 294004 707680
rect 297004 690400 297604 709560
rect 300604 690400 301204 711440
rect 307804 690352 308404 705800
rect 275404 621040 276004 630400
rect 279004 621040 279604 630400
rect 282604 621040 283204 630400
rect 289804 620992 290404 630448
rect 293404 621040 294004 630400
rect 297004 621040 297604 630400
rect 300604 621040 301204 630400
rect 307804 620992 308404 630448
rect 275404 551680 276004 561040
rect 279004 551680 279604 561040
rect 282604 551680 283204 561040
rect 289804 551632 290404 561088
rect 293404 551680 294004 561040
rect 297004 551680 297604 561040
rect 300604 551680 301204 561040
rect 307804 551632 308404 561088
rect 275404 482320 276004 491680
rect 279004 482320 279604 491680
rect 282604 482320 283204 491680
rect 289804 482272 290404 491728
rect 293404 482320 294004 491680
rect 297004 482320 297604 491680
rect 300604 482320 301204 491680
rect 307804 482272 308404 491728
rect 275404 412960 276004 422320
rect 279004 412960 279604 422320
rect 282604 412960 283204 422320
rect 289804 412912 290404 422368
rect 293404 412960 294004 422320
rect 297004 412960 297604 422320
rect 300604 412960 301204 422320
rect 307804 412912 308404 422368
rect 275404 343600 276004 352960
rect 279004 343600 279604 352960
rect 282604 343600 283204 352960
rect 289804 343552 290404 353008
rect 293404 343600 294004 352960
rect 297004 343600 297604 352960
rect 300604 343600 301204 352960
rect 307804 343552 308404 353008
rect 275404 274240 276004 283600
rect 279004 274240 279604 283600
rect 282604 274240 283204 283600
rect 289804 274192 290404 283648
rect 293404 274240 294004 283600
rect 297004 274240 297604 283600
rect 300604 274240 301204 283600
rect 307804 274192 308404 283648
rect 275404 204880 276004 214240
rect 279004 204880 279604 214240
rect 282604 204880 283204 214240
rect 289804 204832 290404 214288
rect 293404 204880 294004 214240
rect 297004 204880 297604 214240
rect 300604 204880 301204 214240
rect 307804 204832 308404 214288
rect 275404 132200 276004 144880
rect 279004 132200 279604 144880
rect 282604 132200 283204 144880
rect 289804 132152 290404 144928
rect 293404 132200 294004 144880
rect 297004 132200 297604 144880
rect 300604 132200 301204 144880
rect 239404 -3744 240004 8200
rect 243004 -5624 243604 8200
rect 246604 -7504 247204 8200
rect 253804 -1864 254404 8248
rect 257404 -3744 258004 8200
rect 261004 -5624 261604 8200
rect 264604 -7504 265204 8200
rect 271804 -1864 272404 8248
rect 275404 -3744 276004 8200
rect 279004 -5624 279604 8200
rect 282604 -7504 283204 8200
rect 289804 -1864 290404 8248
rect 293404 -3744 294004 8200
rect 297004 -5624 297604 8200
rect 300604 -7504 301204 8200
rect 307804 -1864 308404 144928
rect 311404 132200 312004 707680
rect 315004 132200 315604 709560
rect 318604 690400 319204 711440
rect 325804 690352 326404 705800
rect 329404 690400 330004 707680
rect 333004 690400 333604 709560
rect 336604 690400 337204 711440
rect 343804 690352 344404 705800
rect 347404 690400 348004 707680
rect 351004 690400 351604 709560
rect 354604 690400 355204 711440
rect 361804 690352 362404 705800
rect 365404 690400 366004 707680
rect 369004 690400 369604 709560
rect 372604 690400 373204 711440
rect 379804 690352 380404 705800
rect 383404 690400 384004 707680
rect 387004 690400 387604 709560
rect 390604 690400 391204 711440
rect 397804 690352 398404 705800
rect 318604 621040 319204 630400
rect 325804 620992 326404 630448
rect 329404 621040 330004 630400
rect 333004 621040 333604 630400
rect 336604 621040 337204 630400
rect 343804 620992 344404 630448
rect 347404 621040 348004 630400
rect 351004 621040 351604 630400
rect 354604 621040 355204 630400
rect 361804 620992 362404 630448
rect 365404 621040 366004 630400
rect 369004 621040 369604 630400
rect 372604 621040 373204 630400
rect 379804 620992 380404 630448
rect 383404 621040 384004 630400
rect 387004 621040 387604 630400
rect 390604 621040 391204 630400
rect 397804 620992 398404 630448
rect 318604 551680 319204 561040
rect 325804 551632 326404 561088
rect 329404 551680 330004 561040
rect 333004 551680 333604 561040
rect 336604 551680 337204 561040
rect 343804 551632 344404 561088
rect 347404 551680 348004 561040
rect 351004 551680 351604 561040
rect 354604 551680 355204 561040
rect 361804 551632 362404 561088
rect 365404 551680 366004 561040
rect 369004 551680 369604 561040
rect 372604 551680 373204 561040
rect 379804 551632 380404 561088
rect 383404 551680 384004 561040
rect 387004 551680 387604 561040
rect 390604 551680 391204 561040
rect 397804 551632 398404 561088
rect 318604 482320 319204 491680
rect 325804 482272 326404 491728
rect 329404 482320 330004 491680
rect 333004 482320 333604 491680
rect 336604 482320 337204 491680
rect 343804 482272 344404 491728
rect 347404 482320 348004 491680
rect 351004 482320 351604 491680
rect 354604 482320 355204 491680
rect 361804 482272 362404 491728
rect 365404 482320 366004 491680
rect 369004 482320 369604 491680
rect 372604 482320 373204 491680
rect 379804 482272 380404 491728
rect 383404 482320 384004 491680
rect 387004 482320 387604 491680
rect 390604 482320 391204 491680
rect 397804 482272 398404 491728
rect 318604 412960 319204 422320
rect 325804 412912 326404 422368
rect 329404 412960 330004 422320
rect 333004 412960 333604 422320
rect 336604 412960 337204 422320
rect 343804 412912 344404 422368
rect 347404 412960 348004 422320
rect 351004 412960 351604 422320
rect 354604 412960 355204 422320
rect 361804 412912 362404 422368
rect 365404 412960 366004 422320
rect 369004 412960 369604 422320
rect 372604 412960 373204 422320
rect 379804 412912 380404 422368
rect 383404 412960 384004 422320
rect 387004 412960 387604 422320
rect 390604 412960 391204 422320
rect 397804 412912 398404 422368
rect 318604 343600 319204 352960
rect 325804 343552 326404 353008
rect 329404 343600 330004 352960
rect 333004 343600 333604 352960
rect 336604 343600 337204 352960
rect 343804 343552 344404 353008
rect 347404 343600 348004 352960
rect 351004 343600 351604 352960
rect 354604 343600 355204 352960
rect 361804 343552 362404 353008
rect 365404 343600 366004 352960
rect 369004 343600 369604 352960
rect 372604 343600 373204 352960
rect 379804 343552 380404 353008
rect 383404 343600 384004 352960
rect 387004 343600 387604 352960
rect 390604 343600 391204 352960
rect 397804 343552 398404 353008
rect 318604 274240 319204 283600
rect 325804 274192 326404 283648
rect 329404 274240 330004 283600
rect 333004 274240 333604 283600
rect 336604 274240 337204 283600
rect 343804 274192 344404 283648
rect 347404 274240 348004 283600
rect 351004 274240 351604 283600
rect 354604 274240 355204 283600
rect 361804 274192 362404 283648
rect 365404 274240 366004 283600
rect 369004 274240 369604 283600
rect 372604 274240 373204 283600
rect 379804 274192 380404 283648
rect 383404 274240 384004 283600
rect 387004 274240 387604 283600
rect 390604 274240 391204 283600
rect 397804 274192 398404 283648
rect 318604 204880 319204 214240
rect 325804 204832 326404 214288
rect 329404 204880 330004 214240
rect 333004 204880 333604 214240
rect 336604 204880 337204 214240
rect 343804 204832 344404 214288
rect 347404 204880 348004 214240
rect 351004 204880 351604 214240
rect 354604 204880 355204 214240
rect 361804 204832 362404 214288
rect 365404 204880 366004 214240
rect 369004 204880 369604 214240
rect 372604 204880 373204 214240
rect 379804 204832 380404 214288
rect 383404 204880 384004 214240
rect 387004 204880 387604 214240
rect 390604 204880 391204 214240
rect 397804 204832 398404 214288
rect 318604 132200 319204 144880
rect 325804 132152 326404 144928
rect 329404 132200 330004 144880
rect 333004 132200 333604 144880
rect 336604 132200 337204 144880
rect 343804 132152 344404 144928
rect 347404 132200 348004 144880
rect 351004 132200 351604 144880
rect 354604 132200 355204 144880
rect 361804 132152 362404 144928
rect 365404 132200 366004 144880
rect 369004 132200 369604 144880
rect 372604 132200 373204 144880
rect 311404 -3744 312004 8200
rect 315004 -5624 315604 8200
rect 318604 -7504 319204 8200
rect 325804 -1864 326404 8248
rect 329404 -3744 330004 8200
rect 333004 -5624 333604 8200
rect 336604 -7504 337204 8200
rect 343804 -1864 344404 8248
rect 347404 -3744 348004 8200
rect 351004 -5624 351604 8200
rect 354604 -7504 355204 8200
rect 361804 -1864 362404 8248
rect 365404 -3744 366004 8200
rect 369004 -5624 369604 8200
rect 372604 -7504 373204 8200
rect 379804 -1864 380404 144928
rect 383404 -3744 384004 144880
rect 387004 132200 387604 144880
rect 390604 132200 391204 144880
rect 397804 132152 398404 144928
rect 401404 132200 402004 707680
rect 405004 690400 405604 709560
rect 408604 690400 409204 711440
rect 415804 690352 416404 705800
rect 419404 690400 420004 707680
rect 423004 690400 423604 709560
rect 426604 690400 427204 711440
rect 433804 690352 434404 705800
rect 437404 690400 438004 707680
rect 441004 690400 441604 709560
rect 405004 621040 405604 630400
rect 408604 621040 409204 630400
rect 415804 620992 416404 630448
rect 419404 621040 420004 630400
rect 423004 621040 423604 630400
rect 426604 621040 427204 630400
rect 433804 620992 434404 630448
rect 437404 621040 438004 630400
rect 441004 621040 441604 630400
rect 405004 551680 405604 561040
rect 408604 551680 409204 561040
rect 415804 551632 416404 561088
rect 419404 551680 420004 561040
rect 423004 551680 423604 561040
rect 426604 551680 427204 561040
rect 433804 551632 434404 561088
rect 437404 551680 438004 561040
rect 441004 551680 441604 561040
rect 405004 482320 405604 491680
rect 408604 482320 409204 491680
rect 415804 482272 416404 491728
rect 419404 482320 420004 491680
rect 423004 482320 423604 491680
rect 426604 482320 427204 491680
rect 433804 482272 434404 491728
rect 437404 482320 438004 491680
rect 441004 482320 441604 491680
rect 405004 412960 405604 422320
rect 408604 412960 409204 422320
rect 415804 412912 416404 422368
rect 419404 412960 420004 422320
rect 423004 412960 423604 422320
rect 426604 412960 427204 422320
rect 433804 412912 434404 422368
rect 437404 412960 438004 422320
rect 441004 412960 441604 422320
rect 405004 343600 405604 352960
rect 408604 343600 409204 352960
rect 415804 343552 416404 353008
rect 419404 343600 420004 352960
rect 423004 343600 423604 352960
rect 426604 343600 427204 352960
rect 433804 343552 434404 353008
rect 437404 343600 438004 352960
rect 441004 343600 441604 352960
rect 405004 274240 405604 283600
rect 408604 274240 409204 283600
rect 415804 274192 416404 283648
rect 419404 274240 420004 283600
rect 423004 274240 423604 283600
rect 426604 274240 427204 283600
rect 433804 274192 434404 283648
rect 437404 274240 438004 283600
rect 441004 274240 441604 283600
rect 405004 204880 405604 214240
rect 408604 204880 409204 214240
rect 415804 204832 416404 214288
rect 419404 204880 420004 214240
rect 423004 204880 423604 214240
rect 426604 204880 427204 214240
rect 433804 204832 434404 214288
rect 437404 204880 438004 214240
rect 441004 204880 441604 214240
rect 405004 132200 405604 144880
rect 408604 132200 409204 144880
rect 415804 132152 416404 144928
rect 419404 132200 420004 144880
rect 423004 132200 423604 144880
rect 426604 132200 427204 144880
rect 433804 132152 434404 144928
rect 437404 132200 438004 144880
rect 441004 132200 441604 144880
rect 444604 132200 445204 711440
rect 451804 690352 452404 705800
rect 455404 690400 456004 707680
rect 459004 690400 459604 709560
rect 462604 690400 463204 711440
rect 469804 690352 470404 705800
rect 473404 690400 474004 707680
rect 477004 690400 477604 709560
rect 480604 690400 481204 711440
rect 451804 620992 452404 630448
rect 455404 621040 456004 630400
rect 459004 621040 459604 630400
rect 462604 621040 463204 630400
rect 469804 620992 470404 630448
rect 473404 621040 474004 630400
rect 477004 621040 477604 630400
rect 480604 621040 481204 630400
rect 451804 551632 452404 561088
rect 455404 551680 456004 561040
rect 459004 551680 459604 561040
rect 462604 551680 463204 561040
rect 469804 551632 470404 561088
rect 473404 551680 474004 561040
rect 477004 551680 477604 561040
rect 480604 551680 481204 561040
rect 451804 482272 452404 491728
rect 455404 482320 456004 491680
rect 459004 482320 459604 491680
rect 462604 482320 463204 491680
rect 469804 482272 470404 491728
rect 473404 482320 474004 491680
rect 477004 482320 477604 491680
rect 480604 482320 481204 491680
rect 451804 412912 452404 422368
rect 455404 412960 456004 422320
rect 459004 412960 459604 422320
rect 462604 412960 463204 422320
rect 469804 412912 470404 422368
rect 473404 412960 474004 422320
rect 477004 412960 477604 422320
rect 480604 412960 481204 422320
rect 451804 343552 452404 353008
rect 455404 343600 456004 352960
rect 459004 343600 459604 352960
rect 462604 343600 463204 352960
rect 469804 343552 470404 353008
rect 473404 343600 474004 352960
rect 477004 343600 477604 352960
rect 480604 343600 481204 352960
rect 451804 274192 452404 283648
rect 455404 274240 456004 283600
rect 459004 274240 459604 283600
rect 462604 274240 463204 283600
rect 469804 274192 470404 283648
rect 473404 274240 474004 283600
rect 477004 274240 477604 283600
rect 480604 274240 481204 283600
rect 451804 204832 452404 214288
rect 455404 204880 456004 214240
rect 459004 204880 459604 214240
rect 462604 204880 463204 214240
rect 469804 204832 470404 214288
rect 473404 204880 474004 214240
rect 477004 204880 477604 214240
rect 480604 204880 481204 214240
rect 451804 132152 452404 144928
rect 455404 132200 456004 144880
rect 459004 132200 459604 144880
rect 462604 132200 463204 144880
rect 469804 132152 470404 144928
rect 473404 132200 474004 144880
rect 477004 132200 477604 144880
rect 480604 132200 481204 144880
rect 487804 132152 488404 705800
rect 491404 132200 492004 707680
rect 495004 690400 495604 709560
rect 498604 690400 499204 711440
rect 505804 690352 506404 705800
rect 509404 690400 510004 707680
rect 513004 690400 513604 709560
rect 516604 690400 517204 711440
rect 523804 690352 524404 705800
rect 527404 690400 528004 707680
rect 531004 690400 531604 709560
rect 495004 621040 495604 630400
rect 498604 621040 499204 630400
rect 505804 620992 506404 630448
rect 509404 621040 510004 630400
rect 513004 621040 513604 630400
rect 516604 621040 517204 630400
rect 523804 620992 524404 630448
rect 527404 621040 528004 630400
rect 531004 621040 531604 630400
rect 495004 551680 495604 561040
rect 498604 551680 499204 561040
rect 505804 551632 506404 561088
rect 509404 551680 510004 561040
rect 513004 551680 513604 561040
rect 516604 551680 517204 561040
rect 523804 551632 524404 561088
rect 527404 551680 528004 561040
rect 531004 551680 531604 561040
rect 495004 482320 495604 491680
rect 498604 482320 499204 491680
rect 505804 482272 506404 491728
rect 509404 482320 510004 491680
rect 513004 482320 513604 491680
rect 516604 482320 517204 491680
rect 523804 482272 524404 491728
rect 527404 482320 528004 491680
rect 531004 482320 531604 491680
rect 495004 412960 495604 422320
rect 498604 412960 499204 422320
rect 505804 412912 506404 422368
rect 509404 412960 510004 422320
rect 513004 412960 513604 422320
rect 516604 412960 517204 422320
rect 523804 412912 524404 422368
rect 527404 412960 528004 422320
rect 531004 412960 531604 422320
rect 495004 343600 495604 352960
rect 498604 343600 499204 352960
rect 505804 343552 506404 353008
rect 509404 343600 510004 352960
rect 513004 343600 513604 352960
rect 516604 343600 517204 352960
rect 523804 343552 524404 353008
rect 527404 343600 528004 352960
rect 531004 343600 531604 352960
rect 495004 274240 495604 283600
rect 498604 274240 499204 283600
rect 505804 274192 506404 283648
rect 509404 274240 510004 283600
rect 513004 274240 513604 283600
rect 516604 274240 517204 283600
rect 523804 274192 524404 283648
rect 527404 274240 528004 283600
rect 531004 274240 531604 283600
rect 495004 204880 495604 214240
rect 498604 204880 499204 214240
rect 505804 204832 506404 214288
rect 509404 204880 510004 214240
rect 513004 204880 513604 214240
rect 516604 204880 517204 214240
rect 523804 204832 524404 214288
rect 527404 204880 528004 214240
rect 531004 204880 531604 214240
rect 495004 132200 495604 144880
rect 498604 132200 499204 144880
rect 505804 132152 506404 144928
rect 509404 132200 510004 144880
rect 513004 132200 513604 144880
rect 516604 132200 517204 144880
rect 523804 132152 524404 144928
rect 527404 132200 528004 144880
rect 531004 132200 531604 144880
rect 534604 132200 535204 711440
rect 541804 690352 542404 705800
rect 545404 690400 546004 707680
rect 549004 690400 549604 709560
rect 552604 690400 553204 711440
rect 559804 690352 560404 705800
rect 563404 690400 564004 707680
rect 567004 690400 567604 709560
rect 570604 690400 571204 711440
rect 541804 620992 542404 630448
rect 545404 621040 546004 630400
rect 549004 621040 549604 630400
rect 552604 621040 553204 630400
rect 559804 620992 560404 630448
rect 563404 621040 564004 630400
rect 567004 621040 567604 630400
rect 570604 621040 571204 630400
rect 541804 551632 542404 561088
rect 545404 551680 546004 561040
rect 549004 551680 549604 561040
rect 552604 551680 553204 561040
rect 559804 551632 560404 561088
rect 563404 551680 564004 561040
rect 567004 551680 567604 561040
rect 570604 551680 571204 561040
rect 541804 482272 542404 491728
rect 545404 482320 546004 491680
rect 549004 482320 549604 491680
rect 552604 482320 553204 491680
rect 559804 482272 560404 491728
rect 563404 482320 564004 491680
rect 567004 482320 567604 491680
rect 570604 482320 571204 491680
rect 541804 412912 542404 422368
rect 545404 412960 546004 422320
rect 549004 412960 549604 422320
rect 552604 412960 553204 422320
rect 559804 412912 560404 422368
rect 563404 412960 564004 422320
rect 567004 412960 567604 422320
rect 570604 412960 571204 422320
rect 541804 343552 542404 353008
rect 545404 343600 546004 352960
rect 549004 343600 549604 352960
rect 552604 343600 553204 352960
rect 559804 343552 560404 353008
rect 563404 343600 564004 352960
rect 567004 343600 567604 352960
rect 570604 343600 571204 352960
rect 541804 274192 542404 283648
rect 545404 274240 546004 283600
rect 549004 274240 549604 283600
rect 552604 274240 553204 283600
rect 559804 274192 560404 283648
rect 563404 274240 564004 283600
rect 567004 274240 567604 283600
rect 570604 274240 571204 283600
rect 541804 204832 542404 214288
rect 545404 204880 546004 214240
rect 549004 204880 549604 214240
rect 552604 204880 553204 214240
rect 559804 204832 560404 214288
rect 563404 204880 564004 214240
rect 567004 204880 567604 214240
rect 570604 204880 571204 214240
rect 541804 132152 542404 144928
rect 545404 132200 546004 144880
rect 549004 132200 549604 144880
rect 552604 132200 553204 144880
rect 559804 132152 560404 144928
rect 563404 132200 564004 144880
rect 567004 132200 567604 144880
rect 387004 -5624 387604 8200
rect 390604 -7504 391204 8200
rect 397804 -1864 398404 8248
rect 401404 -3744 402004 8200
rect 405004 -5624 405604 8200
rect 408604 -7504 409204 8200
rect 415804 -1864 416404 8248
rect 419404 -3744 420004 8200
rect 423004 -5624 423604 8200
rect 426604 -7504 427204 8200
rect 433804 -1864 434404 8248
rect 437404 -3744 438004 8200
rect 441004 -5624 441604 8200
rect 444604 -7504 445204 8200
rect 451804 -1864 452404 8248
rect 455404 -3744 456004 8200
rect 459004 -5624 459604 8200
rect 462604 -7504 463204 8200
rect 469804 -1864 470404 8248
rect 473404 -3744 474004 8200
rect 477004 -5624 477604 8200
rect 480604 -7504 481204 8200
rect 487804 -1864 488404 8248
rect 491404 -3744 492004 8200
rect 495004 -5624 495604 8200
rect 498604 -7504 499204 8200
rect 505804 -1864 506404 8248
rect 509404 -3744 510004 8200
rect 513004 -5624 513604 8200
rect 516604 -7504 517204 8200
rect 523804 -1864 524404 8248
rect 527404 -3744 528004 8200
rect 531004 -5624 531604 8200
rect 534604 -7504 535204 8200
rect 541804 -1864 542404 8248
rect 545404 -3744 546004 8200
rect 549004 -5624 549604 8200
rect 552604 -7504 553204 8200
rect 559804 -1864 560404 8248
rect 563404 -3744 564004 8200
rect 567004 -5624 567604 8200
rect 570604 -7504 571204 144880
rect 577804 -1864 578404 705800
rect 581404 -3744 582004 707680
rect 585320 -924 585920 704860
rect 586260 -1864 586860 705800
rect 587200 -2804 587800 706740
rect 588140 -3744 588740 707680
rect 589080 -4684 589680 708620
rect 590020 -5624 590620 709560
rect 590960 -6564 591560 710500
rect 591900 -7504 592500 711440
<< obsm4 >>
rect 611 579 1724 700501
rect 2484 579 5324 700501
rect 6084 579 8924 700501
rect 9684 579 12524 700501
rect 13284 690272 19724 700501
rect 20484 690320 23324 700501
rect 24084 690320 26924 700501
rect 27684 690320 30524 700501
rect 31284 690320 37724 700501
rect 20484 690272 37724 690320
rect 38484 690320 41324 700501
rect 42084 690320 44924 700501
rect 45684 690320 48524 700501
rect 49284 690320 55724 700501
rect 38484 690272 55724 690320
rect 56484 690320 59324 700501
rect 60084 690320 62924 700501
rect 63684 690320 66524 700501
rect 67284 690320 73724 700501
rect 56484 690272 73724 690320
rect 74484 690320 77324 700501
rect 78084 690320 80924 700501
rect 74484 690272 80924 690320
rect 13284 630528 80924 690272
rect 13284 620912 19724 630528
rect 20484 630480 37724 630528
rect 20484 620960 23324 630480
rect 24084 620960 26924 630480
rect 27684 620960 30524 630480
rect 31284 620960 37724 630480
rect 38484 630480 55724 630528
rect 20484 620912 37724 620960
rect 38484 620960 41324 630480
rect 42084 620960 44924 630480
rect 45684 620960 48524 630480
rect 49284 620960 55724 630480
rect 56484 630480 73724 630528
rect 38484 620912 55724 620960
rect 56484 620960 59324 630480
rect 60084 620960 62924 630480
rect 63684 620960 66524 630480
rect 67284 620960 73724 630480
rect 74484 630480 80924 630528
rect 56484 620912 73724 620960
rect 74484 620960 77324 630480
rect 78084 620960 80924 630480
rect 74484 620912 80924 620960
rect 13284 561168 80924 620912
rect 13284 551552 19724 561168
rect 20484 561120 37724 561168
rect 20484 551600 23324 561120
rect 24084 551600 26924 561120
rect 27684 551600 30524 561120
rect 31284 551600 37724 561120
rect 38484 561120 55724 561168
rect 20484 551552 37724 551600
rect 38484 551600 41324 561120
rect 42084 551600 44924 561120
rect 45684 551600 48524 561120
rect 49284 551600 55724 561120
rect 56484 561120 73724 561168
rect 38484 551552 55724 551600
rect 56484 551600 59324 561120
rect 60084 551600 62924 561120
rect 63684 551600 66524 561120
rect 67284 551600 73724 561120
rect 74484 561120 80924 561168
rect 56484 551552 73724 551600
rect 74484 551600 77324 561120
rect 78084 551600 80924 561120
rect 74484 551552 80924 551600
rect 13284 491808 80924 551552
rect 13284 482192 19724 491808
rect 20484 491760 37724 491808
rect 20484 482240 23324 491760
rect 24084 482240 26924 491760
rect 27684 482240 30524 491760
rect 31284 482240 37724 491760
rect 38484 491760 55724 491808
rect 20484 482192 37724 482240
rect 38484 482240 41324 491760
rect 42084 482240 44924 491760
rect 45684 482240 48524 491760
rect 49284 482240 55724 491760
rect 56484 491760 73724 491808
rect 38484 482192 55724 482240
rect 56484 482240 59324 491760
rect 60084 482240 62924 491760
rect 63684 482240 66524 491760
rect 67284 482240 73724 491760
rect 74484 491760 80924 491808
rect 56484 482192 73724 482240
rect 74484 482240 77324 491760
rect 78084 482240 80924 491760
rect 74484 482192 80924 482240
rect 13284 422448 80924 482192
rect 13284 412832 19724 422448
rect 20484 422400 37724 422448
rect 20484 412880 23324 422400
rect 24084 412880 26924 422400
rect 27684 412880 30524 422400
rect 31284 412880 37724 422400
rect 38484 422400 55724 422448
rect 20484 412832 37724 412880
rect 38484 412880 41324 422400
rect 42084 412880 44924 422400
rect 45684 412880 48524 422400
rect 49284 412880 55724 422400
rect 56484 422400 73724 422448
rect 38484 412832 55724 412880
rect 56484 412880 59324 422400
rect 60084 412880 62924 422400
rect 63684 412880 66524 422400
rect 67284 412880 73724 422400
rect 74484 422400 80924 422448
rect 56484 412832 73724 412880
rect 74484 412880 77324 422400
rect 78084 412880 80924 422400
rect 74484 412832 80924 412880
rect 13284 353088 80924 412832
rect 13284 343472 19724 353088
rect 20484 353040 37724 353088
rect 20484 343520 23324 353040
rect 24084 343520 26924 353040
rect 27684 343520 30524 353040
rect 31284 343520 37724 353040
rect 38484 353040 55724 353088
rect 20484 343472 37724 343520
rect 38484 343520 41324 353040
rect 42084 343520 44924 353040
rect 45684 343520 48524 353040
rect 49284 343520 55724 353040
rect 56484 353040 73724 353088
rect 38484 343472 55724 343520
rect 56484 343520 59324 353040
rect 60084 343520 62924 353040
rect 63684 343520 66524 353040
rect 67284 343520 73724 353040
rect 74484 353040 80924 353088
rect 56484 343472 73724 343520
rect 74484 343520 77324 353040
rect 78084 343520 80924 353040
rect 74484 343472 80924 343520
rect 13284 283728 80924 343472
rect 13284 274112 19724 283728
rect 20484 283680 37724 283728
rect 20484 274160 23324 283680
rect 24084 274160 26924 283680
rect 27684 274160 30524 283680
rect 31284 274160 37724 283680
rect 38484 283680 55724 283728
rect 20484 274112 37724 274160
rect 38484 274160 41324 283680
rect 42084 274160 44924 283680
rect 45684 274160 48524 283680
rect 49284 274160 55724 283680
rect 56484 283680 73724 283728
rect 38484 274112 55724 274160
rect 56484 274160 59324 283680
rect 60084 274160 62924 283680
rect 63684 274160 66524 283680
rect 67284 274160 73724 283680
rect 74484 283680 80924 283728
rect 56484 274112 73724 274160
rect 74484 274160 77324 283680
rect 78084 274160 80924 283680
rect 74484 274112 80924 274160
rect 13284 214368 80924 274112
rect 13284 204752 19724 214368
rect 20484 214320 37724 214368
rect 20484 204800 23324 214320
rect 24084 204800 26924 214320
rect 27684 204800 30524 214320
rect 31284 204800 37724 214320
rect 38484 214320 55724 214368
rect 20484 204752 37724 204800
rect 38484 204800 41324 214320
rect 42084 204800 44924 214320
rect 45684 204800 48524 214320
rect 49284 204800 55724 214320
rect 56484 214320 73724 214368
rect 38484 204752 55724 204800
rect 56484 204800 59324 214320
rect 60084 204800 62924 214320
rect 63684 204800 66524 214320
rect 67284 204800 73724 214320
rect 74484 214320 80924 214368
rect 56484 204752 73724 204800
rect 74484 204800 77324 214320
rect 78084 204800 80924 214320
rect 74484 204752 80924 204800
rect 13284 145008 80924 204752
rect 13284 579 19724 145008
rect 20484 144960 37724 145008
rect 20484 579 23324 144960
rect 24084 579 26924 144960
rect 27684 579 30524 144960
rect 31284 132072 37724 144960
rect 38484 144960 55724 145008
rect 38484 132120 41324 144960
rect 42084 132120 44924 144960
rect 45684 132120 48524 144960
rect 49284 132120 55724 144960
rect 56484 144960 73724 145008
rect 38484 132072 55724 132120
rect 56484 132120 59324 144960
rect 60084 132120 62924 144960
rect 63684 132120 66524 144960
rect 67284 132120 73724 144960
rect 74484 144960 80924 145008
rect 56484 132072 73724 132120
rect 74484 132120 77324 144960
rect 78084 132120 80924 144960
rect 74484 132072 80924 132120
rect 31284 8328 80924 132072
rect 31284 579 37724 8328
rect 38484 8280 55724 8328
rect 38484 579 41324 8280
rect 42084 579 44924 8280
rect 45684 579 48524 8280
rect 49284 579 55724 8280
rect 56484 8280 73724 8328
rect 56484 579 59324 8280
rect 60084 579 62924 8280
rect 63684 579 66524 8280
rect 67284 579 73724 8280
rect 74484 8280 80924 8328
rect 74484 579 77324 8280
rect 78084 579 80924 8280
rect 81684 579 84524 700501
rect 85284 579 91724 700501
rect 92484 132120 95324 700501
rect 96084 690320 98924 700501
rect 99684 690320 102524 700501
rect 103284 690320 109724 700501
rect 96084 690272 109724 690320
rect 110484 690320 113324 700501
rect 114084 690320 116924 700501
rect 117684 690320 120524 700501
rect 121284 690320 127724 700501
rect 110484 690272 127724 690320
rect 128484 690320 131324 700501
rect 132084 690320 134924 700501
rect 128484 690272 134924 690320
rect 96084 630528 134924 690272
rect 96084 630480 109724 630528
rect 96084 620960 98924 630480
rect 99684 620960 102524 630480
rect 103284 620960 109724 630480
rect 110484 630480 127724 630528
rect 96084 620912 109724 620960
rect 110484 620960 113324 630480
rect 114084 620960 116924 630480
rect 117684 620960 120524 630480
rect 121284 620960 127724 630480
rect 128484 630480 134924 630528
rect 110484 620912 127724 620960
rect 128484 620960 131324 630480
rect 132084 620960 134924 630480
rect 128484 620912 134924 620960
rect 96084 561168 134924 620912
rect 96084 561120 109724 561168
rect 96084 551600 98924 561120
rect 99684 551600 102524 561120
rect 103284 551600 109724 561120
rect 110484 561120 127724 561168
rect 96084 551552 109724 551600
rect 110484 551600 113324 561120
rect 114084 551600 116924 561120
rect 117684 551600 120524 561120
rect 121284 551600 127724 561120
rect 128484 561120 134924 561168
rect 110484 551552 127724 551600
rect 128484 551600 131324 561120
rect 132084 551600 134924 561120
rect 128484 551552 134924 551600
rect 96084 491808 134924 551552
rect 96084 491760 109724 491808
rect 96084 482240 98924 491760
rect 99684 482240 102524 491760
rect 103284 482240 109724 491760
rect 110484 491760 127724 491808
rect 96084 482192 109724 482240
rect 110484 482240 113324 491760
rect 114084 482240 116924 491760
rect 117684 482240 120524 491760
rect 121284 482240 127724 491760
rect 128484 491760 134924 491808
rect 110484 482192 127724 482240
rect 128484 482240 131324 491760
rect 132084 482240 134924 491760
rect 128484 482192 134924 482240
rect 96084 422448 134924 482192
rect 96084 422400 109724 422448
rect 96084 412880 98924 422400
rect 99684 412880 102524 422400
rect 103284 412880 109724 422400
rect 110484 422400 127724 422448
rect 96084 412832 109724 412880
rect 110484 412880 113324 422400
rect 114084 412880 116924 422400
rect 117684 412880 120524 422400
rect 121284 412880 127724 422400
rect 128484 422400 134924 422448
rect 110484 412832 127724 412880
rect 128484 412880 131324 422400
rect 132084 412880 134924 422400
rect 128484 412832 134924 412880
rect 96084 353088 134924 412832
rect 96084 353040 109724 353088
rect 96084 343520 98924 353040
rect 99684 343520 102524 353040
rect 103284 343520 109724 353040
rect 110484 353040 127724 353088
rect 96084 343472 109724 343520
rect 110484 343520 113324 353040
rect 114084 343520 116924 353040
rect 117684 343520 120524 353040
rect 121284 343520 127724 353040
rect 128484 353040 134924 353088
rect 110484 343472 127724 343520
rect 128484 343520 131324 353040
rect 132084 343520 134924 353040
rect 128484 343472 134924 343520
rect 96084 283728 134924 343472
rect 96084 283680 109724 283728
rect 96084 274160 98924 283680
rect 99684 274160 102524 283680
rect 103284 274160 109724 283680
rect 110484 283680 127724 283728
rect 96084 274112 109724 274160
rect 110484 274160 113324 283680
rect 114084 274160 116924 283680
rect 117684 274160 120524 283680
rect 121284 274160 127724 283680
rect 128484 283680 134924 283728
rect 110484 274112 127724 274160
rect 128484 274160 131324 283680
rect 132084 274160 134924 283680
rect 128484 274112 134924 274160
rect 96084 214368 134924 274112
rect 96084 214320 109724 214368
rect 96084 204800 98924 214320
rect 99684 204800 102524 214320
rect 103284 204800 109724 214320
rect 110484 214320 127724 214368
rect 96084 204752 109724 204800
rect 110484 204800 113324 214320
rect 114084 204800 116924 214320
rect 117684 204800 120524 214320
rect 121284 204800 127724 214320
rect 128484 214320 134924 214368
rect 110484 204752 127724 204800
rect 128484 204800 131324 214320
rect 132084 204800 134924 214320
rect 128484 204752 134924 204800
rect 96084 145008 134924 204752
rect 96084 144960 109724 145008
rect 96084 132120 98924 144960
rect 99684 132120 102524 144960
rect 103284 132120 109724 144960
rect 110484 144960 127724 145008
rect 92484 132072 109724 132120
rect 110484 132120 113324 144960
rect 114084 132120 116924 144960
rect 117684 132120 120524 144960
rect 121284 132120 127724 144960
rect 128484 144960 134924 145008
rect 110484 132072 127724 132120
rect 128484 132120 131324 144960
rect 132084 132120 134924 144960
rect 135684 132120 138524 700501
rect 139284 690272 145724 700501
rect 146484 690320 149324 700501
rect 150084 690320 152924 700501
rect 153684 690320 156524 700501
rect 157284 690320 163724 700501
rect 146484 690272 163724 690320
rect 164484 690320 167324 700501
rect 168084 690320 170924 700501
rect 171684 690320 174524 700501
rect 175284 690320 181724 700501
rect 164484 690272 181724 690320
rect 139284 630528 181724 690272
rect 139284 620912 145724 630528
rect 146484 630480 163724 630528
rect 146484 620960 149324 630480
rect 150084 620960 152924 630480
rect 153684 620960 156524 630480
rect 157284 620960 163724 630480
rect 164484 630480 181724 630528
rect 146484 620912 163724 620960
rect 164484 620960 167324 630480
rect 168084 620960 170924 630480
rect 171684 620960 174524 630480
rect 175284 620960 181724 630480
rect 164484 620912 181724 620960
rect 139284 561168 181724 620912
rect 139284 551552 145724 561168
rect 146484 561120 163724 561168
rect 146484 551600 149324 561120
rect 150084 551600 152924 561120
rect 153684 551600 156524 561120
rect 157284 551600 163724 561120
rect 164484 561120 181724 561168
rect 146484 551552 163724 551600
rect 164484 551600 167324 561120
rect 168084 551600 170924 561120
rect 171684 551600 174524 561120
rect 175284 551600 181724 561120
rect 164484 551552 181724 551600
rect 139284 491808 181724 551552
rect 139284 482192 145724 491808
rect 146484 491760 163724 491808
rect 146484 482240 149324 491760
rect 150084 482240 152924 491760
rect 153684 482240 156524 491760
rect 157284 482240 163724 491760
rect 164484 491760 181724 491808
rect 146484 482192 163724 482240
rect 164484 482240 167324 491760
rect 168084 482240 170924 491760
rect 171684 482240 174524 491760
rect 175284 482240 181724 491760
rect 164484 482192 181724 482240
rect 139284 422448 181724 482192
rect 139284 412832 145724 422448
rect 146484 422400 163724 422448
rect 146484 412880 149324 422400
rect 150084 412880 152924 422400
rect 153684 412880 156524 422400
rect 157284 412880 163724 422400
rect 164484 422400 181724 422448
rect 146484 412832 163724 412880
rect 164484 412880 167324 422400
rect 168084 412880 170924 422400
rect 171684 412880 174524 422400
rect 175284 412880 181724 422400
rect 164484 412832 181724 412880
rect 139284 353088 181724 412832
rect 139284 343472 145724 353088
rect 146484 353040 163724 353088
rect 146484 343520 149324 353040
rect 150084 343520 152924 353040
rect 153684 343520 156524 353040
rect 157284 343520 163724 353040
rect 164484 353040 181724 353088
rect 146484 343472 163724 343520
rect 164484 343520 167324 353040
rect 168084 343520 170924 353040
rect 171684 343520 174524 353040
rect 175284 343520 181724 353040
rect 164484 343472 181724 343520
rect 139284 283728 181724 343472
rect 139284 274112 145724 283728
rect 146484 283680 163724 283728
rect 146484 274160 149324 283680
rect 150084 274160 152924 283680
rect 153684 274160 156524 283680
rect 157284 274160 163724 283680
rect 164484 283680 181724 283728
rect 146484 274112 163724 274160
rect 164484 274160 167324 283680
rect 168084 274160 170924 283680
rect 171684 274160 174524 283680
rect 175284 274160 181724 283680
rect 164484 274112 181724 274160
rect 139284 214368 181724 274112
rect 139284 204752 145724 214368
rect 146484 214320 163724 214368
rect 146484 204800 149324 214320
rect 150084 204800 152924 214320
rect 153684 204800 156524 214320
rect 157284 204800 163724 214320
rect 164484 214320 181724 214368
rect 146484 204752 163724 204800
rect 164484 204800 167324 214320
rect 168084 204800 170924 214320
rect 171684 204800 174524 214320
rect 175284 204800 181724 214320
rect 164484 204752 181724 204800
rect 139284 145008 181724 204752
rect 139284 132120 145724 145008
rect 146484 144960 163724 145008
rect 128484 132072 145724 132120
rect 146484 132120 149324 144960
rect 150084 132120 152924 144960
rect 153684 132120 156524 144960
rect 157284 132120 163724 144960
rect 164484 144960 181724 145008
rect 146484 132072 163724 132120
rect 92484 8328 163724 132072
rect 92484 8280 109724 8328
rect 92484 579 95324 8280
rect 96084 579 98924 8280
rect 99684 579 102524 8280
rect 103284 579 109724 8280
rect 110484 8280 127724 8328
rect 110484 579 113324 8280
rect 114084 579 116924 8280
rect 117684 579 120524 8280
rect 121284 579 127724 8280
rect 128484 8280 145724 8328
rect 128484 579 131324 8280
rect 132084 579 134924 8280
rect 135684 579 138524 8280
rect 139284 579 145724 8280
rect 146484 8280 163724 8328
rect 146484 579 149324 8280
rect 150084 579 152924 8280
rect 153684 579 156524 8280
rect 157284 579 163724 8280
rect 164484 132120 167324 144960
rect 168084 132120 170924 144960
rect 171684 132120 174524 144960
rect 175284 132120 181724 144960
rect 182484 690320 185324 700501
rect 186084 690320 188924 700501
rect 189684 690320 192524 700501
rect 193284 690320 199724 700501
rect 182484 690272 199724 690320
rect 200484 690320 203324 700501
rect 204084 690320 206924 700501
rect 207684 690320 210524 700501
rect 211284 690320 217724 700501
rect 200484 690272 217724 690320
rect 218484 690320 221324 700501
rect 222084 690320 224924 700501
rect 218484 690272 224924 690320
rect 182484 630528 224924 690272
rect 182484 630480 199724 630528
rect 182484 620960 185324 630480
rect 186084 620960 188924 630480
rect 189684 620960 192524 630480
rect 193284 620960 199724 630480
rect 200484 630480 217724 630528
rect 182484 620912 199724 620960
rect 200484 620960 203324 630480
rect 204084 620960 206924 630480
rect 207684 620960 210524 630480
rect 211284 620960 217724 630480
rect 218484 630480 224924 630528
rect 200484 620912 217724 620960
rect 218484 620960 221324 630480
rect 222084 620960 224924 630480
rect 218484 620912 224924 620960
rect 182484 561168 224924 620912
rect 182484 561120 199724 561168
rect 182484 551600 185324 561120
rect 186084 551600 188924 561120
rect 189684 551600 192524 561120
rect 193284 551600 199724 561120
rect 200484 561120 217724 561168
rect 182484 551552 199724 551600
rect 200484 551600 203324 561120
rect 204084 551600 206924 561120
rect 207684 551600 210524 561120
rect 211284 551600 217724 561120
rect 218484 561120 224924 561168
rect 200484 551552 217724 551600
rect 218484 551600 221324 561120
rect 222084 551600 224924 561120
rect 218484 551552 224924 551600
rect 182484 491808 224924 551552
rect 182484 491760 199724 491808
rect 182484 482240 185324 491760
rect 186084 482240 188924 491760
rect 189684 482240 192524 491760
rect 193284 482240 199724 491760
rect 200484 491760 217724 491808
rect 182484 482192 199724 482240
rect 200484 482240 203324 491760
rect 204084 482240 206924 491760
rect 207684 482240 210524 491760
rect 211284 482240 217724 491760
rect 218484 491760 224924 491808
rect 200484 482192 217724 482240
rect 218484 482240 221324 491760
rect 222084 482240 224924 491760
rect 218484 482192 224924 482240
rect 182484 422448 224924 482192
rect 182484 422400 199724 422448
rect 182484 412880 185324 422400
rect 186084 412880 188924 422400
rect 189684 412880 192524 422400
rect 193284 412880 199724 422400
rect 200484 422400 217724 422448
rect 182484 412832 199724 412880
rect 200484 412880 203324 422400
rect 204084 412880 206924 422400
rect 207684 412880 210524 422400
rect 211284 412880 217724 422400
rect 218484 422400 224924 422448
rect 200484 412832 217724 412880
rect 218484 412880 221324 422400
rect 222084 412880 224924 422400
rect 218484 412832 224924 412880
rect 182484 353088 224924 412832
rect 182484 353040 199724 353088
rect 182484 343520 185324 353040
rect 186084 343520 188924 353040
rect 189684 343520 192524 353040
rect 193284 343520 199724 353040
rect 200484 353040 217724 353088
rect 182484 343472 199724 343520
rect 200484 343520 203324 353040
rect 204084 343520 206924 353040
rect 207684 343520 210524 353040
rect 211284 343520 217724 353040
rect 218484 353040 224924 353088
rect 200484 343472 217724 343520
rect 218484 343520 221324 353040
rect 222084 343520 224924 353040
rect 218484 343472 224924 343520
rect 182484 283728 224924 343472
rect 182484 283680 199724 283728
rect 182484 274160 185324 283680
rect 186084 274160 188924 283680
rect 189684 274160 192524 283680
rect 193284 274160 199724 283680
rect 200484 283680 217724 283728
rect 182484 274112 199724 274160
rect 200484 274160 203324 283680
rect 204084 274160 206924 283680
rect 207684 274160 210524 283680
rect 211284 274160 217724 283680
rect 218484 283680 224924 283728
rect 200484 274112 217724 274160
rect 218484 274160 221324 283680
rect 222084 274160 224924 283680
rect 218484 274112 224924 274160
rect 182484 214368 224924 274112
rect 182484 214320 199724 214368
rect 182484 204800 185324 214320
rect 186084 204800 188924 214320
rect 189684 204800 192524 214320
rect 193284 204800 199724 214320
rect 200484 214320 217724 214368
rect 182484 204752 199724 204800
rect 200484 204800 203324 214320
rect 204084 204800 206924 214320
rect 207684 204800 210524 214320
rect 211284 204800 217724 214320
rect 218484 214320 224924 214368
rect 200484 204752 217724 204800
rect 218484 204800 221324 214320
rect 222084 204800 224924 214320
rect 218484 204752 224924 204800
rect 182484 145008 224924 204752
rect 182484 144960 199724 145008
rect 164484 132072 181724 132120
rect 182484 132120 185324 144960
rect 186084 132120 188924 144960
rect 189684 132120 192524 144960
rect 193284 132120 199724 144960
rect 200484 144960 217724 145008
rect 182484 132072 199724 132120
rect 200484 132120 203324 144960
rect 204084 132120 206924 144960
rect 207684 132120 210524 144960
rect 211284 132120 217724 144960
rect 218484 144960 224924 145008
rect 200484 132072 217724 132120
rect 218484 132120 221324 144960
rect 222084 132120 224924 144960
rect 225684 690320 228524 700501
rect 229284 690320 235724 700501
rect 225684 690272 235724 690320
rect 236484 690320 239324 700501
rect 240084 690320 242924 700501
rect 243684 690320 246524 700501
rect 247284 690320 253724 700501
rect 236484 690272 253724 690320
rect 254484 690320 257324 700501
rect 258084 690320 260924 700501
rect 261684 690320 264524 700501
rect 265284 690320 271724 700501
rect 254484 690272 271724 690320
rect 225684 630528 271724 690272
rect 225684 630480 235724 630528
rect 225684 620960 228524 630480
rect 229284 620960 235724 630480
rect 236484 630480 253724 630528
rect 225684 620912 235724 620960
rect 236484 620960 239324 630480
rect 240084 620960 242924 630480
rect 243684 620960 246524 630480
rect 247284 620960 253724 630480
rect 254484 630480 271724 630528
rect 236484 620912 253724 620960
rect 254484 620960 257324 630480
rect 258084 620960 260924 630480
rect 261684 620960 264524 630480
rect 265284 620960 271724 630480
rect 254484 620912 271724 620960
rect 225684 561168 271724 620912
rect 225684 561120 235724 561168
rect 225684 551600 228524 561120
rect 229284 551600 235724 561120
rect 236484 561120 253724 561168
rect 225684 551552 235724 551600
rect 236484 551600 239324 561120
rect 240084 551600 242924 561120
rect 243684 551600 246524 561120
rect 247284 551600 253724 561120
rect 254484 561120 271724 561168
rect 236484 551552 253724 551600
rect 254484 551600 257324 561120
rect 258084 551600 260924 561120
rect 261684 551600 264524 561120
rect 265284 551600 271724 561120
rect 254484 551552 271724 551600
rect 225684 491808 271724 551552
rect 225684 491760 235724 491808
rect 225684 482240 228524 491760
rect 229284 482240 235724 491760
rect 236484 491760 253724 491808
rect 225684 482192 235724 482240
rect 236484 482240 239324 491760
rect 240084 482240 242924 491760
rect 243684 482240 246524 491760
rect 247284 482240 253724 491760
rect 254484 491760 271724 491808
rect 236484 482192 253724 482240
rect 254484 482240 257324 491760
rect 258084 482240 260924 491760
rect 261684 482240 264524 491760
rect 265284 482240 271724 491760
rect 254484 482192 271724 482240
rect 225684 422448 271724 482192
rect 225684 422400 235724 422448
rect 225684 412880 228524 422400
rect 229284 412880 235724 422400
rect 236484 422400 253724 422448
rect 225684 412832 235724 412880
rect 236484 412880 239324 422400
rect 240084 412880 242924 422400
rect 243684 412880 246524 422400
rect 247284 412880 253724 422400
rect 254484 422400 271724 422448
rect 236484 412832 253724 412880
rect 254484 412880 257324 422400
rect 258084 412880 260924 422400
rect 261684 412880 264524 422400
rect 265284 412880 271724 422400
rect 254484 412832 271724 412880
rect 225684 353088 271724 412832
rect 225684 353040 235724 353088
rect 225684 343520 228524 353040
rect 229284 343520 235724 353040
rect 236484 353040 253724 353088
rect 225684 343472 235724 343520
rect 236484 343520 239324 353040
rect 240084 343520 242924 353040
rect 243684 343520 246524 353040
rect 247284 343520 253724 353040
rect 254484 353040 271724 353088
rect 236484 343472 253724 343520
rect 254484 343520 257324 353040
rect 258084 343520 260924 353040
rect 261684 343520 264524 353040
rect 265284 343520 271724 353040
rect 254484 343472 271724 343520
rect 225684 283728 271724 343472
rect 225684 283680 235724 283728
rect 225684 274160 228524 283680
rect 229284 274160 235724 283680
rect 236484 283680 253724 283728
rect 225684 274112 235724 274160
rect 236484 274160 239324 283680
rect 240084 274160 242924 283680
rect 243684 274160 246524 283680
rect 247284 274160 253724 283680
rect 254484 283680 271724 283728
rect 236484 274112 253724 274160
rect 254484 274160 257324 283680
rect 258084 274160 260924 283680
rect 261684 274160 264524 283680
rect 265284 274160 271724 283680
rect 254484 274112 271724 274160
rect 225684 214368 271724 274112
rect 225684 214320 235724 214368
rect 225684 204800 228524 214320
rect 229284 204800 235724 214320
rect 236484 214320 253724 214368
rect 225684 204752 235724 204800
rect 236484 204800 239324 214320
rect 240084 204800 242924 214320
rect 243684 204800 246524 214320
rect 247284 204800 253724 214320
rect 254484 214320 271724 214368
rect 236484 204752 253724 204800
rect 254484 204800 257324 214320
rect 258084 204800 260924 214320
rect 261684 204800 264524 214320
rect 265284 204800 271724 214320
rect 254484 204752 271724 204800
rect 225684 145008 271724 204752
rect 225684 144960 235724 145008
rect 225684 132120 228524 144960
rect 229284 132120 235724 144960
rect 236484 144960 253724 145008
rect 218484 132072 235724 132120
rect 164484 8328 235724 132072
rect 164484 8280 181724 8328
rect 164484 579 167324 8280
rect 168084 579 170924 8280
rect 171684 579 174524 8280
rect 175284 579 181724 8280
rect 182484 8280 199724 8328
rect 182484 579 185324 8280
rect 186084 579 188924 8280
rect 189684 579 192524 8280
rect 193284 579 199724 8280
rect 200484 8280 217724 8328
rect 200484 579 203324 8280
rect 204084 579 206924 8280
rect 207684 579 210524 8280
rect 211284 579 217724 8280
rect 218484 8280 235724 8328
rect 218484 579 221324 8280
rect 222084 579 224924 8280
rect 225684 579 228524 8280
rect 229284 579 235724 8280
rect 236484 132120 239324 144960
rect 240084 132120 242924 144960
rect 243684 132120 246524 144960
rect 247284 132120 253724 144960
rect 254484 144960 271724 145008
rect 236484 132072 253724 132120
rect 254484 132120 257324 144960
rect 258084 132120 260924 144960
rect 261684 132120 264524 144960
rect 265284 132120 271724 144960
rect 272484 690320 275324 700501
rect 276084 690320 278924 700501
rect 279684 690320 282524 700501
rect 283284 690320 289724 700501
rect 272484 690272 289724 690320
rect 290484 690320 293324 700501
rect 294084 690320 296924 700501
rect 297684 690320 300524 700501
rect 301284 690320 307724 700501
rect 290484 690272 307724 690320
rect 308484 690272 311324 700501
rect 272484 630528 311324 690272
rect 272484 630480 289724 630528
rect 272484 620960 275324 630480
rect 276084 620960 278924 630480
rect 279684 620960 282524 630480
rect 283284 620960 289724 630480
rect 290484 630480 307724 630528
rect 272484 620912 289724 620960
rect 290484 620960 293324 630480
rect 294084 620960 296924 630480
rect 297684 620960 300524 630480
rect 301284 620960 307724 630480
rect 290484 620912 307724 620960
rect 308484 620912 311324 630528
rect 272484 561168 311324 620912
rect 272484 561120 289724 561168
rect 272484 551600 275324 561120
rect 276084 551600 278924 561120
rect 279684 551600 282524 561120
rect 283284 551600 289724 561120
rect 290484 561120 307724 561168
rect 272484 551552 289724 551600
rect 290484 551600 293324 561120
rect 294084 551600 296924 561120
rect 297684 551600 300524 561120
rect 301284 551600 307724 561120
rect 290484 551552 307724 551600
rect 308484 551552 311324 561168
rect 272484 491808 311324 551552
rect 272484 491760 289724 491808
rect 272484 482240 275324 491760
rect 276084 482240 278924 491760
rect 279684 482240 282524 491760
rect 283284 482240 289724 491760
rect 290484 491760 307724 491808
rect 272484 482192 289724 482240
rect 290484 482240 293324 491760
rect 294084 482240 296924 491760
rect 297684 482240 300524 491760
rect 301284 482240 307724 491760
rect 290484 482192 307724 482240
rect 308484 482192 311324 491808
rect 272484 422448 311324 482192
rect 272484 422400 289724 422448
rect 272484 412880 275324 422400
rect 276084 412880 278924 422400
rect 279684 412880 282524 422400
rect 283284 412880 289724 422400
rect 290484 422400 307724 422448
rect 272484 412832 289724 412880
rect 290484 412880 293324 422400
rect 294084 412880 296924 422400
rect 297684 412880 300524 422400
rect 301284 412880 307724 422400
rect 290484 412832 307724 412880
rect 308484 412832 311324 422448
rect 272484 353088 311324 412832
rect 272484 353040 289724 353088
rect 272484 343520 275324 353040
rect 276084 343520 278924 353040
rect 279684 343520 282524 353040
rect 283284 343520 289724 353040
rect 290484 353040 307724 353088
rect 272484 343472 289724 343520
rect 290484 343520 293324 353040
rect 294084 343520 296924 353040
rect 297684 343520 300524 353040
rect 301284 343520 307724 353040
rect 290484 343472 307724 343520
rect 308484 343472 311324 353088
rect 272484 283728 311324 343472
rect 272484 283680 289724 283728
rect 272484 274160 275324 283680
rect 276084 274160 278924 283680
rect 279684 274160 282524 283680
rect 283284 274160 289724 283680
rect 290484 283680 307724 283728
rect 272484 274112 289724 274160
rect 290484 274160 293324 283680
rect 294084 274160 296924 283680
rect 297684 274160 300524 283680
rect 301284 274160 307724 283680
rect 290484 274112 307724 274160
rect 308484 274112 311324 283728
rect 272484 214368 311324 274112
rect 272484 214320 289724 214368
rect 272484 204800 275324 214320
rect 276084 204800 278924 214320
rect 279684 204800 282524 214320
rect 283284 204800 289724 214320
rect 290484 214320 307724 214368
rect 272484 204752 289724 204800
rect 290484 204800 293324 214320
rect 294084 204800 296924 214320
rect 297684 204800 300524 214320
rect 301284 204800 307724 214320
rect 290484 204752 307724 204800
rect 308484 204752 311324 214368
rect 272484 145008 311324 204752
rect 272484 144960 289724 145008
rect 254484 132072 271724 132120
rect 272484 132120 275324 144960
rect 276084 132120 278924 144960
rect 279684 132120 282524 144960
rect 283284 132120 289724 144960
rect 290484 144960 307724 145008
rect 272484 132072 289724 132120
rect 290484 132120 293324 144960
rect 294084 132120 296924 144960
rect 297684 132120 300524 144960
rect 301284 132120 307724 144960
rect 290484 132072 307724 132120
rect 236484 8328 307724 132072
rect 236484 8280 253724 8328
rect 236484 579 239324 8280
rect 240084 579 242924 8280
rect 243684 579 246524 8280
rect 247284 579 253724 8280
rect 254484 8280 271724 8328
rect 254484 579 257324 8280
rect 258084 579 260924 8280
rect 261684 579 264524 8280
rect 265284 579 271724 8280
rect 272484 8280 289724 8328
rect 272484 579 275324 8280
rect 276084 579 278924 8280
rect 279684 579 282524 8280
rect 283284 579 289724 8280
rect 290484 8280 307724 8328
rect 290484 579 293324 8280
rect 294084 579 296924 8280
rect 297684 579 300524 8280
rect 301284 579 307724 8280
rect 308484 132120 311324 145008
rect 312084 132120 314924 700501
rect 315684 690320 318524 700501
rect 319284 690320 325724 700501
rect 315684 690272 325724 690320
rect 326484 690320 329324 700501
rect 330084 690320 332924 700501
rect 333684 690320 336524 700501
rect 337284 690320 343724 700501
rect 326484 690272 343724 690320
rect 344484 690320 347324 700501
rect 348084 690320 350924 700501
rect 351684 690320 354524 700501
rect 355284 690320 361724 700501
rect 344484 690272 361724 690320
rect 362484 690320 365324 700501
rect 366084 690320 368924 700501
rect 369684 690320 372524 700501
rect 373284 690320 379724 700501
rect 362484 690272 379724 690320
rect 380484 690320 383324 700501
rect 384084 690320 386924 700501
rect 387684 690320 390524 700501
rect 391284 690320 397724 700501
rect 380484 690272 397724 690320
rect 398484 690272 401324 700501
rect 315684 630528 401324 690272
rect 315684 630480 325724 630528
rect 315684 620960 318524 630480
rect 319284 620960 325724 630480
rect 326484 630480 343724 630528
rect 315684 620912 325724 620960
rect 326484 620960 329324 630480
rect 330084 620960 332924 630480
rect 333684 620960 336524 630480
rect 337284 620960 343724 630480
rect 344484 630480 361724 630528
rect 326484 620912 343724 620960
rect 344484 620960 347324 630480
rect 348084 620960 350924 630480
rect 351684 620960 354524 630480
rect 355284 620960 361724 630480
rect 362484 630480 379724 630528
rect 344484 620912 361724 620960
rect 362484 620960 365324 630480
rect 366084 620960 368924 630480
rect 369684 620960 372524 630480
rect 373284 620960 379724 630480
rect 380484 630480 397724 630528
rect 362484 620912 379724 620960
rect 380484 620960 383324 630480
rect 384084 620960 386924 630480
rect 387684 620960 390524 630480
rect 391284 620960 397724 630480
rect 380484 620912 397724 620960
rect 398484 620912 401324 630528
rect 315684 561168 401324 620912
rect 315684 561120 325724 561168
rect 315684 551600 318524 561120
rect 319284 551600 325724 561120
rect 326484 561120 343724 561168
rect 315684 551552 325724 551600
rect 326484 551600 329324 561120
rect 330084 551600 332924 561120
rect 333684 551600 336524 561120
rect 337284 551600 343724 561120
rect 344484 561120 361724 561168
rect 326484 551552 343724 551600
rect 344484 551600 347324 561120
rect 348084 551600 350924 561120
rect 351684 551600 354524 561120
rect 355284 551600 361724 561120
rect 362484 561120 379724 561168
rect 344484 551552 361724 551600
rect 362484 551600 365324 561120
rect 366084 551600 368924 561120
rect 369684 551600 372524 561120
rect 373284 551600 379724 561120
rect 380484 561120 397724 561168
rect 362484 551552 379724 551600
rect 380484 551600 383324 561120
rect 384084 551600 386924 561120
rect 387684 551600 390524 561120
rect 391284 551600 397724 561120
rect 380484 551552 397724 551600
rect 398484 551552 401324 561168
rect 315684 491808 401324 551552
rect 315684 491760 325724 491808
rect 315684 482240 318524 491760
rect 319284 482240 325724 491760
rect 326484 491760 343724 491808
rect 315684 482192 325724 482240
rect 326484 482240 329324 491760
rect 330084 482240 332924 491760
rect 333684 482240 336524 491760
rect 337284 482240 343724 491760
rect 344484 491760 361724 491808
rect 326484 482192 343724 482240
rect 344484 482240 347324 491760
rect 348084 482240 350924 491760
rect 351684 482240 354524 491760
rect 355284 482240 361724 491760
rect 362484 491760 379724 491808
rect 344484 482192 361724 482240
rect 362484 482240 365324 491760
rect 366084 482240 368924 491760
rect 369684 482240 372524 491760
rect 373284 482240 379724 491760
rect 380484 491760 397724 491808
rect 362484 482192 379724 482240
rect 380484 482240 383324 491760
rect 384084 482240 386924 491760
rect 387684 482240 390524 491760
rect 391284 482240 397724 491760
rect 380484 482192 397724 482240
rect 398484 482192 401324 491808
rect 315684 422448 401324 482192
rect 315684 422400 325724 422448
rect 315684 412880 318524 422400
rect 319284 412880 325724 422400
rect 326484 422400 343724 422448
rect 315684 412832 325724 412880
rect 326484 412880 329324 422400
rect 330084 412880 332924 422400
rect 333684 412880 336524 422400
rect 337284 412880 343724 422400
rect 344484 422400 361724 422448
rect 326484 412832 343724 412880
rect 344484 412880 347324 422400
rect 348084 412880 350924 422400
rect 351684 412880 354524 422400
rect 355284 412880 361724 422400
rect 362484 422400 379724 422448
rect 344484 412832 361724 412880
rect 362484 412880 365324 422400
rect 366084 412880 368924 422400
rect 369684 412880 372524 422400
rect 373284 412880 379724 422400
rect 380484 422400 397724 422448
rect 362484 412832 379724 412880
rect 380484 412880 383324 422400
rect 384084 412880 386924 422400
rect 387684 412880 390524 422400
rect 391284 412880 397724 422400
rect 380484 412832 397724 412880
rect 398484 412832 401324 422448
rect 315684 353088 401324 412832
rect 315684 353040 325724 353088
rect 315684 343520 318524 353040
rect 319284 343520 325724 353040
rect 326484 353040 343724 353088
rect 315684 343472 325724 343520
rect 326484 343520 329324 353040
rect 330084 343520 332924 353040
rect 333684 343520 336524 353040
rect 337284 343520 343724 353040
rect 344484 353040 361724 353088
rect 326484 343472 343724 343520
rect 344484 343520 347324 353040
rect 348084 343520 350924 353040
rect 351684 343520 354524 353040
rect 355284 343520 361724 353040
rect 362484 353040 379724 353088
rect 344484 343472 361724 343520
rect 362484 343520 365324 353040
rect 366084 343520 368924 353040
rect 369684 343520 372524 353040
rect 373284 343520 379724 353040
rect 380484 353040 397724 353088
rect 362484 343472 379724 343520
rect 380484 343520 383324 353040
rect 384084 343520 386924 353040
rect 387684 343520 390524 353040
rect 391284 343520 397724 353040
rect 380484 343472 397724 343520
rect 398484 343472 401324 353088
rect 315684 283728 401324 343472
rect 315684 283680 325724 283728
rect 315684 274160 318524 283680
rect 319284 274160 325724 283680
rect 326484 283680 343724 283728
rect 315684 274112 325724 274160
rect 326484 274160 329324 283680
rect 330084 274160 332924 283680
rect 333684 274160 336524 283680
rect 337284 274160 343724 283680
rect 344484 283680 361724 283728
rect 326484 274112 343724 274160
rect 344484 274160 347324 283680
rect 348084 274160 350924 283680
rect 351684 274160 354524 283680
rect 355284 274160 361724 283680
rect 362484 283680 379724 283728
rect 344484 274112 361724 274160
rect 362484 274160 365324 283680
rect 366084 274160 368924 283680
rect 369684 274160 372524 283680
rect 373284 274160 379724 283680
rect 380484 283680 397724 283728
rect 362484 274112 379724 274160
rect 380484 274160 383324 283680
rect 384084 274160 386924 283680
rect 387684 274160 390524 283680
rect 391284 274160 397724 283680
rect 380484 274112 397724 274160
rect 398484 274112 401324 283728
rect 315684 214368 401324 274112
rect 315684 214320 325724 214368
rect 315684 204800 318524 214320
rect 319284 204800 325724 214320
rect 326484 214320 343724 214368
rect 315684 204752 325724 204800
rect 326484 204800 329324 214320
rect 330084 204800 332924 214320
rect 333684 204800 336524 214320
rect 337284 204800 343724 214320
rect 344484 214320 361724 214368
rect 326484 204752 343724 204800
rect 344484 204800 347324 214320
rect 348084 204800 350924 214320
rect 351684 204800 354524 214320
rect 355284 204800 361724 214320
rect 362484 214320 379724 214368
rect 344484 204752 361724 204800
rect 362484 204800 365324 214320
rect 366084 204800 368924 214320
rect 369684 204800 372524 214320
rect 373284 204800 379724 214320
rect 380484 214320 397724 214368
rect 362484 204752 379724 204800
rect 380484 204800 383324 214320
rect 384084 204800 386924 214320
rect 387684 204800 390524 214320
rect 391284 204800 397724 214320
rect 380484 204752 397724 204800
rect 398484 204752 401324 214368
rect 315684 145008 401324 204752
rect 315684 144960 325724 145008
rect 315684 132120 318524 144960
rect 319284 132120 325724 144960
rect 326484 144960 343724 145008
rect 308484 132072 325724 132120
rect 326484 132120 329324 144960
rect 330084 132120 332924 144960
rect 333684 132120 336524 144960
rect 337284 132120 343724 144960
rect 344484 144960 361724 145008
rect 326484 132072 343724 132120
rect 344484 132120 347324 144960
rect 348084 132120 350924 144960
rect 351684 132120 354524 144960
rect 355284 132120 361724 144960
rect 362484 144960 379724 145008
rect 344484 132072 361724 132120
rect 362484 132120 365324 144960
rect 366084 132120 368924 144960
rect 369684 132120 372524 144960
rect 373284 132120 379724 144960
rect 380484 144960 397724 145008
rect 362484 132072 379724 132120
rect 308484 8328 379724 132072
rect 308484 8280 325724 8328
rect 308484 579 311324 8280
rect 312084 579 314924 8280
rect 315684 579 318524 8280
rect 319284 579 325724 8280
rect 326484 8280 343724 8328
rect 326484 579 329324 8280
rect 330084 579 332924 8280
rect 333684 579 336524 8280
rect 337284 579 343724 8280
rect 344484 8280 361724 8328
rect 344484 579 347324 8280
rect 348084 579 350924 8280
rect 351684 579 354524 8280
rect 355284 579 361724 8280
rect 362484 8280 379724 8328
rect 362484 579 365324 8280
rect 366084 579 368924 8280
rect 369684 579 372524 8280
rect 373284 579 379724 8280
rect 380484 579 383324 144960
rect 384084 132120 386924 144960
rect 387684 132120 390524 144960
rect 391284 132120 397724 144960
rect 384084 132072 397724 132120
rect 398484 132120 401324 145008
rect 402084 690320 404924 700501
rect 405684 690320 408524 700501
rect 409284 690320 415724 700501
rect 402084 690272 415724 690320
rect 416484 690320 419324 700501
rect 420084 690320 422924 700501
rect 423684 690320 426524 700501
rect 427284 690320 433724 700501
rect 416484 690272 433724 690320
rect 434484 690320 437324 700501
rect 438084 690320 440924 700501
rect 441684 690320 444524 700501
rect 434484 690272 444524 690320
rect 402084 630528 444524 690272
rect 402084 630480 415724 630528
rect 402084 620960 404924 630480
rect 405684 620960 408524 630480
rect 409284 620960 415724 630480
rect 416484 630480 433724 630528
rect 402084 620912 415724 620960
rect 416484 620960 419324 630480
rect 420084 620960 422924 630480
rect 423684 620960 426524 630480
rect 427284 620960 433724 630480
rect 434484 630480 444524 630528
rect 416484 620912 433724 620960
rect 434484 620960 437324 630480
rect 438084 620960 440924 630480
rect 441684 620960 444524 630480
rect 434484 620912 444524 620960
rect 402084 561168 444524 620912
rect 402084 561120 415724 561168
rect 402084 551600 404924 561120
rect 405684 551600 408524 561120
rect 409284 551600 415724 561120
rect 416484 561120 433724 561168
rect 402084 551552 415724 551600
rect 416484 551600 419324 561120
rect 420084 551600 422924 561120
rect 423684 551600 426524 561120
rect 427284 551600 433724 561120
rect 434484 561120 444524 561168
rect 416484 551552 433724 551600
rect 434484 551600 437324 561120
rect 438084 551600 440924 561120
rect 441684 551600 444524 561120
rect 434484 551552 444524 551600
rect 402084 491808 444524 551552
rect 402084 491760 415724 491808
rect 402084 482240 404924 491760
rect 405684 482240 408524 491760
rect 409284 482240 415724 491760
rect 416484 491760 433724 491808
rect 402084 482192 415724 482240
rect 416484 482240 419324 491760
rect 420084 482240 422924 491760
rect 423684 482240 426524 491760
rect 427284 482240 433724 491760
rect 434484 491760 444524 491808
rect 416484 482192 433724 482240
rect 434484 482240 437324 491760
rect 438084 482240 440924 491760
rect 441684 482240 444524 491760
rect 434484 482192 444524 482240
rect 402084 422448 444524 482192
rect 402084 422400 415724 422448
rect 402084 412880 404924 422400
rect 405684 412880 408524 422400
rect 409284 412880 415724 422400
rect 416484 422400 433724 422448
rect 402084 412832 415724 412880
rect 416484 412880 419324 422400
rect 420084 412880 422924 422400
rect 423684 412880 426524 422400
rect 427284 412880 433724 422400
rect 434484 422400 444524 422448
rect 416484 412832 433724 412880
rect 434484 412880 437324 422400
rect 438084 412880 440924 422400
rect 441684 412880 444524 422400
rect 434484 412832 444524 412880
rect 402084 353088 444524 412832
rect 402084 353040 415724 353088
rect 402084 343520 404924 353040
rect 405684 343520 408524 353040
rect 409284 343520 415724 353040
rect 416484 353040 433724 353088
rect 402084 343472 415724 343520
rect 416484 343520 419324 353040
rect 420084 343520 422924 353040
rect 423684 343520 426524 353040
rect 427284 343520 433724 353040
rect 434484 353040 444524 353088
rect 416484 343472 433724 343520
rect 434484 343520 437324 353040
rect 438084 343520 440924 353040
rect 441684 343520 444524 353040
rect 434484 343472 444524 343520
rect 402084 283728 444524 343472
rect 402084 283680 415724 283728
rect 402084 274160 404924 283680
rect 405684 274160 408524 283680
rect 409284 274160 415724 283680
rect 416484 283680 433724 283728
rect 402084 274112 415724 274160
rect 416484 274160 419324 283680
rect 420084 274160 422924 283680
rect 423684 274160 426524 283680
rect 427284 274160 433724 283680
rect 434484 283680 444524 283728
rect 416484 274112 433724 274160
rect 434484 274160 437324 283680
rect 438084 274160 440924 283680
rect 441684 274160 444524 283680
rect 434484 274112 444524 274160
rect 402084 214368 444524 274112
rect 402084 214320 415724 214368
rect 402084 204800 404924 214320
rect 405684 204800 408524 214320
rect 409284 204800 415724 214320
rect 416484 214320 433724 214368
rect 402084 204752 415724 204800
rect 416484 204800 419324 214320
rect 420084 204800 422924 214320
rect 423684 204800 426524 214320
rect 427284 204800 433724 214320
rect 434484 214320 444524 214368
rect 416484 204752 433724 204800
rect 434484 204800 437324 214320
rect 438084 204800 440924 214320
rect 441684 204800 444524 214320
rect 434484 204752 444524 204800
rect 402084 145008 444524 204752
rect 402084 144960 415724 145008
rect 402084 132120 404924 144960
rect 405684 132120 408524 144960
rect 409284 132120 415724 144960
rect 416484 144960 433724 145008
rect 398484 132072 415724 132120
rect 416484 132120 419324 144960
rect 420084 132120 422924 144960
rect 423684 132120 426524 144960
rect 427284 132120 433724 144960
rect 434484 144960 444524 145008
rect 416484 132072 433724 132120
rect 434484 132120 437324 144960
rect 438084 132120 440924 144960
rect 441684 132120 444524 144960
rect 445284 690272 451724 700501
rect 452484 690320 455324 700501
rect 456084 690320 458924 700501
rect 459684 690320 462524 700501
rect 463284 690320 469724 700501
rect 452484 690272 469724 690320
rect 470484 690320 473324 700501
rect 474084 690320 476924 700501
rect 477684 690320 480524 700501
rect 481284 690320 487724 700501
rect 470484 690272 487724 690320
rect 445284 630528 487724 690272
rect 445284 620912 451724 630528
rect 452484 630480 469724 630528
rect 452484 620960 455324 630480
rect 456084 620960 458924 630480
rect 459684 620960 462524 630480
rect 463284 620960 469724 630480
rect 470484 630480 487724 630528
rect 452484 620912 469724 620960
rect 470484 620960 473324 630480
rect 474084 620960 476924 630480
rect 477684 620960 480524 630480
rect 481284 620960 487724 630480
rect 470484 620912 487724 620960
rect 445284 561168 487724 620912
rect 445284 551552 451724 561168
rect 452484 561120 469724 561168
rect 452484 551600 455324 561120
rect 456084 551600 458924 561120
rect 459684 551600 462524 561120
rect 463284 551600 469724 561120
rect 470484 561120 487724 561168
rect 452484 551552 469724 551600
rect 470484 551600 473324 561120
rect 474084 551600 476924 561120
rect 477684 551600 480524 561120
rect 481284 551600 487724 561120
rect 470484 551552 487724 551600
rect 445284 491808 487724 551552
rect 445284 482192 451724 491808
rect 452484 491760 469724 491808
rect 452484 482240 455324 491760
rect 456084 482240 458924 491760
rect 459684 482240 462524 491760
rect 463284 482240 469724 491760
rect 470484 491760 487724 491808
rect 452484 482192 469724 482240
rect 470484 482240 473324 491760
rect 474084 482240 476924 491760
rect 477684 482240 480524 491760
rect 481284 482240 487724 491760
rect 470484 482192 487724 482240
rect 445284 422448 487724 482192
rect 445284 412832 451724 422448
rect 452484 422400 469724 422448
rect 452484 412880 455324 422400
rect 456084 412880 458924 422400
rect 459684 412880 462524 422400
rect 463284 412880 469724 422400
rect 470484 422400 487724 422448
rect 452484 412832 469724 412880
rect 470484 412880 473324 422400
rect 474084 412880 476924 422400
rect 477684 412880 480524 422400
rect 481284 412880 487724 422400
rect 470484 412832 487724 412880
rect 445284 353088 487724 412832
rect 445284 343472 451724 353088
rect 452484 353040 469724 353088
rect 452484 343520 455324 353040
rect 456084 343520 458924 353040
rect 459684 343520 462524 353040
rect 463284 343520 469724 353040
rect 470484 353040 487724 353088
rect 452484 343472 469724 343520
rect 470484 343520 473324 353040
rect 474084 343520 476924 353040
rect 477684 343520 480524 353040
rect 481284 343520 487724 353040
rect 470484 343472 487724 343520
rect 445284 283728 487724 343472
rect 445284 274112 451724 283728
rect 452484 283680 469724 283728
rect 452484 274160 455324 283680
rect 456084 274160 458924 283680
rect 459684 274160 462524 283680
rect 463284 274160 469724 283680
rect 470484 283680 487724 283728
rect 452484 274112 469724 274160
rect 470484 274160 473324 283680
rect 474084 274160 476924 283680
rect 477684 274160 480524 283680
rect 481284 274160 487724 283680
rect 470484 274112 487724 274160
rect 445284 214368 487724 274112
rect 445284 204752 451724 214368
rect 452484 214320 469724 214368
rect 452484 204800 455324 214320
rect 456084 204800 458924 214320
rect 459684 204800 462524 214320
rect 463284 204800 469724 214320
rect 470484 214320 487724 214368
rect 452484 204752 469724 204800
rect 470484 204800 473324 214320
rect 474084 204800 476924 214320
rect 477684 204800 480524 214320
rect 481284 204800 487724 214320
rect 470484 204752 487724 204800
rect 445284 145008 487724 204752
rect 445284 132120 451724 145008
rect 452484 144960 469724 145008
rect 434484 132072 451724 132120
rect 452484 132120 455324 144960
rect 456084 132120 458924 144960
rect 459684 132120 462524 144960
rect 463284 132120 469724 144960
rect 470484 144960 487724 145008
rect 452484 132072 469724 132120
rect 470484 132120 473324 144960
rect 474084 132120 476924 144960
rect 477684 132120 480524 144960
rect 481284 132120 487724 144960
rect 470484 132072 487724 132120
rect 488484 132120 491324 700501
rect 492084 690320 494924 700501
rect 495684 690320 498524 700501
rect 499284 690320 505724 700501
rect 492084 690272 505724 690320
rect 506484 690320 509324 700501
rect 510084 690320 512924 700501
rect 513684 690320 516524 700501
rect 517284 690320 523724 700501
rect 506484 690272 523724 690320
rect 524484 690320 527324 700501
rect 528084 690320 530924 700501
rect 531684 690320 534524 700501
rect 524484 690272 534524 690320
rect 492084 630528 534524 690272
rect 492084 630480 505724 630528
rect 492084 620960 494924 630480
rect 495684 620960 498524 630480
rect 499284 620960 505724 630480
rect 506484 630480 523724 630528
rect 492084 620912 505724 620960
rect 506484 620960 509324 630480
rect 510084 620960 512924 630480
rect 513684 620960 516524 630480
rect 517284 620960 523724 630480
rect 524484 630480 534524 630528
rect 506484 620912 523724 620960
rect 524484 620960 527324 630480
rect 528084 620960 530924 630480
rect 531684 620960 534524 630480
rect 524484 620912 534524 620960
rect 492084 561168 534524 620912
rect 492084 561120 505724 561168
rect 492084 551600 494924 561120
rect 495684 551600 498524 561120
rect 499284 551600 505724 561120
rect 506484 561120 523724 561168
rect 492084 551552 505724 551600
rect 506484 551600 509324 561120
rect 510084 551600 512924 561120
rect 513684 551600 516524 561120
rect 517284 551600 523724 561120
rect 524484 561120 534524 561168
rect 506484 551552 523724 551600
rect 524484 551600 527324 561120
rect 528084 551600 530924 561120
rect 531684 551600 534524 561120
rect 524484 551552 534524 551600
rect 492084 491808 534524 551552
rect 492084 491760 505724 491808
rect 492084 482240 494924 491760
rect 495684 482240 498524 491760
rect 499284 482240 505724 491760
rect 506484 491760 523724 491808
rect 492084 482192 505724 482240
rect 506484 482240 509324 491760
rect 510084 482240 512924 491760
rect 513684 482240 516524 491760
rect 517284 482240 523724 491760
rect 524484 491760 534524 491808
rect 506484 482192 523724 482240
rect 524484 482240 527324 491760
rect 528084 482240 530924 491760
rect 531684 482240 534524 491760
rect 524484 482192 534524 482240
rect 492084 422448 534524 482192
rect 492084 422400 505724 422448
rect 492084 412880 494924 422400
rect 495684 412880 498524 422400
rect 499284 412880 505724 422400
rect 506484 422400 523724 422448
rect 492084 412832 505724 412880
rect 506484 412880 509324 422400
rect 510084 412880 512924 422400
rect 513684 412880 516524 422400
rect 517284 412880 523724 422400
rect 524484 422400 534524 422448
rect 506484 412832 523724 412880
rect 524484 412880 527324 422400
rect 528084 412880 530924 422400
rect 531684 412880 534524 422400
rect 524484 412832 534524 412880
rect 492084 353088 534524 412832
rect 492084 353040 505724 353088
rect 492084 343520 494924 353040
rect 495684 343520 498524 353040
rect 499284 343520 505724 353040
rect 506484 353040 523724 353088
rect 492084 343472 505724 343520
rect 506484 343520 509324 353040
rect 510084 343520 512924 353040
rect 513684 343520 516524 353040
rect 517284 343520 523724 353040
rect 524484 353040 534524 353088
rect 506484 343472 523724 343520
rect 524484 343520 527324 353040
rect 528084 343520 530924 353040
rect 531684 343520 534524 353040
rect 524484 343472 534524 343520
rect 492084 283728 534524 343472
rect 492084 283680 505724 283728
rect 492084 274160 494924 283680
rect 495684 274160 498524 283680
rect 499284 274160 505724 283680
rect 506484 283680 523724 283728
rect 492084 274112 505724 274160
rect 506484 274160 509324 283680
rect 510084 274160 512924 283680
rect 513684 274160 516524 283680
rect 517284 274160 523724 283680
rect 524484 283680 534524 283728
rect 506484 274112 523724 274160
rect 524484 274160 527324 283680
rect 528084 274160 530924 283680
rect 531684 274160 534524 283680
rect 524484 274112 534524 274160
rect 492084 214368 534524 274112
rect 492084 214320 505724 214368
rect 492084 204800 494924 214320
rect 495684 204800 498524 214320
rect 499284 204800 505724 214320
rect 506484 214320 523724 214368
rect 492084 204752 505724 204800
rect 506484 204800 509324 214320
rect 510084 204800 512924 214320
rect 513684 204800 516524 214320
rect 517284 204800 523724 214320
rect 524484 214320 534524 214368
rect 506484 204752 523724 204800
rect 524484 204800 527324 214320
rect 528084 204800 530924 214320
rect 531684 204800 534524 214320
rect 524484 204752 534524 204800
rect 492084 145008 534524 204752
rect 492084 144960 505724 145008
rect 492084 132120 494924 144960
rect 495684 132120 498524 144960
rect 499284 132120 505724 144960
rect 506484 144960 523724 145008
rect 488484 132072 505724 132120
rect 506484 132120 509324 144960
rect 510084 132120 512924 144960
rect 513684 132120 516524 144960
rect 517284 132120 523724 144960
rect 524484 144960 534524 145008
rect 506484 132072 523724 132120
rect 524484 132120 527324 144960
rect 528084 132120 530924 144960
rect 531684 132120 534524 144960
rect 535284 690272 541724 700501
rect 542484 690320 545324 700501
rect 546084 690320 548924 700501
rect 549684 690320 552524 700501
rect 553284 690320 559724 700501
rect 542484 690272 559724 690320
rect 560484 690320 563324 700501
rect 564084 690320 566924 700501
rect 567684 690320 570524 700501
rect 571284 690320 577724 700501
rect 560484 690272 577724 690320
rect 535284 630528 577724 690272
rect 535284 620912 541724 630528
rect 542484 630480 559724 630528
rect 542484 620960 545324 630480
rect 546084 620960 548924 630480
rect 549684 620960 552524 630480
rect 553284 620960 559724 630480
rect 560484 630480 577724 630528
rect 542484 620912 559724 620960
rect 560484 620960 563324 630480
rect 564084 620960 566924 630480
rect 567684 620960 570524 630480
rect 571284 620960 577724 630480
rect 560484 620912 577724 620960
rect 535284 561168 577724 620912
rect 535284 551552 541724 561168
rect 542484 561120 559724 561168
rect 542484 551600 545324 561120
rect 546084 551600 548924 561120
rect 549684 551600 552524 561120
rect 553284 551600 559724 561120
rect 560484 561120 577724 561168
rect 542484 551552 559724 551600
rect 560484 551600 563324 561120
rect 564084 551600 566924 561120
rect 567684 551600 570524 561120
rect 571284 551600 577724 561120
rect 560484 551552 577724 551600
rect 535284 491808 577724 551552
rect 535284 482192 541724 491808
rect 542484 491760 559724 491808
rect 542484 482240 545324 491760
rect 546084 482240 548924 491760
rect 549684 482240 552524 491760
rect 553284 482240 559724 491760
rect 560484 491760 577724 491808
rect 542484 482192 559724 482240
rect 560484 482240 563324 491760
rect 564084 482240 566924 491760
rect 567684 482240 570524 491760
rect 571284 482240 577724 491760
rect 560484 482192 577724 482240
rect 535284 422448 577724 482192
rect 535284 412832 541724 422448
rect 542484 422400 559724 422448
rect 542484 412880 545324 422400
rect 546084 412880 548924 422400
rect 549684 412880 552524 422400
rect 553284 412880 559724 422400
rect 560484 422400 577724 422448
rect 542484 412832 559724 412880
rect 560484 412880 563324 422400
rect 564084 412880 566924 422400
rect 567684 412880 570524 422400
rect 571284 412880 577724 422400
rect 560484 412832 577724 412880
rect 535284 353088 577724 412832
rect 535284 343472 541724 353088
rect 542484 353040 559724 353088
rect 542484 343520 545324 353040
rect 546084 343520 548924 353040
rect 549684 343520 552524 353040
rect 553284 343520 559724 353040
rect 560484 353040 577724 353088
rect 542484 343472 559724 343520
rect 560484 343520 563324 353040
rect 564084 343520 566924 353040
rect 567684 343520 570524 353040
rect 571284 343520 577724 353040
rect 560484 343472 577724 343520
rect 535284 283728 577724 343472
rect 535284 274112 541724 283728
rect 542484 283680 559724 283728
rect 542484 274160 545324 283680
rect 546084 274160 548924 283680
rect 549684 274160 552524 283680
rect 553284 274160 559724 283680
rect 560484 283680 577724 283728
rect 542484 274112 559724 274160
rect 560484 274160 563324 283680
rect 564084 274160 566924 283680
rect 567684 274160 570524 283680
rect 571284 274160 577724 283680
rect 560484 274112 577724 274160
rect 535284 214368 577724 274112
rect 535284 204752 541724 214368
rect 542484 214320 559724 214368
rect 542484 204800 545324 214320
rect 546084 204800 548924 214320
rect 549684 204800 552524 214320
rect 553284 204800 559724 214320
rect 560484 214320 577724 214368
rect 542484 204752 559724 204800
rect 560484 204800 563324 214320
rect 564084 204800 566924 214320
rect 567684 204800 570524 214320
rect 571284 204800 577724 214320
rect 560484 204752 577724 204800
rect 535284 145008 577724 204752
rect 535284 132120 541724 145008
rect 542484 144960 559724 145008
rect 524484 132072 541724 132120
rect 542484 132120 545324 144960
rect 546084 132120 548924 144960
rect 549684 132120 552524 144960
rect 553284 132120 559724 144960
rect 560484 144960 577724 145008
rect 542484 132072 559724 132120
rect 560484 132120 563324 144960
rect 564084 132120 566924 144960
rect 567684 132120 570524 144960
rect 560484 132072 570524 132120
rect 384084 8328 570524 132072
rect 384084 8280 397724 8328
rect 384084 579 386924 8280
rect 387684 579 390524 8280
rect 391284 579 397724 8280
rect 398484 8280 415724 8328
rect 398484 579 401324 8280
rect 402084 579 404924 8280
rect 405684 579 408524 8280
rect 409284 579 415724 8280
rect 416484 8280 433724 8328
rect 416484 579 419324 8280
rect 420084 579 422924 8280
rect 423684 579 426524 8280
rect 427284 579 433724 8280
rect 434484 8280 451724 8328
rect 434484 579 437324 8280
rect 438084 579 440924 8280
rect 441684 579 444524 8280
rect 445284 579 451724 8280
rect 452484 8280 469724 8328
rect 452484 579 455324 8280
rect 456084 579 458924 8280
rect 459684 579 462524 8280
rect 463284 579 469724 8280
rect 470484 8280 487724 8328
rect 470484 579 473324 8280
rect 474084 579 476924 8280
rect 477684 579 480524 8280
rect 481284 579 487724 8280
rect 488484 8280 505724 8328
rect 488484 579 491324 8280
rect 492084 579 494924 8280
rect 495684 579 498524 8280
rect 499284 579 505724 8280
rect 506484 8280 523724 8328
rect 506484 579 509324 8280
rect 510084 579 512924 8280
rect 513684 579 516524 8280
rect 517284 579 523724 8280
rect 524484 8280 541724 8328
rect 524484 579 527324 8280
rect 528084 579 530924 8280
rect 531684 579 534524 8280
rect 535284 579 541724 8280
rect 542484 8280 559724 8328
rect 542484 579 545324 8280
rect 546084 579 548924 8280
rect 549684 579 552524 8280
rect 553284 579 559724 8280
rect 560484 8280 570524 8328
rect 560484 579 563324 8280
rect 564084 579 566924 8280
rect 567684 579 570524 8280
rect 571284 579 577724 144960
rect 578484 579 580277 700501
<< metal5 >>
rect -8576 710840 592500 711440
rect -7636 709900 591560 710500
rect -6696 708960 590620 709560
rect -5756 708020 589680 708620
rect -4816 707080 588740 707680
rect -3876 706140 587800 706740
rect -2936 705200 586860 705800
rect -1996 704260 585920 704860
rect -8576 697676 592500 698276
rect -6696 694076 590620 694676
rect -4816 690476 588740 691076
rect -2936 686828 586860 687428
rect -8576 679676 592500 680276
rect -6696 676076 590620 676676
rect -4816 672476 588740 673076
rect -2936 668828 586860 669428
rect -8576 661676 592500 662276
rect -6696 658076 590620 658676
rect -4816 654476 588740 655076
rect -2936 650828 586860 651428
rect -8576 643676 592500 644276
rect -6696 640076 590620 640676
rect -4816 636476 588740 637076
rect -2936 632828 586860 633428
rect -8576 625676 592500 626276
rect -6696 622076 590620 622676
rect -4816 618476 588740 619076
rect -2936 614828 586860 615428
rect -8576 607676 592500 608276
rect -6696 604076 590620 604676
rect -4816 600476 588740 601076
rect -2936 596828 586860 597428
rect -8576 589676 592500 590276
rect -6696 586076 590620 586676
rect -4816 582476 588740 583076
rect -2936 578828 586860 579428
rect -8576 571676 592500 572276
rect -6696 568076 590620 568676
rect -4816 564476 588740 565076
rect -2936 560828 586860 561428
rect -8576 553676 592500 554276
rect -6696 550076 590620 550676
rect -4816 546476 588740 547076
rect -2936 542828 586860 543428
rect -8576 535676 592500 536276
rect -6696 532076 590620 532676
rect -4816 528476 588740 529076
rect -2936 524828 586860 525428
rect -8576 517676 592500 518276
rect -6696 514076 590620 514676
rect -4816 510476 588740 511076
rect -2936 506828 586860 507428
rect -8576 499676 592500 500276
rect -6696 496076 590620 496676
rect -4816 492476 588740 493076
rect -2936 488828 586860 489428
rect -8576 481676 592500 482276
rect -6696 478076 590620 478676
rect -4816 474476 588740 475076
rect -2936 470828 586860 471428
rect -8576 463676 592500 464276
rect -6696 460076 590620 460676
rect -4816 456476 588740 457076
rect -2936 452828 586860 453428
rect -8576 445676 592500 446276
rect -6696 442076 590620 442676
rect -4816 438476 588740 439076
rect -2936 434828 586860 435428
rect -8576 427676 592500 428276
rect -6696 424076 590620 424676
rect -4816 420476 588740 421076
rect -2936 416828 586860 417428
rect -8576 409676 592500 410276
rect -6696 406076 590620 406676
rect -4816 402476 588740 403076
rect -2936 398828 586860 399428
rect -8576 391676 592500 392276
rect -6696 388076 590620 388676
rect -4816 384476 588740 385076
rect -2936 380828 586860 381428
rect -8576 373676 592500 374276
rect -6696 370076 590620 370676
rect -4816 366476 588740 367076
rect -2936 362828 586860 363428
rect -8576 355676 592500 356276
rect -6696 352076 590620 352676
rect -4816 348476 588740 349076
rect -2936 344828 586860 345428
rect -8576 337676 592500 338276
rect -6696 334076 590620 334676
rect -4816 330476 588740 331076
rect -2936 326828 586860 327428
rect -8576 319676 592500 320276
rect -6696 316076 590620 316676
rect -4816 312476 588740 313076
rect -2936 308828 586860 309428
rect -8576 301676 592500 302276
rect -6696 298076 590620 298676
rect -4816 294476 588740 295076
rect -2936 290828 586860 291428
rect -8576 283676 592500 284276
rect -6696 280076 590620 280676
rect -4816 276476 588740 277076
rect -2936 272828 586860 273428
rect -8576 265676 592500 266276
rect -6696 262076 590620 262676
rect -4816 258476 588740 259076
rect -2936 254828 586860 255428
rect -8576 247676 592500 248276
rect -6696 244076 590620 244676
rect -4816 240476 588740 241076
rect -2936 236828 586860 237428
rect -8576 229676 592500 230276
rect -6696 226076 590620 226676
rect -4816 222476 588740 223076
rect -2936 218828 586860 219428
rect -8576 211676 592500 212276
rect -6696 208076 590620 208676
rect -4816 204476 588740 205076
rect -2936 200828 586860 201428
rect -8576 193676 592500 194276
rect -6696 190076 590620 190676
rect -4816 186476 588740 187076
rect -2936 182828 586860 183428
rect -8576 175676 592500 176276
rect -6696 172076 590620 172676
rect -4816 168476 588740 169076
rect -2936 164828 586860 165428
rect -8576 157676 592500 158276
rect -6696 154076 590620 154676
rect -4816 150476 588740 151076
rect -2936 146828 586860 147428
rect -8576 139676 592500 140276
rect -6696 136076 590620 136676
rect -4816 132476 588740 133076
rect -2936 128828 586860 129428
rect -8576 121676 592500 122276
rect -6696 118076 590620 118676
rect -4816 114476 588740 115076
rect -2936 110828 586860 111428
rect -8576 103676 592500 104276
rect -6696 100076 590620 100676
rect -4816 96476 588740 97076
rect -2936 92828 586860 93428
rect -8576 85676 592500 86276
rect -6696 82076 590620 82676
rect -4816 78476 588740 79076
rect -2936 74828 586860 75428
rect -8576 67676 592500 68276
rect -6696 64076 590620 64676
rect -4816 60476 588740 61076
rect -2936 56828 586860 57428
rect -8576 49676 592500 50276
rect -6696 46076 590620 46676
rect -4816 42476 588740 43076
rect -2936 38828 586860 39428
rect -8576 31676 592500 32276
rect -6696 28076 590620 28676
rect -4816 24476 588740 25076
rect -2936 20828 586860 21428
rect -8576 13676 592500 14276
rect -6696 10076 590620 10676
rect -4816 6476 588740 7076
rect -2936 2828 586860 3428
rect -1996 -924 585920 -324
rect -2936 -1864 586860 -1264
rect -3876 -2804 587800 -2204
rect -4816 -3744 588740 -3144
rect -5756 -4684 589680 -4084
rect -6696 -5624 590620 -5024
rect -7636 -6564 591560 -5964
rect -8576 -7504 592500 -6904
<< obsm5 >>
rect -8576 711440 -7976 711442
rect 30604 711440 31204 711442
rect 66604 711440 67204 711442
rect 102604 711440 103204 711442
rect 138604 711440 139204 711442
rect 174604 711440 175204 711442
rect 210604 711440 211204 711442
rect 246604 711440 247204 711442
rect 282604 711440 283204 711442
rect 318604 711440 319204 711442
rect 354604 711440 355204 711442
rect 390604 711440 391204 711442
rect 426604 711440 427204 711442
rect 462604 711440 463204 711442
rect 498604 711440 499204 711442
rect 534604 711440 535204 711442
rect 570604 711440 571204 711442
rect 591900 711440 592500 711442
rect -8576 710838 -7976 710840
rect 30604 710838 31204 710840
rect 66604 710838 67204 710840
rect 102604 710838 103204 710840
rect 138604 710838 139204 710840
rect 174604 710838 175204 710840
rect 210604 710838 211204 710840
rect 246604 710838 247204 710840
rect 282604 710838 283204 710840
rect 318604 710838 319204 710840
rect 354604 710838 355204 710840
rect 390604 710838 391204 710840
rect 426604 710838 427204 710840
rect 462604 710838 463204 710840
rect 498604 710838 499204 710840
rect 534604 710838 535204 710840
rect 570604 710838 571204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 12604 710500 13204 710502
rect 48604 710500 49204 710502
rect 84604 710500 85204 710502
rect 120604 710500 121204 710502
rect 156604 710500 157204 710502
rect 192604 710500 193204 710502
rect 228604 710500 229204 710502
rect 264604 710500 265204 710502
rect 300604 710500 301204 710502
rect 336604 710500 337204 710502
rect 372604 710500 373204 710502
rect 408604 710500 409204 710502
rect 444604 710500 445204 710502
rect 480604 710500 481204 710502
rect 516604 710500 517204 710502
rect 552604 710500 553204 710502
rect 590960 710500 591560 710502
rect -7636 709898 -7036 709900
rect 12604 709898 13204 709900
rect 48604 709898 49204 709900
rect 84604 709898 85204 709900
rect 120604 709898 121204 709900
rect 156604 709898 157204 709900
rect 192604 709898 193204 709900
rect 228604 709898 229204 709900
rect 264604 709898 265204 709900
rect 300604 709898 301204 709900
rect 336604 709898 337204 709900
rect 372604 709898 373204 709900
rect 408604 709898 409204 709900
rect 444604 709898 445204 709900
rect 480604 709898 481204 709900
rect 516604 709898 517204 709900
rect 552604 709898 553204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 27004 709560 27604 709562
rect 63004 709560 63604 709562
rect 99004 709560 99604 709562
rect 135004 709560 135604 709562
rect 171004 709560 171604 709562
rect 207004 709560 207604 709562
rect 243004 709560 243604 709562
rect 279004 709560 279604 709562
rect 315004 709560 315604 709562
rect 351004 709560 351604 709562
rect 387004 709560 387604 709562
rect 423004 709560 423604 709562
rect 459004 709560 459604 709562
rect 495004 709560 495604 709562
rect 531004 709560 531604 709562
rect 567004 709560 567604 709562
rect 590020 709560 590620 709562
rect -6696 708958 -6096 708960
rect 27004 708958 27604 708960
rect 63004 708958 63604 708960
rect 99004 708958 99604 708960
rect 135004 708958 135604 708960
rect 171004 708958 171604 708960
rect 207004 708958 207604 708960
rect 243004 708958 243604 708960
rect 279004 708958 279604 708960
rect 315004 708958 315604 708960
rect 351004 708958 351604 708960
rect 387004 708958 387604 708960
rect 423004 708958 423604 708960
rect 459004 708958 459604 708960
rect 495004 708958 495604 708960
rect 531004 708958 531604 708960
rect 567004 708958 567604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 9004 708620 9604 708622
rect 45004 708620 45604 708622
rect 81004 708620 81604 708622
rect 117004 708620 117604 708622
rect 153004 708620 153604 708622
rect 189004 708620 189604 708622
rect 225004 708620 225604 708622
rect 261004 708620 261604 708622
rect 297004 708620 297604 708622
rect 333004 708620 333604 708622
rect 369004 708620 369604 708622
rect 405004 708620 405604 708622
rect 441004 708620 441604 708622
rect 477004 708620 477604 708622
rect 513004 708620 513604 708622
rect 549004 708620 549604 708622
rect 589080 708620 589680 708622
rect -5756 708018 -5156 708020
rect 9004 708018 9604 708020
rect 45004 708018 45604 708020
rect 81004 708018 81604 708020
rect 117004 708018 117604 708020
rect 153004 708018 153604 708020
rect 189004 708018 189604 708020
rect 225004 708018 225604 708020
rect 261004 708018 261604 708020
rect 297004 708018 297604 708020
rect 333004 708018 333604 708020
rect 369004 708018 369604 708020
rect 405004 708018 405604 708020
rect 441004 708018 441604 708020
rect 477004 708018 477604 708020
rect 513004 708018 513604 708020
rect 549004 708018 549604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 23404 707680 24004 707682
rect 59404 707680 60004 707682
rect 95404 707680 96004 707682
rect 131404 707680 132004 707682
rect 167404 707680 168004 707682
rect 203404 707680 204004 707682
rect 239404 707680 240004 707682
rect 275404 707680 276004 707682
rect 311404 707680 312004 707682
rect 347404 707680 348004 707682
rect 383404 707680 384004 707682
rect 419404 707680 420004 707682
rect 455404 707680 456004 707682
rect 491404 707680 492004 707682
rect 527404 707680 528004 707682
rect 563404 707680 564004 707682
rect 588140 707680 588740 707682
rect -4816 707078 -4216 707080
rect 23404 707078 24004 707080
rect 59404 707078 60004 707080
rect 95404 707078 96004 707080
rect 131404 707078 132004 707080
rect 167404 707078 168004 707080
rect 203404 707078 204004 707080
rect 239404 707078 240004 707080
rect 275404 707078 276004 707080
rect 311404 707078 312004 707080
rect 347404 707078 348004 707080
rect 383404 707078 384004 707080
rect 419404 707078 420004 707080
rect 455404 707078 456004 707080
rect 491404 707078 492004 707080
rect 527404 707078 528004 707080
rect 563404 707078 564004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 5404 706740 6004 706742
rect 41404 706740 42004 706742
rect 77404 706740 78004 706742
rect 113404 706740 114004 706742
rect 149404 706740 150004 706742
rect 185404 706740 186004 706742
rect 221404 706740 222004 706742
rect 257404 706740 258004 706742
rect 293404 706740 294004 706742
rect 329404 706740 330004 706742
rect 365404 706740 366004 706742
rect 401404 706740 402004 706742
rect 437404 706740 438004 706742
rect 473404 706740 474004 706742
rect 509404 706740 510004 706742
rect 545404 706740 546004 706742
rect 581404 706740 582004 706742
rect 587200 706740 587800 706742
rect -3876 706138 -3276 706140
rect 5404 706138 6004 706140
rect 41404 706138 42004 706140
rect 77404 706138 78004 706140
rect 113404 706138 114004 706140
rect 149404 706138 150004 706140
rect 185404 706138 186004 706140
rect 221404 706138 222004 706140
rect 257404 706138 258004 706140
rect 293404 706138 294004 706140
rect 329404 706138 330004 706140
rect 365404 706138 366004 706140
rect 401404 706138 402004 706140
rect 437404 706138 438004 706140
rect 473404 706138 474004 706140
rect 509404 706138 510004 706140
rect 545404 706138 546004 706140
rect 581404 706138 582004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 19804 705800 20404 705802
rect 55804 705800 56404 705802
rect 91804 705800 92404 705802
rect 127804 705800 128404 705802
rect 163804 705800 164404 705802
rect 199804 705800 200404 705802
rect 235804 705800 236404 705802
rect 271804 705800 272404 705802
rect 307804 705800 308404 705802
rect 343804 705800 344404 705802
rect 379804 705800 380404 705802
rect 415804 705800 416404 705802
rect 451804 705800 452404 705802
rect 487804 705800 488404 705802
rect 523804 705800 524404 705802
rect 559804 705800 560404 705802
rect 586260 705800 586860 705802
rect -2936 705198 -2336 705200
rect 19804 705198 20404 705200
rect 55804 705198 56404 705200
rect 91804 705198 92404 705200
rect 127804 705198 128404 705200
rect 163804 705198 164404 705200
rect 199804 705198 200404 705200
rect 235804 705198 236404 705200
rect 271804 705198 272404 705200
rect 307804 705198 308404 705200
rect 343804 705198 344404 705200
rect 379804 705198 380404 705200
rect 415804 705198 416404 705200
rect 451804 705198 452404 705200
rect 487804 705198 488404 705200
rect 523804 705198 524404 705200
rect 559804 705198 560404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 1804 704860 2404 704862
rect 37804 704860 38404 704862
rect 73804 704860 74404 704862
rect 109804 704860 110404 704862
rect 145804 704860 146404 704862
rect 181804 704860 182404 704862
rect 217804 704860 218404 704862
rect 253804 704860 254404 704862
rect 289804 704860 290404 704862
rect 325804 704860 326404 704862
rect 361804 704860 362404 704862
rect 397804 704860 398404 704862
rect 433804 704860 434404 704862
rect 469804 704860 470404 704862
rect 505804 704860 506404 704862
rect 541804 704860 542404 704862
rect 577804 704860 578404 704862
rect 585320 704860 585920 704862
rect -1996 704258 -1396 704260
rect 1804 704258 2404 704260
rect 37804 704258 38404 704260
rect 73804 704258 74404 704260
rect 109804 704258 110404 704260
rect 145804 704258 146404 704260
rect 181804 704258 182404 704260
rect 217804 704258 218404 704260
rect 253804 704258 254404 704260
rect 289804 704258 290404 704260
rect 325804 704258 326404 704260
rect 361804 704258 362404 704260
rect 397804 704258 398404 704260
rect 433804 704258 434404 704260
rect 469804 704258 470404 704260
rect 505804 704258 506404 704260
rect 541804 704258 542404 704260
rect 577804 704258 578404 704260
rect 585320 704258 585920 704260
rect 0 698596 584000 703940
rect -7636 698276 -7036 698278
rect 590960 698276 591560 698278
rect -7636 697674 -7036 697676
rect 590960 697674 591560 697676
rect 0 694996 584000 697356
rect -5756 694676 -5156 694678
rect 589080 694676 589680 694678
rect -5756 694074 -5156 694076
rect 589080 694074 589680 694076
rect 0 691396 584000 693756
rect -3876 691076 -3276 691078
rect 587200 691076 587800 691078
rect -3876 690474 -3276 690476
rect 587200 690474 587800 690476
rect 0 687748 584000 690156
rect -1996 687428 -1396 687430
rect 585320 687428 585920 687430
rect -1996 686826 -1396 686828
rect 585320 686826 585920 686828
rect 0 680596 584000 686508
rect -8576 680276 -7976 680278
rect 591900 680276 592500 680278
rect -8576 679674 -7976 679676
rect 591900 679674 592500 679676
rect 0 676996 584000 679356
rect -6696 676676 -6096 676678
rect 590020 676676 590620 676678
rect -6696 676074 -6096 676076
rect 590020 676074 590620 676076
rect 0 673396 584000 675756
rect -4816 673076 -4216 673078
rect 588140 673076 588740 673078
rect -4816 672474 -4216 672476
rect 588140 672474 588740 672476
rect 0 669748 584000 672156
rect -2936 669428 -2336 669430
rect 586260 669428 586860 669430
rect -2936 668826 -2336 668828
rect 586260 668826 586860 668828
rect 0 662596 584000 668508
rect -7636 662276 -7036 662278
rect 590960 662276 591560 662278
rect -7636 661674 -7036 661676
rect 590960 661674 591560 661676
rect 0 658996 584000 661356
rect -5756 658676 -5156 658678
rect 589080 658676 589680 658678
rect -5756 658074 -5156 658076
rect 589080 658074 589680 658076
rect 0 655396 584000 657756
rect -3876 655076 -3276 655078
rect 587200 655076 587800 655078
rect -3876 654474 -3276 654476
rect 587200 654474 587800 654476
rect 0 651748 584000 654156
rect -1996 651428 -1396 651430
rect 585320 651428 585920 651430
rect -1996 650826 -1396 650828
rect 585320 650826 585920 650828
rect 0 644596 584000 650508
rect -8576 644276 -7976 644278
rect 591900 644276 592500 644278
rect -8576 643674 -7976 643676
rect 591900 643674 592500 643676
rect 0 640996 584000 643356
rect -6696 640676 -6096 640678
rect 590020 640676 590620 640678
rect -6696 640074 -6096 640076
rect 590020 640074 590620 640076
rect 0 637396 584000 639756
rect -4816 637076 -4216 637078
rect 588140 637076 588740 637078
rect -4816 636474 -4216 636476
rect 588140 636474 588740 636476
rect 0 633748 584000 636156
rect -2936 633428 -2336 633430
rect 586260 633428 586860 633430
rect -2936 632826 -2336 632828
rect 586260 632826 586860 632828
rect 0 626596 584000 632508
rect -7636 626276 -7036 626278
rect 590960 626276 591560 626278
rect -7636 625674 -7036 625676
rect 590960 625674 591560 625676
rect 0 622996 584000 625356
rect -5756 622676 -5156 622678
rect 589080 622676 589680 622678
rect -5756 622074 -5156 622076
rect 589080 622074 589680 622076
rect 0 619396 584000 621756
rect -3876 619076 -3276 619078
rect 587200 619076 587800 619078
rect -3876 618474 -3276 618476
rect 587200 618474 587800 618476
rect 0 615748 584000 618156
rect -1996 615428 -1396 615430
rect 585320 615428 585920 615430
rect -1996 614826 -1396 614828
rect 585320 614826 585920 614828
rect 0 608596 584000 614508
rect -8576 608276 -7976 608278
rect 591900 608276 592500 608278
rect -8576 607674 -7976 607676
rect 591900 607674 592500 607676
rect 0 604996 584000 607356
rect -6696 604676 -6096 604678
rect 590020 604676 590620 604678
rect -6696 604074 -6096 604076
rect 590020 604074 590620 604076
rect 0 601396 584000 603756
rect -4816 601076 -4216 601078
rect 588140 601076 588740 601078
rect -4816 600474 -4216 600476
rect 588140 600474 588740 600476
rect 0 597748 584000 600156
rect -2936 597428 -2336 597430
rect 586260 597428 586860 597430
rect -2936 596826 -2336 596828
rect 586260 596826 586860 596828
rect 0 590596 584000 596508
rect -7636 590276 -7036 590278
rect 590960 590276 591560 590278
rect -7636 589674 -7036 589676
rect 590960 589674 591560 589676
rect 0 586996 584000 589356
rect -5756 586676 -5156 586678
rect 589080 586676 589680 586678
rect -5756 586074 -5156 586076
rect 589080 586074 589680 586076
rect 0 583396 584000 585756
rect -3876 583076 -3276 583078
rect 587200 583076 587800 583078
rect -3876 582474 -3276 582476
rect 587200 582474 587800 582476
rect 0 579748 584000 582156
rect -1996 579428 -1396 579430
rect 585320 579428 585920 579430
rect -1996 578826 -1396 578828
rect 585320 578826 585920 578828
rect 0 572596 584000 578508
rect -8576 572276 -7976 572278
rect 591900 572276 592500 572278
rect -8576 571674 -7976 571676
rect 591900 571674 592500 571676
rect 0 568996 584000 571356
rect -6696 568676 -6096 568678
rect 590020 568676 590620 568678
rect -6696 568074 -6096 568076
rect 590020 568074 590620 568076
rect 0 565396 584000 567756
rect -4816 565076 -4216 565078
rect 588140 565076 588740 565078
rect -4816 564474 -4216 564476
rect 588140 564474 588740 564476
rect 0 561748 584000 564156
rect -2936 561428 -2336 561430
rect 586260 561428 586860 561430
rect -2936 560826 -2336 560828
rect 586260 560826 586860 560828
rect 0 554596 584000 560508
rect -7636 554276 -7036 554278
rect 590960 554276 591560 554278
rect -7636 553674 -7036 553676
rect 590960 553674 591560 553676
rect 0 550996 584000 553356
rect -5756 550676 -5156 550678
rect 589080 550676 589680 550678
rect -5756 550074 -5156 550076
rect 589080 550074 589680 550076
rect 0 547396 584000 549756
rect -3876 547076 -3276 547078
rect 587200 547076 587800 547078
rect -3876 546474 -3276 546476
rect 587200 546474 587800 546476
rect 0 543748 584000 546156
rect -1996 543428 -1396 543430
rect 585320 543428 585920 543430
rect -1996 542826 -1396 542828
rect 585320 542826 585920 542828
rect 0 536596 584000 542508
rect -8576 536276 -7976 536278
rect 591900 536276 592500 536278
rect -8576 535674 -7976 535676
rect 591900 535674 592500 535676
rect 0 532996 584000 535356
rect -6696 532676 -6096 532678
rect 590020 532676 590620 532678
rect -6696 532074 -6096 532076
rect 590020 532074 590620 532076
rect 0 529396 584000 531756
rect -4816 529076 -4216 529078
rect 588140 529076 588740 529078
rect -4816 528474 -4216 528476
rect 588140 528474 588740 528476
rect 0 525748 584000 528156
rect -2936 525428 -2336 525430
rect 586260 525428 586860 525430
rect -2936 524826 -2336 524828
rect 586260 524826 586860 524828
rect 0 518596 584000 524508
rect -7636 518276 -7036 518278
rect 590960 518276 591560 518278
rect -7636 517674 -7036 517676
rect 590960 517674 591560 517676
rect 0 514996 584000 517356
rect -5756 514676 -5156 514678
rect 589080 514676 589680 514678
rect -5756 514074 -5156 514076
rect 589080 514074 589680 514076
rect 0 511396 584000 513756
rect -3876 511076 -3276 511078
rect 587200 511076 587800 511078
rect -3876 510474 -3276 510476
rect 587200 510474 587800 510476
rect 0 507748 584000 510156
rect -1996 507428 -1396 507430
rect 585320 507428 585920 507430
rect -1996 506826 -1396 506828
rect 585320 506826 585920 506828
rect 0 500596 584000 506508
rect -8576 500276 -7976 500278
rect 591900 500276 592500 500278
rect -8576 499674 -7976 499676
rect 591900 499674 592500 499676
rect 0 496996 584000 499356
rect -6696 496676 -6096 496678
rect 590020 496676 590620 496678
rect -6696 496074 -6096 496076
rect 590020 496074 590620 496076
rect 0 493396 584000 495756
rect -4816 493076 -4216 493078
rect 588140 493076 588740 493078
rect -4816 492474 -4216 492476
rect 588140 492474 588740 492476
rect 0 489748 584000 492156
rect -2936 489428 -2336 489430
rect 586260 489428 586860 489430
rect -2936 488826 -2336 488828
rect 586260 488826 586860 488828
rect 0 482596 584000 488508
rect -7636 482276 -7036 482278
rect 590960 482276 591560 482278
rect -7636 481674 -7036 481676
rect 590960 481674 591560 481676
rect 0 478996 584000 481356
rect -5756 478676 -5156 478678
rect 589080 478676 589680 478678
rect -5756 478074 -5156 478076
rect 589080 478074 589680 478076
rect 0 475396 584000 477756
rect -3876 475076 -3276 475078
rect 587200 475076 587800 475078
rect -3876 474474 -3276 474476
rect 587200 474474 587800 474476
rect 0 471748 584000 474156
rect -1996 471428 -1396 471430
rect 585320 471428 585920 471430
rect -1996 470826 -1396 470828
rect 585320 470826 585920 470828
rect 0 464596 584000 470508
rect -8576 464276 -7976 464278
rect 591900 464276 592500 464278
rect -8576 463674 -7976 463676
rect 591900 463674 592500 463676
rect 0 460996 584000 463356
rect -6696 460676 -6096 460678
rect 590020 460676 590620 460678
rect -6696 460074 -6096 460076
rect 590020 460074 590620 460076
rect 0 457396 584000 459756
rect -4816 457076 -4216 457078
rect 588140 457076 588740 457078
rect -4816 456474 -4216 456476
rect 588140 456474 588740 456476
rect 0 453748 584000 456156
rect -2936 453428 -2336 453430
rect 586260 453428 586860 453430
rect -2936 452826 -2336 452828
rect 586260 452826 586860 452828
rect 0 446596 584000 452508
rect -7636 446276 -7036 446278
rect 590960 446276 591560 446278
rect -7636 445674 -7036 445676
rect 590960 445674 591560 445676
rect 0 442996 584000 445356
rect -5756 442676 -5156 442678
rect 589080 442676 589680 442678
rect -5756 442074 -5156 442076
rect 589080 442074 589680 442076
rect 0 439396 584000 441756
rect -3876 439076 -3276 439078
rect 587200 439076 587800 439078
rect -3876 438474 -3276 438476
rect 587200 438474 587800 438476
rect 0 435748 584000 438156
rect -1996 435428 -1396 435430
rect 585320 435428 585920 435430
rect -1996 434826 -1396 434828
rect 585320 434826 585920 434828
rect 0 428596 584000 434508
rect -8576 428276 -7976 428278
rect 591900 428276 592500 428278
rect -8576 427674 -7976 427676
rect 591900 427674 592500 427676
rect 0 424996 584000 427356
rect -6696 424676 -6096 424678
rect 590020 424676 590620 424678
rect -6696 424074 -6096 424076
rect 590020 424074 590620 424076
rect 0 421396 584000 423756
rect -4816 421076 -4216 421078
rect 588140 421076 588740 421078
rect -4816 420474 -4216 420476
rect 588140 420474 588740 420476
rect 0 417748 584000 420156
rect -2936 417428 -2336 417430
rect 586260 417428 586860 417430
rect -2936 416826 -2336 416828
rect 586260 416826 586860 416828
rect 0 410596 584000 416508
rect -7636 410276 -7036 410278
rect 590960 410276 591560 410278
rect -7636 409674 -7036 409676
rect 590960 409674 591560 409676
rect 0 406996 584000 409356
rect -5756 406676 -5156 406678
rect 589080 406676 589680 406678
rect -5756 406074 -5156 406076
rect 589080 406074 589680 406076
rect 0 403396 584000 405756
rect -3876 403076 -3276 403078
rect 587200 403076 587800 403078
rect -3876 402474 -3276 402476
rect 587200 402474 587800 402476
rect 0 399748 584000 402156
rect -1996 399428 -1396 399430
rect 585320 399428 585920 399430
rect -1996 398826 -1396 398828
rect 585320 398826 585920 398828
rect 0 392596 584000 398508
rect -8576 392276 -7976 392278
rect 591900 392276 592500 392278
rect -8576 391674 -7976 391676
rect 591900 391674 592500 391676
rect 0 388996 584000 391356
rect -6696 388676 -6096 388678
rect 590020 388676 590620 388678
rect -6696 388074 -6096 388076
rect 590020 388074 590620 388076
rect 0 385396 584000 387756
rect -4816 385076 -4216 385078
rect 588140 385076 588740 385078
rect -4816 384474 -4216 384476
rect 588140 384474 588740 384476
rect 0 381748 584000 384156
rect -2936 381428 -2336 381430
rect 586260 381428 586860 381430
rect -2936 380826 -2336 380828
rect 586260 380826 586860 380828
rect 0 374596 584000 380508
rect -7636 374276 -7036 374278
rect 590960 374276 591560 374278
rect -7636 373674 -7036 373676
rect 590960 373674 591560 373676
rect 0 370996 584000 373356
rect -5756 370676 -5156 370678
rect 589080 370676 589680 370678
rect -5756 370074 -5156 370076
rect 589080 370074 589680 370076
rect 0 367396 584000 369756
rect -3876 367076 -3276 367078
rect 587200 367076 587800 367078
rect -3876 366474 -3276 366476
rect 587200 366474 587800 366476
rect 0 363748 584000 366156
rect -1996 363428 -1396 363430
rect 585320 363428 585920 363430
rect -1996 362826 -1396 362828
rect 585320 362826 585920 362828
rect 0 356596 584000 362508
rect -8576 356276 -7976 356278
rect 591900 356276 592500 356278
rect -8576 355674 -7976 355676
rect 591900 355674 592500 355676
rect 0 352996 584000 355356
rect -6696 352676 -6096 352678
rect 590020 352676 590620 352678
rect -6696 352074 -6096 352076
rect 590020 352074 590620 352076
rect 0 349396 584000 351756
rect -4816 349076 -4216 349078
rect 588140 349076 588740 349078
rect -4816 348474 -4216 348476
rect 588140 348474 588740 348476
rect 0 345748 584000 348156
rect -2936 345428 -2336 345430
rect 586260 345428 586860 345430
rect -2936 344826 -2336 344828
rect 586260 344826 586860 344828
rect 0 338596 584000 344508
rect -7636 338276 -7036 338278
rect 590960 338276 591560 338278
rect -7636 337674 -7036 337676
rect 590960 337674 591560 337676
rect 0 334996 584000 337356
rect -5756 334676 -5156 334678
rect 589080 334676 589680 334678
rect -5756 334074 -5156 334076
rect 589080 334074 589680 334076
rect 0 331396 584000 333756
rect -3876 331076 -3276 331078
rect 587200 331076 587800 331078
rect -3876 330474 -3276 330476
rect 587200 330474 587800 330476
rect 0 327748 584000 330156
rect -1996 327428 -1396 327430
rect 585320 327428 585920 327430
rect -1996 326826 -1396 326828
rect 585320 326826 585920 326828
rect 0 320596 584000 326508
rect -8576 320276 -7976 320278
rect 591900 320276 592500 320278
rect -8576 319674 -7976 319676
rect 591900 319674 592500 319676
rect 0 316996 584000 319356
rect -6696 316676 -6096 316678
rect 590020 316676 590620 316678
rect -6696 316074 -6096 316076
rect 590020 316074 590620 316076
rect 0 313396 584000 315756
rect -4816 313076 -4216 313078
rect 588140 313076 588740 313078
rect -4816 312474 -4216 312476
rect 588140 312474 588740 312476
rect 0 309748 584000 312156
rect -2936 309428 -2336 309430
rect 586260 309428 586860 309430
rect -2936 308826 -2336 308828
rect 586260 308826 586860 308828
rect 0 302596 584000 308508
rect -7636 302276 -7036 302278
rect 590960 302276 591560 302278
rect -7636 301674 -7036 301676
rect 590960 301674 591560 301676
rect 0 298996 584000 301356
rect -5756 298676 -5156 298678
rect 589080 298676 589680 298678
rect -5756 298074 -5156 298076
rect 589080 298074 589680 298076
rect 0 295396 584000 297756
rect -3876 295076 -3276 295078
rect 587200 295076 587800 295078
rect -3876 294474 -3276 294476
rect 587200 294474 587800 294476
rect 0 291748 584000 294156
rect -1996 291428 -1396 291430
rect 585320 291428 585920 291430
rect -1996 290826 -1396 290828
rect 585320 290826 585920 290828
rect 0 284596 584000 290508
rect -8576 284276 -7976 284278
rect 591900 284276 592500 284278
rect -8576 283674 -7976 283676
rect 591900 283674 592500 283676
rect 0 280996 584000 283356
rect -6696 280676 -6096 280678
rect 590020 280676 590620 280678
rect -6696 280074 -6096 280076
rect 590020 280074 590620 280076
rect 0 277396 584000 279756
rect -4816 277076 -4216 277078
rect 588140 277076 588740 277078
rect -4816 276474 -4216 276476
rect 588140 276474 588740 276476
rect 0 273748 584000 276156
rect -2936 273428 -2336 273430
rect 586260 273428 586860 273430
rect -2936 272826 -2336 272828
rect 586260 272826 586860 272828
rect 0 266596 584000 272508
rect -7636 266276 -7036 266278
rect 590960 266276 591560 266278
rect -7636 265674 -7036 265676
rect 590960 265674 591560 265676
rect 0 262996 584000 265356
rect -5756 262676 -5156 262678
rect 589080 262676 589680 262678
rect -5756 262074 -5156 262076
rect 589080 262074 589680 262076
rect 0 259396 584000 261756
rect -3876 259076 -3276 259078
rect 587200 259076 587800 259078
rect -3876 258474 -3276 258476
rect 587200 258474 587800 258476
rect 0 255748 584000 258156
rect -1996 255428 -1396 255430
rect 585320 255428 585920 255430
rect -1996 254826 -1396 254828
rect 585320 254826 585920 254828
rect 0 248596 584000 254508
rect -8576 248276 -7976 248278
rect 591900 248276 592500 248278
rect -8576 247674 -7976 247676
rect 591900 247674 592500 247676
rect 0 244996 584000 247356
rect -6696 244676 -6096 244678
rect 590020 244676 590620 244678
rect -6696 244074 -6096 244076
rect 590020 244074 590620 244076
rect 0 241396 584000 243756
rect -4816 241076 -4216 241078
rect 588140 241076 588740 241078
rect -4816 240474 -4216 240476
rect 588140 240474 588740 240476
rect 0 237748 584000 240156
rect -2936 237428 -2336 237430
rect 586260 237428 586860 237430
rect -2936 236826 -2336 236828
rect 586260 236826 586860 236828
rect 0 230596 584000 236508
rect -7636 230276 -7036 230278
rect 590960 230276 591560 230278
rect -7636 229674 -7036 229676
rect 590960 229674 591560 229676
rect 0 226996 584000 229356
rect -5756 226676 -5156 226678
rect 589080 226676 589680 226678
rect -5756 226074 -5156 226076
rect 589080 226074 589680 226076
rect 0 223396 584000 225756
rect -3876 223076 -3276 223078
rect 587200 223076 587800 223078
rect -3876 222474 -3276 222476
rect 587200 222474 587800 222476
rect 0 219748 584000 222156
rect -1996 219428 -1396 219430
rect 585320 219428 585920 219430
rect -1996 218826 -1396 218828
rect 585320 218826 585920 218828
rect 0 212596 584000 218508
rect -8576 212276 -7976 212278
rect 591900 212276 592500 212278
rect -8576 211674 -7976 211676
rect 591900 211674 592500 211676
rect 0 208996 584000 211356
rect -6696 208676 -6096 208678
rect 590020 208676 590620 208678
rect -6696 208074 -6096 208076
rect 590020 208074 590620 208076
rect 0 205396 584000 207756
rect -4816 205076 -4216 205078
rect 588140 205076 588740 205078
rect -4816 204474 -4216 204476
rect 588140 204474 588740 204476
rect 0 201748 584000 204156
rect -2936 201428 -2336 201430
rect 586260 201428 586860 201430
rect -2936 200826 -2336 200828
rect 586260 200826 586860 200828
rect 0 194596 584000 200508
rect -7636 194276 -7036 194278
rect 590960 194276 591560 194278
rect -7636 193674 -7036 193676
rect 590960 193674 591560 193676
rect 0 190996 584000 193356
rect -5756 190676 -5156 190678
rect 589080 190676 589680 190678
rect -5756 190074 -5156 190076
rect 589080 190074 589680 190076
rect 0 187396 584000 189756
rect -3876 187076 -3276 187078
rect 587200 187076 587800 187078
rect -3876 186474 -3276 186476
rect 587200 186474 587800 186476
rect 0 183748 584000 186156
rect -1996 183428 -1396 183430
rect 585320 183428 585920 183430
rect -1996 182826 -1396 182828
rect 585320 182826 585920 182828
rect 0 176596 584000 182508
rect -8576 176276 -7976 176278
rect 591900 176276 592500 176278
rect -8576 175674 -7976 175676
rect 591900 175674 592500 175676
rect 0 172996 584000 175356
rect -6696 172676 -6096 172678
rect 590020 172676 590620 172678
rect -6696 172074 -6096 172076
rect 590020 172074 590620 172076
rect 0 169396 584000 171756
rect -4816 169076 -4216 169078
rect 588140 169076 588740 169078
rect -4816 168474 -4216 168476
rect 588140 168474 588740 168476
rect 0 165748 584000 168156
rect -2936 165428 -2336 165430
rect 586260 165428 586860 165430
rect -2936 164826 -2336 164828
rect 586260 164826 586860 164828
rect 0 158596 584000 164508
rect -7636 158276 -7036 158278
rect 590960 158276 591560 158278
rect -7636 157674 -7036 157676
rect 590960 157674 591560 157676
rect 0 154996 584000 157356
rect -5756 154676 -5156 154678
rect 589080 154676 589680 154678
rect -5756 154074 -5156 154076
rect 589080 154074 589680 154076
rect 0 151396 584000 153756
rect -3876 151076 -3276 151078
rect 587200 151076 587800 151078
rect -3876 150474 -3276 150476
rect 587200 150474 587800 150476
rect 0 147748 584000 150156
rect -1996 147428 -1396 147430
rect 585320 147428 585920 147430
rect -1996 146826 -1396 146828
rect 585320 146826 585920 146828
rect 0 140596 584000 146508
rect -8576 140276 -7976 140278
rect 591900 140276 592500 140278
rect -8576 139674 -7976 139676
rect 591900 139674 592500 139676
rect 0 136996 584000 139356
rect -6696 136676 -6096 136678
rect 590020 136676 590620 136678
rect -6696 136074 -6096 136076
rect 590020 136074 590620 136076
rect 0 133396 584000 135756
rect -4816 133076 -4216 133078
rect 588140 133076 588740 133078
rect -4816 132474 -4216 132476
rect 588140 132474 588740 132476
rect 0 129748 584000 132156
rect -2936 129428 -2336 129430
rect 586260 129428 586860 129430
rect -2936 128826 -2336 128828
rect 586260 128826 586860 128828
rect 0 122596 584000 128508
rect -7636 122276 -7036 122278
rect 590960 122276 591560 122278
rect -7636 121674 -7036 121676
rect 590960 121674 591560 121676
rect 0 118996 584000 121356
rect -5756 118676 -5156 118678
rect 589080 118676 589680 118678
rect -5756 118074 -5156 118076
rect 589080 118074 589680 118076
rect 0 115396 584000 117756
rect -3876 115076 -3276 115078
rect 587200 115076 587800 115078
rect -3876 114474 -3276 114476
rect 587200 114474 587800 114476
rect 0 111748 584000 114156
rect -1996 111428 -1396 111430
rect 585320 111428 585920 111430
rect -1996 110826 -1396 110828
rect 585320 110826 585920 110828
rect 0 104596 584000 110508
rect -8576 104276 -7976 104278
rect 591900 104276 592500 104278
rect -8576 103674 -7976 103676
rect 591900 103674 592500 103676
rect 0 100996 584000 103356
rect -6696 100676 -6096 100678
rect 590020 100676 590620 100678
rect -6696 100074 -6096 100076
rect 590020 100074 590620 100076
rect 0 97396 584000 99756
rect -4816 97076 -4216 97078
rect 588140 97076 588740 97078
rect -4816 96474 -4216 96476
rect 588140 96474 588740 96476
rect 0 93748 584000 96156
rect -2936 93428 -2336 93430
rect 586260 93428 586860 93430
rect -2936 92826 -2336 92828
rect 586260 92826 586860 92828
rect 0 86596 584000 92508
rect -7636 86276 -7036 86278
rect 590960 86276 591560 86278
rect -7636 85674 -7036 85676
rect 590960 85674 591560 85676
rect 0 82996 584000 85356
rect -5756 82676 -5156 82678
rect 589080 82676 589680 82678
rect -5756 82074 -5156 82076
rect 589080 82074 589680 82076
rect 0 79396 584000 81756
rect -3876 79076 -3276 79078
rect 587200 79076 587800 79078
rect -3876 78474 -3276 78476
rect 587200 78474 587800 78476
rect 0 75748 584000 78156
rect -1996 75428 -1396 75430
rect 585320 75428 585920 75430
rect -1996 74826 -1396 74828
rect 585320 74826 585920 74828
rect 0 68596 584000 74508
rect -8576 68276 -7976 68278
rect 591900 68276 592500 68278
rect -8576 67674 -7976 67676
rect 591900 67674 592500 67676
rect 0 64996 584000 67356
rect -6696 64676 -6096 64678
rect 590020 64676 590620 64678
rect -6696 64074 -6096 64076
rect 590020 64074 590620 64076
rect 0 61396 584000 63756
rect -4816 61076 -4216 61078
rect 588140 61076 588740 61078
rect -4816 60474 -4216 60476
rect 588140 60474 588740 60476
rect 0 57748 584000 60156
rect -2936 57428 -2336 57430
rect 586260 57428 586860 57430
rect -2936 56826 -2336 56828
rect 586260 56826 586860 56828
rect 0 50596 584000 56508
rect -7636 50276 -7036 50278
rect 590960 50276 591560 50278
rect -7636 49674 -7036 49676
rect 590960 49674 591560 49676
rect 0 46996 584000 49356
rect -5756 46676 -5156 46678
rect 589080 46676 589680 46678
rect -5756 46074 -5156 46076
rect 589080 46074 589680 46076
rect 0 43396 584000 45756
rect -3876 43076 -3276 43078
rect 587200 43076 587800 43078
rect -3876 42474 -3276 42476
rect 587200 42474 587800 42476
rect 0 39748 584000 42156
rect -1996 39428 -1396 39430
rect 585320 39428 585920 39430
rect -1996 38826 -1396 38828
rect 585320 38826 585920 38828
rect 0 32596 584000 38508
rect -8576 32276 -7976 32278
rect 591900 32276 592500 32278
rect -8576 31674 -7976 31676
rect 591900 31674 592500 31676
rect 0 28996 584000 31356
rect -6696 28676 -6096 28678
rect 590020 28676 590620 28678
rect -6696 28074 -6096 28076
rect 590020 28074 590620 28076
rect 0 25396 584000 27756
rect -4816 25076 -4216 25078
rect 588140 25076 588740 25078
rect -4816 24474 -4216 24476
rect 588140 24474 588740 24476
rect 0 21748 584000 24156
rect -2936 21428 -2336 21430
rect 586260 21428 586860 21430
rect -2936 20826 -2336 20828
rect 586260 20826 586860 20828
rect 0 14596 584000 20508
rect -7636 14276 -7036 14278
rect 590960 14276 591560 14278
rect -7636 13674 -7036 13676
rect 590960 13674 591560 13676
rect 0 10996 584000 13356
rect -5756 10676 -5156 10678
rect 589080 10676 589680 10678
rect -5756 10074 -5156 10076
rect 589080 10074 589680 10076
rect 0 7396 584000 9756
rect -3876 7076 -3276 7078
rect 587200 7076 587800 7078
rect -3876 6474 -3276 6476
rect 587200 6474 587800 6476
rect 0 3748 584000 6156
rect -1996 3428 -1396 3430
rect 585320 3428 585920 3430
rect -1996 2826 -1396 2828
rect 585320 2826 585920 2828
rect 0 0 584000 2508
rect -1996 -324 -1396 -322
rect 1804 -324 2404 -322
rect 37804 -324 38404 -322
rect 73804 -324 74404 -322
rect 109804 -324 110404 -322
rect 145804 -324 146404 -322
rect 181804 -324 182404 -322
rect 217804 -324 218404 -322
rect 253804 -324 254404 -322
rect 289804 -324 290404 -322
rect 325804 -324 326404 -322
rect 361804 -324 362404 -322
rect 397804 -324 398404 -322
rect 433804 -324 434404 -322
rect 469804 -324 470404 -322
rect 505804 -324 506404 -322
rect 541804 -324 542404 -322
rect 577804 -324 578404 -322
rect 585320 -324 585920 -322
rect -1996 -926 -1396 -924
rect 1804 -926 2404 -924
rect 37804 -926 38404 -924
rect 73804 -926 74404 -924
rect 109804 -926 110404 -924
rect 145804 -926 146404 -924
rect 181804 -926 182404 -924
rect 217804 -926 218404 -924
rect 253804 -926 254404 -924
rect 289804 -926 290404 -924
rect 325804 -926 326404 -924
rect 361804 -926 362404 -924
rect 397804 -926 398404 -924
rect 433804 -926 434404 -924
rect 469804 -926 470404 -924
rect 505804 -926 506404 -924
rect 541804 -926 542404 -924
rect 577804 -926 578404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 19804 -1264 20404 -1262
rect 55804 -1264 56404 -1262
rect 91804 -1264 92404 -1262
rect 127804 -1264 128404 -1262
rect 163804 -1264 164404 -1262
rect 199804 -1264 200404 -1262
rect 235804 -1264 236404 -1262
rect 271804 -1264 272404 -1262
rect 307804 -1264 308404 -1262
rect 343804 -1264 344404 -1262
rect 379804 -1264 380404 -1262
rect 415804 -1264 416404 -1262
rect 451804 -1264 452404 -1262
rect 487804 -1264 488404 -1262
rect 523804 -1264 524404 -1262
rect 559804 -1264 560404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1866 -2336 -1864
rect 19804 -1866 20404 -1864
rect 55804 -1866 56404 -1864
rect 91804 -1866 92404 -1864
rect 127804 -1866 128404 -1864
rect 163804 -1866 164404 -1864
rect 199804 -1866 200404 -1864
rect 235804 -1866 236404 -1864
rect 271804 -1866 272404 -1864
rect 307804 -1866 308404 -1864
rect 343804 -1866 344404 -1864
rect 379804 -1866 380404 -1864
rect 415804 -1866 416404 -1864
rect 451804 -1866 452404 -1864
rect 487804 -1866 488404 -1864
rect 523804 -1866 524404 -1864
rect 559804 -1866 560404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 5404 -2204 6004 -2202
rect 41404 -2204 42004 -2202
rect 77404 -2204 78004 -2202
rect 113404 -2204 114004 -2202
rect 149404 -2204 150004 -2202
rect 185404 -2204 186004 -2202
rect 221404 -2204 222004 -2202
rect 257404 -2204 258004 -2202
rect 293404 -2204 294004 -2202
rect 329404 -2204 330004 -2202
rect 365404 -2204 366004 -2202
rect 401404 -2204 402004 -2202
rect 437404 -2204 438004 -2202
rect 473404 -2204 474004 -2202
rect 509404 -2204 510004 -2202
rect 545404 -2204 546004 -2202
rect 581404 -2204 582004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2806 -3276 -2804
rect 5404 -2806 6004 -2804
rect 41404 -2806 42004 -2804
rect 77404 -2806 78004 -2804
rect 113404 -2806 114004 -2804
rect 149404 -2806 150004 -2804
rect 185404 -2806 186004 -2804
rect 221404 -2806 222004 -2804
rect 257404 -2806 258004 -2804
rect 293404 -2806 294004 -2804
rect 329404 -2806 330004 -2804
rect 365404 -2806 366004 -2804
rect 401404 -2806 402004 -2804
rect 437404 -2806 438004 -2804
rect 473404 -2806 474004 -2804
rect 509404 -2806 510004 -2804
rect 545404 -2806 546004 -2804
rect 581404 -2806 582004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 23404 -3144 24004 -3142
rect 59404 -3144 60004 -3142
rect 95404 -3144 96004 -3142
rect 131404 -3144 132004 -3142
rect 167404 -3144 168004 -3142
rect 203404 -3144 204004 -3142
rect 239404 -3144 240004 -3142
rect 275404 -3144 276004 -3142
rect 311404 -3144 312004 -3142
rect 347404 -3144 348004 -3142
rect 383404 -3144 384004 -3142
rect 419404 -3144 420004 -3142
rect 455404 -3144 456004 -3142
rect 491404 -3144 492004 -3142
rect 527404 -3144 528004 -3142
rect 563404 -3144 564004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3746 -4216 -3744
rect 23404 -3746 24004 -3744
rect 59404 -3746 60004 -3744
rect 95404 -3746 96004 -3744
rect 131404 -3746 132004 -3744
rect 167404 -3746 168004 -3744
rect 203404 -3746 204004 -3744
rect 239404 -3746 240004 -3744
rect 275404 -3746 276004 -3744
rect 311404 -3746 312004 -3744
rect 347404 -3746 348004 -3744
rect 383404 -3746 384004 -3744
rect 419404 -3746 420004 -3744
rect 455404 -3746 456004 -3744
rect 491404 -3746 492004 -3744
rect 527404 -3746 528004 -3744
rect 563404 -3746 564004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 9004 -4084 9604 -4082
rect 45004 -4084 45604 -4082
rect 81004 -4084 81604 -4082
rect 117004 -4084 117604 -4082
rect 153004 -4084 153604 -4082
rect 189004 -4084 189604 -4082
rect 225004 -4084 225604 -4082
rect 261004 -4084 261604 -4082
rect 297004 -4084 297604 -4082
rect 333004 -4084 333604 -4082
rect 369004 -4084 369604 -4082
rect 405004 -4084 405604 -4082
rect 441004 -4084 441604 -4082
rect 477004 -4084 477604 -4082
rect 513004 -4084 513604 -4082
rect 549004 -4084 549604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4686 -5156 -4684
rect 9004 -4686 9604 -4684
rect 45004 -4686 45604 -4684
rect 81004 -4686 81604 -4684
rect 117004 -4686 117604 -4684
rect 153004 -4686 153604 -4684
rect 189004 -4686 189604 -4684
rect 225004 -4686 225604 -4684
rect 261004 -4686 261604 -4684
rect 297004 -4686 297604 -4684
rect 333004 -4686 333604 -4684
rect 369004 -4686 369604 -4684
rect 405004 -4686 405604 -4684
rect 441004 -4686 441604 -4684
rect 477004 -4686 477604 -4684
rect 513004 -4686 513604 -4684
rect 549004 -4686 549604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 27004 -5024 27604 -5022
rect 63004 -5024 63604 -5022
rect 99004 -5024 99604 -5022
rect 135004 -5024 135604 -5022
rect 171004 -5024 171604 -5022
rect 207004 -5024 207604 -5022
rect 243004 -5024 243604 -5022
rect 279004 -5024 279604 -5022
rect 315004 -5024 315604 -5022
rect 351004 -5024 351604 -5022
rect 387004 -5024 387604 -5022
rect 423004 -5024 423604 -5022
rect 459004 -5024 459604 -5022
rect 495004 -5024 495604 -5022
rect 531004 -5024 531604 -5022
rect 567004 -5024 567604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5626 -6096 -5624
rect 27004 -5626 27604 -5624
rect 63004 -5626 63604 -5624
rect 99004 -5626 99604 -5624
rect 135004 -5626 135604 -5624
rect 171004 -5626 171604 -5624
rect 207004 -5626 207604 -5624
rect 243004 -5626 243604 -5624
rect 279004 -5626 279604 -5624
rect 315004 -5626 315604 -5624
rect 351004 -5626 351604 -5624
rect 387004 -5626 387604 -5624
rect 423004 -5626 423604 -5624
rect 459004 -5626 459604 -5624
rect 495004 -5626 495604 -5624
rect 531004 -5626 531604 -5624
rect 567004 -5626 567604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 12604 -5964 13204 -5962
rect 48604 -5964 49204 -5962
rect 84604 -5964 85204 -5962
rect 120604 -5964 121204 -5962
rect 156604 -5964 157204 -5962
rect 192604 -5964 193204 -5962
rect 228604 -5964 229204 -5962
rect 264604 -5964 265204 -5962
rect 300604 -5964 301204 -5962
rect 336604 -5964 337204 -5962
rect 372604 -5964 373204 -5962
rect 408604 -5964 409204 -5962
rect 444604 -5964 445204 -5962
rect 480604 -5964 481204 -5962
rect 516604 -5964 517204 -5962
rect 552604 -5964 553204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -6566 -7036 -6564
rect 12604 -6566 13204 -6564
rect 48604 -6566 49204 -6564
rect 84604 -6566 85204 -6564
rect 120604 -6566 121204 -6564
rect 156604 -6566 157204 -6564
rect 192604 -6566 193204 -6564
rect 228604 -6566 229204 -6564
rect 264604 -6566 265204 -6564
rect 300604 -6566 301204 -6564
rect 336604 -6566 337204 -6564
rect 372604 -6566 373204 -6564
rect 408604 -6566 409204 -6564
rect 444604 -6566 445204 -6564
rect 480604 -6566 481204 -6564
rect 516604 -6566 517204 -6564
rect 552604 -6566 553204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 30604 -6904 31204 -6902
rect 66604 -6904 67204 -6902
rect 102604 -6904 103204 -6902
rect 138604 -6904 139204 -6902
rect 174604 -6904 175204 -6902
rect 210604 -6904 211204 -6902
rect 246604 -6904 247204 -6902
rect 282604 -6904 283204 -6902
rect 318604 -6904 319204 -6902
rect 354604 -6904 355204 -6902
rect 390604 -6904 391204 -6902
rect 426604 -6904 427204 -6902
rect 462604 -6904 463204 -6902
rect 498604 -6904 499204 -6902
rect 534604 -6904 535204 -6902
rect 570604 -6904 571204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -7506 -7976 -7504
rect 30604 -7506 31204 -7504
rect 66604 -7506 67204 -7504
rect 102604 -7506 103204 -7504
rect 138604 -7506 139204 -7504
rect 174604 -7506 175204 -7504
rect 210604 -7506 211204 -7504
rect 246604 -7506 247204 -7504
rect 282604 -7506 283204 -7504
rect 318604 -7506 319204 -7504
rect 354604 -7506 355204 -7504
rect 390604 -7506 391204 -7504
rect 426604 -7506 427204 -7504
rect 462604 -7506 463204 -7504
rect 498604 -7506 499204 -7504
rect 534604 -7506 535204 -7504
rect 570604 -7506 571204 -7504
rect 591900 -7506 592500 -7504
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 532 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 533 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 534 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 535 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 536 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 537 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 538 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 539 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 540 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 541 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 542 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 543 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 544 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 545 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 546 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 547 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 548 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 549 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 550 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 551 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 552 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 553 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 554 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 555 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 556 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 557 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 558 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 559 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 560 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 561 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 562 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 563 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 564 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 565 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 566 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 567 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 568 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 569 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 570 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 571 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 572 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 573 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 574 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 575 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 576 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 577 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 578 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 579 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 580 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 581 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 582 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 583 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 584 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 585 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 586 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 587 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 588 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 589 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 590 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 591 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 592 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 593 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 594 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 595 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 596 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 597 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 598 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 599 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 600 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 601 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 602 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 603 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 604 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 605 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 606 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 607 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 608 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 609 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 610 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 611 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 612 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 613 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 614 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 615 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 616 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 617 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 618 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 619 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 620 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 621 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 622 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 623 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 624 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 625 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 626 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 627 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 628 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 629 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 630 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 631 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 632 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 633 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 634 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 635 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 636 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 637 nsew signal input
rlabel metal4 s 577804 -1864 578404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 541804 690352 542404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 505804 690352 506404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 469804 690352 470404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 433804 690352 434404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 397804 690352 398404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 361804 690352 362404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 325804 690352 326404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 289804 690352 290404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 253804 690352 254404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 217804 690352 218404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 181804 132152 182404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 145804 690352 146404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 109804 690352 110404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 73804 690352 74404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 37804 690352 38404 705800 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s 1804 -1864 2404 705800 6 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 541804 620992 542404 630448 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 505804 620992 506404 630448 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 469804 620992 470404 630448 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 433804 620992 434404 630448 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 397804 620992 398404 630448 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 361804 620992 362404 630448 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 325804 620992 326404 630448 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 289804 620992 290404 630448 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 253804 620992 254404 630448 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 217804 620992 218404 630448 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 145804 620992 146404 630448 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 109804 620992 110404 630448 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 73804 620992 74404 630448 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 37804 620992 38404 630448 6 vccd1
port 670 nsew power bidirectional
rlabel metal4 s 541804 551632 542404 561088 6 vccd1
port 671 nsew power bidirectional
rlabel metal4 s 505804 551632 506404 561088 6 vccd1
port 672 nsew power bidirectional
rlabel metal4 s 469804 551632 470404 561088 6 vccd1
port 673 nsew power bidirectional
rlabel metal4 s 433804 551632 434404 561088 6 vccd1
port 674 nsew power bidirectional
rlabel metal4 s 397804 551632 398404 561088 6 vccd1
port 675 nsew power bidirectional
rlabel metal4 s 361804 551632 362404 561088 6 vccd1
port 676 nsew power bidirectional
rlabel metal4 s 325804 551632 326404 561088 6 vccd1
port 677 nsew power bidirectional
rlabel metal4 s 289804 551632 290404 561088 6 vccd1
port 678 nsew power bidirectional
rlabel metal4 s 253804 551632 254404 561088 6 vccd1
port 679 nsew power bidirectional
rlabel metal4 s 217804 551632 218404 561088 6 vccd1
port 680 nsew power bidirectional
rlabel metal4 s 145804 551632 146404 561088 6 vccd1
port 681 nsew power bidirectional
rlabel metal4 s 109804 551632 110404 561088 6 vccd1
port 682 nsew power bidirectional
rlabel metal4 s 73804 551632 74404 561088 6 vccd1
port 683 nsew power bidirectional
rlabel metal4 s 37804 551632 38404 561088 6 vccd1
port 684 nsew power bidirectional
rlabel metal4 s 541804 482272 542404 491728 6 vccd1
port 685 nsew power bidirectional
rlabel metal4 s 505804 482272 506404 491728 6 vccd1
port 686 nsew power bidirectional
rlabel metal4 s 469804 482272 470404 491728 6 vccd1
port 687 nsew power bidirectional
rlabel metal4 s 433804 482272 434404 491728 6 vccd1
port 688 nsew power bidirectional
rlabel metal4 s 397804 482272 398404 491728 6 vccd1
port 689 nsew power bidirectional
rlabel metal4 s 361804 482272 362404 491728 6 vccd1
port 690 nsew power bidirectional
rlabel metal4 s 325804 482272 326404 491728 6 vccd1
port 691 nsew power bidirectional
rlabel metal4 s 289804 482272 290404 491728 6 vccd1
port 692 nsew power bidirectional
rlabel metal4 s 253804 482272 254404 491728 6 vccd1
port 693 nsew power bidirectional
rlabel metal4 s 217804 482272 218404 491728 6 vccd1
port 694 nsew power bidirectional
rlabel metal4 s 145804 482272 146404 491728 6 vccd1
port 695 nsew power bidirectional
rlabel metal4 s 109804 482272 110404 491728 6 vccd1
port 696 nsew power bidirectional
rlabel metal4 s 73804 482272 74404 491728 6 vccd1
port 697 nsew power bidirectional
rlabel metal4 s 37804 482272 38404 491728 6 vccd1
port 698 nsew power bidirectional
rlabel metal4 s 541804 412912 542404 422368 6 vccd1
port 699 nsew power bidirectional
rlabel metal4 s 505804 412912 506404 422368 6 vccd1
port 700 nsew power bidirectional
rlabel metal4 s 469804 412912 470404 422368 6 vccd1
port 701 nsew power bidirectional
rlabel metal4 s 433804 412912 434404 422368 6 vccd1
port 702 nsew power bidirectional
rlabel metal4 s 397804 412912 398404 422368 6 vccd1
port 703 nsew power bidirectional
rlabel metal4 s 361804 412912 362404 422368 6 vccd1
port 704 nsew power bidirectional
rlabel metal4 s 325804 412912 326404 422368 6 vccd1
port 705 nsew power bidirectional
rlabel metal4 s 289804 412912 290404 422368 6 vccd1
port 706 nsew power bidirectional
rlabel metal4 s 253804 412912 254404 422368 6 vccd1
port 707 nsew power bidirectional
rlabel metal4 s 217804 412912 218404 422368 6 vccd1
port 708 nsew power bidirectional
rlabel metal4 s 145804 412912 146404 422368 6 vccd1
port 709 nsew power bidirectional
rlabel metal4 s 109804 412912 110404 422368 6 vccd1
port 710 nsew power bidirectional
rlabel metal4 s 73804 412912 74404 422368 6 vccd1
port 711 nsew power bidirectional
rlabel metal4 s 37804 412912 38404 422368 6 vccd1
port 712 nsew power bidirectional
rlabel metal4 s 541804 343552 542404 353008 6 vccd1
port 713 nsew power bidirectional
rlabel metal4 s 505804 343552 506404 353008 6 vccd1
port 714 nsew power bidirectional
rlabel metal4 s 469804 343552 470404 353008 6 vccd1
port 715 nsew power bidirectional
rlabel metal4 s 433804 343552 434404 353008 6 vccd1
port 716 nsew power bidirectional
rlabel metal4 s 397804 343552 398404 353008 6 vccd1
port 717 nsew power bidirectional
rlabel metal4 s 361804 343552 362404 353008 6 vccd1
port 718 nsew power bidirectional
rlabel metal4 s 325804 343552 326404 353008 6 vccd1
port 719 nsew power bidirectional
rlabel metal4 s 289804 343552 290404 353008 6 vccd1
port 720 nsew power bidirectional
rlabel metal4 s 253804 343552 254404 353008 6 vccd1
port 721 nsew power bidirectional
rlabel metal4 s 217804 343552 218404 353008 6 vccd1
port 722 nsew power bidirectional
rlabel metal4 s 145804 343552 146404 353008 6 vccd1
port 723 nsew power bidirectional
rlabel metal4 s 109804 343552 110404 353008 6 vccd1
port 724 nsew power bidirectional
rlabel metal4 s 73804 343552 74404 353008 6 vccd1
port 725 nsew power bidirectional
rlabel metal4 s 37804 343552 38404 353008 6 vccd1
port 726 nsew power bidirectional
rlabel metal4 s 541804 274192 542404 283648 6 vccd1
port 727 nsew power bidirectional
rlabel metal4 s 505804 274192 506404 283648 6 vccd1
port 728 nsew power bidirectional
rlabel metal4 s 469804 274192 470404 283648 6 vccd1
port 729 nsew power bidirectional
rlabel metal4 s 433804 274192 434404 283648 6 vccd1
port 730 nsew power bidirectional
rlabel metal4 s 397804 274192 398404 283648 6 vccd1
port 731 nsew power bidirectional
rlabel metal4 s 361804 274192 362404 283648 6 vccd1
port 732 nsew power bidirectional
rlabel metal4 s 325804 274192 326404 283648 6 vccd1
port 733 nsew power bidirectional
rlabel metal4 s 289804 274192 290404 283648 6 vccd1
port 734 nsew power bidirectional
rlabel metal4 s 253804 274192 254404 283648 6 vccd1
port 735 nsew power bidirectional
rlabel metal4 s 217804 274192 218404 283648 6 vccd1
port 736 nsew power bidirectional
rlabel metal4 s 145804 274192 146404 283648 6 vccd1
port 737 nsew power bidirectional
rlabel metal4 s 109804 274192 110404 283648 6 vccd1
port 738 nsew power bidirectional
rlabel metal4 s 73804 274192 74404 283648 6 vccd1
port 739 nsew power bidirectional
rlabel metal4 s 37804 274192 38404 283648 6 vccd1
port 740 nsew power bidirectional
rlabel metal4 s 541804 204832 542404 214288 6 vccd1
port 741 nsew power bidirectional
rlabel metal4 s 505804 204832 506404 214288 6 vccd1
port 742 nsew power bidirectional
rlabel metal4 s 469804 204832 470404 214288 6 vccd1
port 743 nsew power bidirectional
rlabel metal4 s 433804 204832 434404 214288 6 vccd1
port 744 nsew power bidirectional
rlabel metal4 s 397804 204832 398404 214288 6 vccd1
port 745 nsew power bidirectional
rlabel metal4 s 361804 204832 362404 214288 6 vccd1
port 746 nsew power bidirectional
rlabel metal4 s 325804 204832 326404 214288 6 vccd1
port 747 nsew power bidirectional
rlabel metal4 s 289804 204832 290404 214288 6 vccd1
port 748 nsew power bidirectional
rlabel metal4 s 253804 204832 254404 214288 6 vccd1
port 749 nsew power bidirectional
rlabel metal4 s 217804 204832 218404 214288 6 vccd1
port 750 nsew power bidirectional
rlabel metal4 s 145804 204832 146404 214288 6 vccd1
port 751 nsew power bidirectional
rlabel metal4 s 109804 204832 110404 214288 6 vccd1
port 752 nsew power bidirectional
rlabel metal4 s 73804 204832 74404 214288 6 vccd1
port 753 nsew power bidirectional
rlabel metal4 s 37804 204832 38404 214288 6 vccd1
port 754 nsew power bidirectional
rlabel metal4 s 541804 132152 542404 144928 6 vccd1
port 755 nsew power bidirectional
rlabel metal4 s 505804 132152 506404 144928 6 vccd1
port 756 nsew power bidirectional
rlabel metal4 s 469804 132152 470404 144928 6 vccd1
port 757 nsew power bidirectional
rlabel metal4 s 433804 132152 434404 144928 6 vccd1
port 758 nsew power bidirectional
rlabel metal4 s 397804 132152 398404 144928 6 vccd1
port 759 nsew power bidirectional
rlabel metal4 s 361804 132152 362404 144928 6 vccd1
port 760 nsew power bidirectional
rlabel metal4 s 325804 132152 326404 144928 6 vccd1
port 761 nsew power bidirectional
rlabel metal4 s 289804 132152 290404 144928 6 vccd1
port 762 nsew power bidirectional
rlabel metal4 s 253804 132152 254404 144928 6 vccd1
port 763 nsew power bidirectional
rlabel metal4 s 217804 132152 218404 144928 6 vccd1
port 764 nsew power bidirectional
rlabel metal4 s 145804 132152 146404 144928 6 vccd1
port 765 nsew power bidirectional
rlabel metal4 s 109804 132152 110404 144928 6 vccd1
port 766 nsew power bidirectional
rlabel metal4 s 73804 132152 74404 144928 6 vccd1
port 767 nsew power bidirectional
rlabel metal4 s 37804 132152 38404 144928 6 vccd1
port 768 nsew power bidirectional
rlabel metal4 s 541804 -1864 542404 8248 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 505804 -1864 506404 8248 6 vccd1
port 770 nsew power bidirectional
rlabel metal4 s 469804 -1864 470404 8248 6 vccd1
port 771 nsew power bidirectional
rlabel metal4 s 433804 -1864 434404 8248 6 vccd1
port 772 nsew power bidirectional
rlabel metal4 s 397804 -1864 398404 8248 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 361804 -1864 362404 8248 6 vccd1
port 774 nsew power bidirectional
rlabel metal4 s 325804 -1864 326404 8248 6 vccd1
port 775 nsew power bidirectional
rlabel metal4 s 289804 -1864 290404 8248 6 vccd1
port 776 nsew power bidirectional
rlabel metal4 s 253804 -1864 254404 8248 6 vccd1
port 777 nsew power bidirectional
rlabel metal4 s 217804 -1864 218404 8248 6 vccd1
port 778 nsew power bidirectional
rlabel metal4 s 181804 -1864 182404 8248 6 vccd1
port 779 nsew power bidirectional
rlabel metal4 s 145804 -1864 146404 8248 6 vccd1
port 780 nsew power bidirectional
rlabel metal4 s 109804 -1864 110404 8248 6 vccd1
port 781 nsew power bidirectional
rlabel metal4 s 73804 -1864 74404 8248 6 vccd1
port 782 nsew power bidirectional
rlabel metal4 s 37804 -1864 38404 8248 6 vccd1
port 783 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 784 nsew power bidirectional
rlabel metal5 s -2936 686828 586860 687428 6 vccd1
port 785 nsew power bidirectional
rlabel metal5 s -2936 650828 586860 651428 6 vccd1
port 786 nsew power bidirectional
rlabel metal5 s -2936 614828 586860 615428 6 vccd1
port 787 nsew power bidirectional
rlabel metal5 s -2936 578828 586860 579428 6 vccd1
port 788 nsew power bidirectional
rlabel metal5 s -2936 542828 586860 543428 6 vccd1
port 789 nsew power bidirectional
rlabel metal5 s -2936 506828 586860 507428 6 vccd1
port 790 nsew power bidirectional
rlabel metal5 s -2936 470828 586860 471428 6 vccd1
port 791 nsew power bidirectional
rlabel metal5 s -2936 434828 586860 435428 6 vccd1
port 792 nsew power bidirectional
rlabel metal5 s -2936 398828 586860 399428 6 vccd1
port 793 nsew power bidirectional
rlabel metal5 s -2936 362828 586860 363428 6 vccd1
port 794 nsew power bidirectional
rlabel metal5 s -2936 326828 586860 327428 6 vccd1
port 795 nsew power bidirectional
rlabel metal5 s -2936 290828 586860 291428 6 vccd1
port 796 nsew power bidirectional
rlabel metal5 s -2936 254828 586860 255428 6 vccd1
port 797 nsew power bidirectional
rlabel metal5 s -2936 218828 586860 219428 6 vccd1
port 798 nsew power bidirectional
rlabel metal5 s -2936 182828 586860 183428 6 vccd1
port 799 nsew power bidirectional
rlabel metal5 s -2936 146828 586860 147428 6 vccd1
port 800 nsew power bidirectional
rlabel metal5 s -2936 110828 586860 111428 6 vccd1
port 801 nsew power bidirectional
rlabel metal5 s -2936 74828 586860 75428 6 vccd1
port 802 nsew power bidirectional
rlabel metal5 s -2936 38828 586860 39428 6 vccd1
port 803 nsew power bidirectional
rlabel metal5 s -2936 2828 586860 3428 6 vccd1
port 804 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 559804 690352 560404 705800 6 vssd1
port 807 nsew ground bidirectional
rlabel metal4 s 523804 690352 524404 705800 6 vssd1
port 808 nsew ground bidirectional
rlabel metal4 s 487804 132152 488404 705800 6 vssd1
port 809 nsew ground bidirectional
rlabel metal4 s 451804 690352 452404 705800 6 vssd1
port 810 nsew ground bidirectional
rlabel metal4 s 415804 690352 416404 705800 6 vssd1
port 811 nsew ground bidirectional
rlabel metal4 s 379804 690352 380404 705800 6 vssd1
port 812 nsew ground bidirectional
rlabel metal4 s 343804 690352 344404 705800 6 vssd1
port 813 nsew ground bidirectional
rlabel metal4 s 307804 690352 308404 705800 6 vssd1
port 814 nsew ground bidirectional
rlabel metal4 s 271804 132152 272404 705800 6 vssd1
port 815 nsew ground bidirectional
rlabel metal4 s 235804 690352 236404 705800 6 vssd1
port 816 nsew ground bidirectional
rlabel metal4 s 199804 690352 200404 705800 6 vssd1
port 817 nsew ground bidirectional
rlabel metal4 s 163804 690352 164404 705800 6 vssd1
port 818 nsew ground bidirectional
rlabel metal4 s 127804 690352 128404 705800 6 vssd1
port 819 nsew ground bidirectional
rlabel metal4 s 91804 -1864 92404 705800 6 vssd1
port 820 nsew ground bidirectional
rlabel metal4 s 55804 690352 56404 705800 6 vssd1
port 821 nsew ground bidirectional
rlabel metal4 s 19804 690352 20404 705800 6 vssd1
port 822 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 823 nsew ground bidirectional
rlabel metal4 s 559804 620992 560404 630448 6 vssd1
port 824 nsew ground bidirectional
rlabel metal4 s 523804 620992 524404 630448 6 vssd1
port 825 nsew ground bidirectional
rlabel metal4 s 451804 620992 452404 630448 6 vssd1
port 826 nsew ground bidirectional
rlabel metal4 s 415804 620992 416404 630448 6 vssd1
port 827 nsew ground bidirectional
rlabel metal4 s 379804 620992 380404 630448 6 vssd1
port 828 nsew ground bidirectional
rlabel metal4 s 343804 620992 344404 630448 6 vssd1
port 829 nsew ground bidirectional
rlabel metal4 s 307804 620992 308404 630448 6 vssd1
port 830 nsew ground bidirectional
rlabel metal4 s 235804 620992 236404 630448 6 vssd1
port 831 nsew ground bidirectional
rlabel metal4 s 199804 620992 200404 630448 6 vssd1
port 832 nsew ground bidirectional
rlabel metal4 s 163804 620992 164404 630448 6 vssd1
port 833 nsew ground bidirectional
rlabel metal4 s 127804 620992 128404 630448 6 vssd1
port 834 nsew ground bidirectional
rlabel metal4 s 55804 620992 56404 630448 6 vssd1
port 835 nsew ground bidirectional
rlabel metal4 s 19804 620992 20404 630448 6 vssd1
port 836 nsew ground bidirectional
rlabel metal4 s 559804 551632 560404 561088 6 vssd1
port 837 nsew ground bidirectional
rlabel metal4 s 523804 551632 524404 561088 6 vssd1
port 838 nsew ground bidirectional
rlabel metal4 s 451804 551632 452404 561088 6 vssd1
port 839 nsew ground bidirectional
rlabel metal4 s 415804 551632 416404 561088 6 vssd1
port 840 nsew ground bidirectional
rlabel metal4 s 379804 551632 380404 561088 6 vssd1
port 841 nsew ground bidirectional
rlabel metal4 s 343804 551632 344404 561088 6 vssd1
port 842 nsew ground bidirectional
rlabel metal4 s 307804 551632 308404 561088 6 vssd1
port 843 nsew ground bidirectional
rlabel metal4 s 235804 551632 236404 561088 6 vssd1
port 844 nsew ground bidirectional
rlabel metal4 s 199804 551632 200404 561088 6 vssd1
port 845 nsew ground bidirectional
rlabel metal4 s 163804 551632 164404 561088 6 vssd1
port 846 nsew ground bidirectional
rlabel metal4 s 127804 551632 128404 561088 6 vssd1
port 847 nsew ground bidirectional
rlabel metal4 s 55804 551632 56404 561088 6 vssd1
port 848 nsew ground bidirectional
rlabel metal4 s 19804 551632 20404 561088 6 vssd1
port 849 nsew ground bidirectional
rlabel metal4 s 559804 482272 560404 491728 6 vssd1
port 850 nsew ground bidirectional
rlabel metal4 s 523804 482272 524404 491728 6 vssd1
port 851 nsew ground bidirectional
rlabel metal4 s 451804 482272 452404 491728 6 vssd1
port 852 nsew ground bidirectional
rlabel metal4 s 415804 482272 416404 491728 6 vssd1
port 853 nsew ground bidirectional
rlabel metal4 s 379804 482272 380404 491728 6 vssd1
port 854 nsew ground bidirectional
rlabel metal4 s 343804 482272 344404 491728 6 vssd1
port 855 nsew ground bidirectional
rlabel metal4 s 307804 482272 308404 491728 6 vssd1
port 856 nsew ground bidirectional
rlabel metal4 s 235804 482272 236404 491728 6 vssd1
port 857 nsew ground bidirectional
rlabel metal4 s 199804 482272 200404 491728 6 vssd1
port 858 nsew ground bidirectional
rlabel metal4 s 163804 482272 164404 491728 6 vssd1
port 859 nsew ground bidirectional
rlabel metal4 s 127804 482272 128404 491728 6 vssd1
port 860 nsew ground bidirectional
rlabel metal4 s 55804 482272 56404 491728 6 vssd1
port 861 nsew ground bidirectional
rlabel metal4 s 19804 482272 20404 491728 6 vssd1
port 862 nsew ground bidirectional
rlabel metal4 s 559804 412912 560404 422368 6 vssd1
port 863 nsew ground bidirectional
rlabel metal4 s 523804 412912 524404 422368 6 vssd1
port 864 nsew ground bidirectional
rlabel metal4 s 451804 412912 452404 422368 6 vssd1
port 865 nsew ground bidirectional
rlabel metal4 s 415804 412912 416404 422368 6 vssd1
port 866 nsew ground bidirectional
rlabel metal4 s 379804 412912 380404 422368 6 vssd1
port 867 nsew ground bidirectional
rlabel metal4 s 343804 412912 344404 422368 6 vssd1
port 868 nsew ground bidirectional
rlabel metal4 s 307804 412912 308404 422368 6 vssd1
port 869 nsew ground bidirectional
rlabel metal4 s 235804 412912 236404 422368 6 vssd1
port 870 nsew ground bidirectional
rlabel metal4 s 199804 412912 200404 422368 6 vssd1
port 871 nsew ground bidirectional
rlabel metal4 s 163804 412912 164404 422368 6 vssd1
port 872 nsew ground bidirectional
rlabel metal4 s 127804 412912 128404 422368 6 vssd1
port 873 nsew ground bidirectional
rlabel metal4 s 55804 412912 56404 422368 6 vssd1
port 874 nsew ground bidirectional
rlabel metal4 s 19804 412912 20404 422368 6 vssd1
port 875 nsew ground bidirectional
rlabel metal4 s 559804 343552 560404 353008 6 vssd1
port 876 nsew ground bidirectional
rlabel metal4 s 523804 343552 524404 353008 6 vssd1
port 877 nsew ground bidirectional
rlabel metal4 s 451804 343552 452404 353008 6 vssd1
port 878 nsew ground bidirectional
rlabel metal4 s 415804 343552 416404 353008 6 vssd1
port 879 nsew ground bidirectional
rlabel metal4 s 379804 343552 380404 353008 6 vssd1
port 880 nsew ground bidirectional
rlabel metal4 s 343804 343552 344404 353008 6 vssd1
port 881 nsew ground bidirectional
rlabel metal4 s 307804 343552 308404 353008 6 vssd1
port 882 nsew ground bidirectional
rlabel metal4 s 235804 343552 236404 353008 6 vssd1
port 883 nsew ground bidirectional
rlabel metal4 s 199804 343552 200404 353008 6 vssd1
port 884 nsew ground bidirectional
rlabel metal4 s 163804 343552 164404 353008 6 vssd1
port 885 nsew ground bidirectional
rlabel metal4 s 127804 343552 128404 353008 6 vssd1
port 886 nsew ground bidirectional
rlabel metal4 s 55804 343552 56404 353008 6 vssd1
port 887 nsew ground bidirectional
rlabel metal4 s 19804 343552 20404 353008 6 vssd1
port 888 nsew ground bidirectional
rlabel metal4 s 559804 274192 560404 283648 6 vssd1
port 889 nsew ground bidirectional
rlabel metal4 s 523804 274192 524404 283648 6 vssd1
port 890 nsew ground bidirectional
rlabel metal4 s 451804 274192 452404 283648 6 vssd1
port 891 nsew ground bidirectional
rlabel metal4 s 415804 274192 416404 283648 6 vssd1
port 892 nsew ground bidirectional
rlabel metal4 s 379804 274192 380404 283648 6 vssd1
port 893 nsew ground bidirectional
rlabel metal4 s 343804 274192 344404 283648 6 vssd1
port 894 nsew ground bidirectional
rlabel metal4 s 307804 274192 308404 283648 6 vssd1
port 895 nsew ground bidirectional
rlabel metal4 s 235804 274192 236404 283648 6 vssd1
port 896 nsew ground bidirectional
rlabel metal4 s 199804 274192 200404 283648 6 vssd1
port 897 nsew ground bidirectional
rlabel metal4 s 163804 274192 164404 283648 6 vssd1
port 898 nsew ground bidirectional
rlabel metal4 s 127804 274192 128404 283648 6 vssd1
port 899 nsew ground bidirectional
rlabel metal4 s 55804 274192 56404 283648 6 vssd1
port 900 nsew ground bidirectional
rlabel metal4 s 19804 274192 20404 283648 6 vssd1
port 901 nsew ground bidirectional
rlabel metal4 s 559804 204832 560404 214288 6 vssd1
port 902 nsew ground bidirectional
rlabel metal4 s 523804 204832 524404 214288 6 vssd1
port 903 nsew ground bidirectional
rlabel metal4 s 451804 204832 452404 214288 6 vssd1
port 904 nsew ground bidirectional
rlabel metal4 s 415804 204832 416404 214288 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 379804 204832 380404 214288 6 vssd1
port 906 nsew ground bidirectional
rlabel metal4 s 343804 204832 344404 214288 6 vssd1
port 907 nsew ground bidirectional
rlabel metal4 s 307804 204832 308404 214288 6 vssd1
port 908 nsew ground bidirectional
rlabel metal4 s 235804 204832 236404 214288 6 vssd1
port 909 nsew ground bidirectional
rlabel metal4 s 199804 204832 200404 214288 6 vssd1
port 910 nsew ground bidirectional
rlabel metal4 s 163804 204832 164404 214288 6 vssd1
port 911 nsew ground bidirectional
rlabel metal4 s 127804 204832 128404 214288 6 vssd1
port 912 nsew ground bidirectional
rlabel metal4 s 55804 204832 56404 214288 6 vssd1
port 913 nsew ground bidirectional
rlabel metal4 s 19804 204832 20404 214288 6 vssd1
port 914 nsew ground bidirectional
rlabel metal4 s 559804 132152 560404 144928 6 vssd1
port 915 nsew ground bidirectional
rlabel metal4 s 523804 132152 524404 144928 6 vssd1
port 916 nsew ground bidirectional
rlabel metal4 s 451804 132152 452404 144928 6 vssd1
port 917 nsew ground bidirectional
rlabel metal4 s 415804 132152 416404 144928 6 vssd1
port 918 nsew ground bidirectional
rlabel metal4 s 379804 -1864 380404 144928 6 vssd1
port 919 nsew ground bidirectional
rlabel metal4 s 343804 132152 344404 144928 6 vssd1
port 920 nsew ground bidirectional
rlabel metal4 s 307804 -1864 308404 144928 6 vssd1
port 921 nsew ground bidirectional
rlabel metal4 s 235804 -1864 236404 144928 6 vssd1
port 922 nsew ground bidirectional
rlabel metal4 s 199804 132152 200404 144928 6 vssd1
port 923 nsew ground bidirectional
rlabel metal4 s 163804 -1864 164404 144928 6 vssd1
port 924 nsew ground bidirectional
rlabel metal4 s 127804 132152 128404 144928 6 vssd1
port 925 nsew ground bidirectional
rlabel metal4 s 55804 132152 56404 144928 6 vssd1
port 926 nsew ground bidirectional
rlabel metal4 s 19804 -1864 20404 144928 6 vssd1
port 927 nsew ground bidirectional
rlabel metal4 s 559804 -1864 560404 8248 6 vssd1
port 928 nsew ground bidirectional
rlabel metal4 s 523804 -1864 524404 8248 6 vssd1
port 929 nsew ground bidirectional
rlabel metal4 s 487804 -1864 488404 8248 6 vssd1
port 930 nsew ground bidirectional
rlabel metal4 s 451804 -1864 452404 8248 6 vssd1
port 931 nsew ground bidirectional
rlabel metal4 s 415804 -1864 416404 8248 6 vssd1
port 932 nsew ground bidirectional
rlabel metal4 s 343804 -1864 344404 8248 6 vssd1
port 933 nsew ground bidirectional
rlabel metal4 s 271804 -1864 272404 8248 6 vssd1
port 934 nsew ground bidirectional
rlabel metal4 s 199804 -1864 200404 8248 6 vssd1
port 935 nsew ground bidirectional
rlabel metal4 s 127804 -1864 128404 8248 6 vssd1
port 936 nsew ground bidirectional
rlabel metal4 s 55804 -1864 56404 8248 6 vssd1
port 937 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 938 nsew ground bidirectional
rlabel metal5 s -2936 668828 586860 669428 6 vssd1
port 939 nsew ground bidirectional
rlabel metal5 s -2936 632828 586860 633428 6 vssd1
port 940 nsew ground bidirectional
rlabel metal5 s -2936 596828 586860 597428 6 vssd1
port 941 nsew ground bidirectional
rlabel metal5 s -2936 560828 586860 561428 6 vssd1
port 942 nsew ground bidirectional
rlabel metal5 s -2936 524828 586860 525428 6 vssd1
port 943 nsew ground bidirectional
rlabel metal5 s -2936 488828 586860 489428 6 vssd1
port 944 nsew ground bidirectional
rlabel metal5 s -2936 452828 586860 453428 6 vssd1
port 945 nsew ground bidirectional
rlabel metal5 s -2936 416828 586860 417428 6 vssd1
port 946 nsew ground bidirectional
rlabel metal5 s -2936 380828 586860 381428 6 vssd1
port 947 nsew ground bidirectional
rlabel metal5 s -2936 344828 586860 345428 6 vssd1
port 948 nsew ground bidirectional
rlabel metal5 s -2936 308828 586860 309428 6 vssd1
port 949 nsew ground bidirectional
rlabel metal5 s -2936 272828 586860 273428 6 vssd1
port 950 nsew ground bidirectional
rlabel metal5 s -2936 236828 586860 237428 6 vssd1
port 951 nsew ground bidirectional
rlabel metal5 s -2936 200828 586860 201428 6 vssd1
port 952 nsew ground bidirectional
rlabel metal5 s -2936 164828 586860 165428 6 vssd1
port 953 nsew ground bidirectional
rlabel metal5 s -2936 128828 586860 129428 6 vssd1
port 954 nsew ground bidirectional
rlabel metal5 s -2936 92828 586860 93428 6 vssd1
port 955 nsew ground bidirectional
rlabel metal5 s -2936 56828 586860 57428 6 vssd1
port 956 nsew ground bidirectional
rlabel metal5 s -2936 20828 586860 21428 6 vssd1
port 957 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 958 nsew ground bidirectional
rlabel metal4 s 581404 -3744 582004 707680 6 vccd2
port 959 nsew power bidirectional
rlabel metal4 s 545404 690400 546004 707680 6 vccd2
port 960 nsew power bidirectional
rlabel metal4 s 509404 690400 510004 707680 6 vccd2
port 961 nsew power bidirectional
rlabel metal4 s 473404 690400 474004 707680 6 vccd2
port 962 nsew power bidirectional
rlabel metal4 s 437404 690400 438004 707680 6 vccd2
port 963 nsew power bidirectional
rlabel metal4 s 401404 132200 402004 707680 6 vccd2
port 964 nsew power bidirectional
rlabel metal4 s 365404 690400 366004 707680 6 vccd2
port 965 nsew power bidirectional
rlabel metal4 s 329404 690400 330004 707680 6 vccd2
port 966 nsew power bidirectional
rlabel metal4 s 293404 690400 294004 707680 6 vccd2
port 967 nsew power bidirectional
rlabel metal4 s 257404 690400 258004 707680 6 vccd2
port 968 nsew power bidirectional
rlabel metal4 s 221404 690400 222004 707680 6 vccd2
port 969 nsew power bidirectional
rlabel metal4 s 185404 690400 186004 707680 6 vccd2
port 970 nsew power bidirectional
rlabel metal4 s 149404 690400 150004 707680 6 vccd2
port 971 nsew power bidirectional
rlabel metal4 s 113404 690400 114004 707680 6 vccd2
port 972 nsew power bidirectional
rlabel metal4 s 77404 690400 78004 707680 6 vccd2
port 973 nsew power bidirectional
rlabel metal4 s 41404 690400 42004 707680 6 vccd2
port 974 nsew power bidirectional
rlabel metal4 s 5404 -3744 6004 707680 6 vccd2
port 975 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 976 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 977 nsew power bidirectional
rlabel metal4 s 545404 621040 546004 630400 6 vccd2
port 978 nsew power bidirectional
rlabel metal4 s 509404 621040 510004 630400 6 vccd2
port 979 nsew power bidirectional
rlabel metal4 s 473404 621040 474004 630400 6 vccd2
port 980 nsew power bidirectional
rlabel metal4 s 437404 621040 438004 630400 6 vccd2
port 981 nsew power bidirectional
rlabel metal4 s 365404 621040 366004 630400 6 vccd2
port 982 nsew power bidirectional
rlabel metal4 s 329404 621040 330004 630400 6 vccd2
port 983 nsew power bidirectional
rlabel metal4 s 293404 621040 294004 630400 6 vccd2
port 984 nsew power bidirectional
rlabel metal4 s 257404 621040 258004 630400 6 vccd2
port 985 nsew power bidirectional
rlabel metal4 s 221404 621040 222004 630400 6 vccd2
port 986 nsew power bidirectional
rlabel metal4 s 185404 621040 186004 630400 6 vccd2
port 987 nsew power bidirectional
rlabel metal4 s 149404 621040 150004 630400 6 vccd2
port 988 nsew power bidirectional
rlabel metal4 s 113404 621040 114004 630400 6 vccd2
port 989 nsew power bidirectional
rlabel metal4 s 77404 621040 78004 630400 6 vccd2
port 990 nsew power bidirectional
rlabel metal4 s 41404 621040 42004 630400 6 vccd2
port 991 nsew power bidirectional
rlabel metal4 s 545404 551680 546004 561040 6 vccd2
port 992 nsew power bidirectional
rlabel metal4 s 509404 551680 510004 561040 6 vccd2
port 993 nsew power bidirectional
rlabel metal4 s 473404 551680 474004 561040 6 vccd2
port 994 nsew power bidirectional
rlabel metal4 s 437404 551680 438004 561040 6 vccd2
port 995 nsew power bidirectional
rlabel metal4 s 365404 551680 366004 561040 6 vccd2
port 996 nsew power bidirectional
rlabel metal4 s 329404 551680 330004 561040 6 vccd2
port 997 nsew power bidirectional
rlabel metal4 s 293404 551680 294004 561040 6 vccd2
port 998 nsew power bidirectional
rlabel metal4 s 257404 551680 258004 561040 6 vccd2
port 999 nsew power bidirectional
rlabel metal4 s 221404 551680 222004 561040 6 vccd2
port 1000 nsew power bidirectional
rlabel metal4 s 185404 551680 186004 561040 6 vccd2
port 1001 nsew power bidirectional
rlabel metal4 s 149404 551680 150004 561040 6 vccd2
port 1002 nsew power bidirectional
rlabel metal4 s 113404 551680 114004 561040 6 vccd2
port 1003 nsew power bidirectional
rlabel metal4 s 77404 551680 78004 561040 6 vccd2
port 1004 nsew power bidirectional
rlabel metal4 s 41404 551680 42004 561040 6 vccd2
port 1005 nsew power bidirectional
rlabel metal4 s 545404 482320 546004 491680 6 vccd2
port 1006 nsew power bidirectional
rlabel metal4 s 509404 482320 510004 491680 6 vccd2
port 1007 nsew power bidirectional
rlabel metal4 s 473404 482320 474004 491680 6 vccd2
port 1008 nsew power bidirectional
rlabel metal4 s 437404 482320 438004 491680 6 vccd2
port 1009 nsew power bidirectional
rlabel metal4 s 365404 482320 366004 491680 6 vccd2
port 1010 nsew power bidirectional
rlabel metal4 s 329404 482320 330004 491680 6 vccd2
port 1011 nsew power bidirectional
rlabel metal4 s 293404 482320 294004 491680 6 vccd2
port 1012 nsew power bidirectional
rlabel metal4 s 257404 482320 258004 491680 6 vccd2
port 1013 nsew power bidirectional
rlabel metal4 s 221404 482320 222004 491680 6 vccd2
port 1014 nsew power bidirectional
rlabel metal4 s 185404 482320 186004 491680 6 vccd2
port 1015 nsew power bidirectional
rlabel metal4 s 149404 482320 150004 491680 6 vccd2
port 1016 nsew power bidirectional
rlabel metal4 s 113404 482320 114004 491680 6 vccd2
port 1017 nsew power bidirectional
rlabel metal4 s 77404 482320 78004 491680 6 vccd2
port 1018 nsew power bidirectional
rlabel metal4 s 41404 482320 42004 491680 6 vccd2
port 1019 nsew power bidirectional
rlabel metal4 s 545404 412960 546004 422320 6 vccd2
port 1020 nsew power bidirectional
rlabel metal4 s 509404 412960 510004 422320 6 vccd2
port 1021 nsew power bidirectional
rlabel metal4 s 473404 412960 474004 422320 6 vccd2
port 1022 nsew power bidirectional
rlabel metal4 s 437404 412960 438004 422320 6 vccd2
port 1023 nsew power bidirectional
rlabel metal4 s 365404 412960 366004 422320 6 vccd2
port 1024 nsew power bidirectional
rlabel metal4 s 329404 412960 330004 422320 6 vccd2
port 1025 nsew power bidirectional
rlabel metal4 s 293404 412960 294004 422320 6 vccd2
port 1026 nsew power bidirectional
rlabel metal4 s 257404 412960 258004 422320 6 vccd2
port 1027 nsew power bidirectional
rlabel metal4 s 221404 412960 222004 422320 6 vccd2
port 1028 nsew power bidirectional
rlabel metal4 s 185404 412960 186004 422320 6 vccd2
port 1029 nsew power bidirectional
rlabel metal4 s 149404 412960 150004 422320 6 vccd2
port 1030 nsew power bidirectional
rlabel metal4 s 113404 412960 114004 422320 6 vccd2
port 1031 nsew power bidirectional
rlabel metal4 s 77404 412960 78004 422320 6 vccd2
port 1032 nsew power bidirectional
rlabel metal4 s 41404 412960 42004 422320 6 vccd2
port 1033 nsew power bidirectional
rlabel metal4 s 545404 343600 546004 352960 6 vccd2
port 1034 nsew power bidirectional
rlabel metal4 s 509404 343600 510004 352960 6 vccd2
port 1035 nsew power bidirectional
rlabel metal4 s 473404 343600 474004 352960 6 vccd2
port 1036 nsew power bidirectional
rlabel metal4 s 437404 343600 438004 352960 6 vccd2
port 1037 nsew power bidirectional
rlabel metal4 s 365404 343600 366004 352960 6 vccd2
port 1038 nsew power bidirectional
rlabel metal4 s 329404 343600 330004 352960 6 vccd2
port 1039 nsew power bidirectional
rlabel metal4 s 293404 343600 294004 352960 6 vccd2
port 1040 nsew power bidirectional
rlabel metal4 s 257404 343600 258004 352960 6 vccd2
port 1041 nsew power bidirectional
rlabel metal4 s 221404 343600 222004 352960 6 vccd2
port 1042 nsew power bidirectional
rlabel metal4 s 185404 343600 186004 352960 6 vccd2
port 1043 nsew power bidirectional
rlabel metal4 s 149404 343600 150004 352960 6 vccd2
port 1044 nsew power bidirectional
rlabel metal4 s 113404 343600 114004 352960 6 vccd2
port 1045 nsew power bidirectional
rlabel metal4 s 77404 343600 78004 352960 6 vccd2
port 1046 nsew power bidirectional
rlabel metal4 s 41404 343600 42004 352960 6 vccd2
port 1047 nsew power bidirectional
rlabel metal4 s 545404 274240 546004 283600 6 vccd2
port 1048 nsew power bidirectional
rlabel metal4 s 509404 274240 510004 283600 6 vccd2
port 1049 nsew power bidirectional
rlabel metal4 s 473404 274240 474004 283600 6 vccd2
port 1050 nsew power bidirectional
rlabel metal4 s 437404 274240 438004 283600 6 vccd2
port 1051 nsew power bidirectional
rlabel metal4 s 365404 274240 366004 283600 6 vccd2
port 1052 nsew power bidirectional
rlabel metal4 s 329404 274240 330004 283600 6 vccd2
port 1053 nsew power bidirectional
rlabel metal4 s 293404 274240 294004 283600 6 vccd2
port 1054 nsew power bidirectional
rlabel metal4 s 257404 274240 258004 283600 6 vccd2
port 1055 nsew power bidirectional
rlabel metal4 s 221404 274240 222004 283600 6 vccd2
port 1056 nsew power bidirectional
rlabel metal4 s 185404 274240 186004 283600 6 vccd2
port 1057 nsew power bidirectional
rlabel metal4 s 149404 274240 150004 283600 6 vccd2
port 1058 nsew power bidirectional
rlabel metal4 s 113404 274240 114004 283600 6 vccd2
port 1059 nsew power bidirectional
rlabel metal4 s 77404 274240 78004 283600 6 vccd2
port 1060 nsew power bidirectional
rlabel metal4 s 41404 274240 42004 283600 6 vccd2
port 1061 nsew power bidirectional
rlabel metal4 s 545404 204880 546004 214240 6 vccd2
port 1062 nsew power bidirectional
rlabel metal4 s 509404 204880 510004 214240 6 vccd2
port 1063 nsew power bidirectional
rlabel metal4 s 473404 204880 474004 214240 6 vccd2
port 1064 nsew power bidirectional
rlabel metal4 s 437404 204880 438004 214240 6 vccd2
port 1065 nsew power bidirectional
rlabel metal4 s 365404 204880 366004 214240 6 vccd2
port 1066 nsew power bidirectional
rlabel metal4 s 329404 204880 330004 214240 6 vccd2
port 1067 nsew power bidirectional
rlabel metal4 s 293404 204880 294004 214240 6 vccd2
port 1068 nsew power bidirectional
rlabel metal4 s 257404 204880 258004 214240 6 vccd2
port 1069 nsew power bidirectional
rlabel metal4 s 221404 204880 222004 214240 6 vccd2
port 1070 nsew power bidirectional
rlabel metal4 s 185404 204880 186004 214240 6 vccd2
port 1071 nsew power bidirectional
rlabel metal4 s 149404 204880 150004 214240 6 vccd2
port 1072 nsew power bidirectional
rlabel metal4 s 113404 204880 114004 214240 6 vccd2
port 1073 nsew power bidirectional
rlabel metal4 s 77404 204880 78004 214240 6 vccd2
port 1074 nsew power bidirectional
rlabel metal4 s 41404 204880 42004 214240 6 vccd2
port 1075 nsew power bidirectional
rlabel metal4 s 545404 132200 546004 144880 6 vccd2
port 1076 nsew power bidirectional
rlabel metal4 s 509404 132200 510004 144880 6 vccd2
port 1077 nsew power bidirectional
rlabel metal4 s 473404 132200 474004 144880 6 vccd2
port 1078 nsew power bidirectional
rlabel metal4 s 437404 132200 438004 144880 6 vccd2
port 1079 nsew power bidirectional
rlabel metal4 s 365404 132200 366004 144880 6 vccd2
port 1080 nsew power bidirectional
rlabel metal4 s 329404 132200 330004 144880 6 vccd2
port 1081 nsew power bidirectional
rlabel metal4 s 293404 132200 294004 144880 6 vccd2
port 1082 nsew power bidirectional
rlabel metal4 s 257404 132200 258004 144880 6 vccd2
port 1083 nsew power bidirectional
rlabel metal4 s 221404 132200 222004 144880 6 vccd2
port 1084 nsew power bidirectional
rlabel metal4 s 185404 132200 186004 144880 6 vccd2
port 1085 nsew power bidirectional
rlabel metal4 s 149404 132200 150004 144880 6 vccd2
port 1086 nsew power bidirectional
rlabel metal4 s 113404 132200 114004 144880 6 vccd2
port 1087 nsew power bidirectional
rlabel metal4 s 77404 132200 78004 144880 6 vccd2
port 1088 nsew power bidirectional
rlabel metal4 s 41404 132200 42004 144880 6 vccd2
port 1089 nsew power bidirectional
rlabel metal4 s 545404 -3744 546004 8200 6 vccd2
port 1090 nsew power bidirectional
rlabel metal4 s 509404 -3744 510004 8200 6 vccd2
port 1091 nsew power bidirectional
rlabel metal4 s 473404 -3744 474004 8200 6 vccd2
port 1092 nsew power bidirectional
rlabel metal4 s 437404 -3744 438004 8200 6 vccd2
port 1093 nsew power bidirectional
rlabel metal4 s 401404 -3744 402004 8200 6 vccd2
port 1094 nsew power bidirectional
rlabel metal4 s 365404 -3744 366004 8200 6 vccd2
port 1095 nsew power bidirectional
rlabel metal4 s 329404 -3744 330004 8200 6 vccd2
port 1096 nsew power bidirectional
rlabel metal4 s 293404 -3744 294004 8200 6 vccd2
port 1097 nsew power bidirectional
rlabel metal4 s 257404 -3744 258004 8200 6 vccd2
port 1098 nsew power bidirectional
rlabel metal4 s 221404 -3744 222004 8200 6 vccd2
port 1099 nsew power bidirectional
rlabel metal4 s 185404 -3744 186004 8200 6 vccd2
port 1100 nsew power bidirectional
rlabel metal4 s 149404 -3744 150004 8200 6 vccd2
port 1101 nsew power bidirectional
rlabel metal4 s 113404 -3744 114004 8200 6 vccd2
port 1102 nsew power bidirectional
rlabel metal4 s 77404 -3744 78004 8200 6 vccd2
port 1103 nsew power bidirectional
rlabel metal4 s 41404 -3744 42004 8200 6 vccd2
port 1104 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 1105 nsew power bidirectional
rlabel metal5 s -4816 690476 588740 691076 6 vccd2
port 1106 nsew power bidirectional
rlabel metal5 s -4816 654476 588740 655076 6 vccd2
port 1107 nsew power bidirectional
rlabel metal5 s -4816 618476 588740 619076 6 vccd2
port 1108 nsew power bidirectional
rlabel metal5 s -4816 582476 588740 583076 6 vccd2
port 1109 nsew power bidirectional
rlabel metal5 s -4816 546476 588740 547076 6 vccd2
port 1110 nsew power bidirectional
rlabel metal5 s -4816 510476 588740 511076 6 vccd2
port 1111 nsew power bidirectional
rlabel metal5 s -4816 474476 588740 475076 6 vccd2
port 1112 nsew power bidirectional
rlabel metal5 s -4816 438476 588740 439076 6 vccd2
port 1113 nsew power bidirectional
rlabel metal5 s -4816 402476 588740 403076 6 vccd2
port 1114 nsew power bidirectional
rlabel metal5 s -4816 366476 588740 367076 6 vccd2
port 1115 nsew power bidirectional
rlabel metal5 s -4816 330476 588740 331076 6 vccd2
port 1116 nsew power bidirectional
rlabel metal5 s -4816 294476 588740 295076 6 vccd2
port 1117 nsew power bidirectional
rlabel metal5 s -4816 258476 588740 259076 6 vccd2
port 1118 nsew power bidirectional
rlabel metal5 s -4816 222476 588740 223076 6 vccd2
port 1119 nsew power bidirectional
rlabel metal5 s -4816 186476 588740 187076 6 vccd2
port 1120 nsew power bidirectional
rlabel metal5 s -4816 150476 588740 151076 6 vccd2
port 1121 nsew power bidirectional
rlabel metal5 s -4816 114476 588740 115076 6 vccd2
port 1122 nsew power bidirectional
rlabel metal5 s -4816 78476 588740 79076 6 vccd2
port 1123 nsew power bidirectional
rlabel metal5 s -4816 42476 588740 43076 6 vccd2
port 1124 nsew power bidirectional
rlabel metal5 s -4816 6476 588740 7076 6 vccd2
port 1125 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 1126 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 1127 nsew ground bidirectional
rlabel metal4 s 563404 690400 564004 707680 6 vssd2
port 1128 nsew ground bidirectional
rlabel metal4 s 527404 690400 528004 707680 6 vssd2
port 1129 nsew ground bidirectional
rlabel metal4 s 491404 132200 492004 707680 6 vssd2
port 1130 nsew ground bidirectional
rlabel metal4 s 455404 690400 456004 707680 6 vssd2
port 1131 nsew ground bidirectional
rlabel metal4 s 419404 690400 420004 707680 6 vssd2
port 1132 nsew ground bidirectional
rlabel metal4 s 383404 690400 384004 707680 6 vssd2
port 1133 nsew ground bidirectional
rlabel metal4 s 347404 690400 348004 707680 6 vssd2
port 1134 nsew ground bidirectional
rlabel metal4 s 311404 132200 312004 707680 6 vssd2
port 1135 nsew ground bidirectional
rlabel metal4 s 275404 690400 276004 707680 6 vssd2
port 1136 nsew ground bidirectional
rlabel metal4 s 239404 690400 240004 707680 6 vssd2
port 1137 nsew ground bidirectional
rlabel metal4 s 203404 690400 204004 707680 6 vssd2
port 1138 nsew ground bidirectional
rlabel metal4 s 167404 690400 168004 707680 6 vssd2
port 1139 nsew ground bidirectional
rlabel metal4 s 131404 690400 132004 707680 6 vssd2
port 1140 nsew ground bidirectional
rlabel metal4 s 95404 132200 96004 707680 6 vssd2
port 1141 nsew ground bidirectional
rlabel metal4 s 59404 690400 60004 707680 6 vssd2
port 1142 nsew ground bidirectional
rlabel metal4 s 23404 690400 24004 707680 6 vssd2
port 1143 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 1144 nsew ground bidirectional
rlabel metal4 s 563404 621040 564004 630400 6 vssd2
port 1145 nsew ground bidirectional
rlabel metal4 s 527404 621040 528004 630400 6 vssd2
port 1146 nsew ground bidirectional
rlabel metal4 s 455404 621040 456004 630400 6 vssd2
port 1147 nsew ground bidirectional
rlabel metal4 s 419404 621040 420004 630400 6 vssd2
port 1148 nsew ground bidirectional
rlabel metal4 s 383404 621040 384004 630400 6 vssd2
port 1149 nsew ground bidirectional
rlabel metal4 s 347404 621040 348004 630400 6 vssd2
port 1150 nsew ground bidirectional
rlabel metal4 s 275404 621040 276004 630400 6 vssd2
port 1151 nsew ground bidirectional
rlabel metal4 s 239404 621040 240004 630400 6 vssd2
port 1152 nsew ground bidirectional
rlabel metal4 s 203404 621040 204004 630400 6 vssd2
port 1153 nsew ground bidirectional
rlabel metal4 s 167404 621040 168004 630400 6 vssd2
port 1154 nsew ground bidirectional
rlabel metal4 s 131404 621040 132004 630400 6 vssd2
port 1155 nsew ground bidirectional
rlabel metal4 s 59404 621040 60004 630400 6 vssd2
port 1156 nsew ground bidirectional
rlabel metal4 s 23404 621040 24004 630400 6 vssd2
port 1157 nsew ground bidirectional
rlabel metal4 s 563404 551680 564004 561040 6 vssd2
port 1158 nsew ground bidirectional
rlabel metal4 s 527404 551680 528004 561040 6 vssd2
port 1159 nsew ground bidirectional
rlabel metal4 s 455404 551680 456004 561040 6 vssd2
port 1160 nsew ground bidirectional
rlabel metal4 s 419404 551680 420004 561040 6 vssd2
port 1161 nsew ground bidirectional
rlabel metal4 s 383404 551680 384004 561040 6 vssd2
port 1162 nsew ground bidirectional
rlabel metal4 s 347404 551680 348004 561040 6 vssd2
port 1163 nsew ground bidirectional
rlabel metal4 s 275404 551680 276004 561040 6 vssd2
port 1164 nsew ground bidirectional
rlabel metal4 s 239404 551680 240004 561040 6 vssd2
port 1165 nsew ground bidirectional
rlabel metal4 s 203404 551680 204004 561040 6 vssd2
port 1166 nsew ground bidirectional
rlabel metal4 s 167404 551680 168004 561040 6 vssd2
port 1167 nsew ground bidirectional
rlabel metal4 s 131404 551680 132004 561040 6 vssd2
port 1168 nsew ground bidirectional
rlabel metal4 s 59404 551680 60004 561040 6 vssd2
port 1169 nsew ground bidirectional
rlabel metal4 s 23404 551680 24004 561040 6 vssd2
port 1170 nsew ground bidirectional
rlabel metal4 s 563404 482320 564004 491680 6 vssd2
port 1171 nsew ground bidirectional
rlabel metal4 s 527404 482320 528004 491680 6 vssd2
port 1172 nsew ground bidirectional
rlabel metal4 s 455404 482320 456004 491680 6 vssd2
port 1173 nsew ground bidirectional
rlabel metal4 s 419404 482320 420004 491680 6 vssd2
port 1174 nsew ground bidirectional
rlabel metal4 s 383404 482320 384004 491680 6 vssd2
port 1175 nsew ground bidirectional
rlabel metal4 s 347404 482320 348004 491680 6 vssd2
port 1176 nsew ground bidirectional
rlabel metal4 s 275404 482320 276004 491680 6 vssd2
port 1177 nsew ground bidirectional
rlabel metal4 s 239404 482320 240004 491680 6 vssd2
port 1178 nsew ground bidirectional
rlabel metal4 s 203404 482320 204004 491680 6 vssd2
port 1179 nsew ground bidirectional
rlabel metal4 s 167404 482320 168004 491680 6 vssd2
port 1180 nsew ground bidirectional
rlabel metal4 s 131404 482320 132004 491680 6 vssd2
port 1181 nsew ground bidirectional
rlabel metal4 s 59404 482320 60004 491680 6 vssd2
port 1182 nsew ground bidirectional
rlabel metal4 s 23404 482320 24004 491680 6 vssd2
port 1183 nsew ground bidirectional
rlabel metal4 s 563404 412960 564004 422320 6 vssd2
port 1184 nsew ground bidirectional
rlabel metal4 s 527404 412960 528004 422320 6 vssd2
port 1185 nsew ground bidirectional
rlabel metal4 s 455404 412960 456004 422320 6 vssd2
port 1186 nsew ground bidirectional
rlabel metal4 s 419404 412960 420004 422320 6 vssd2
port 1187 nsew ground bidirectional
rlabel metal4 s 383404 412960 384004 422320 6 vssd2
port 1188 nsew ground bidirectional
rlabel metal4 s 347404 412960 348004 422320 6 vssd2
port 1189 nsew ground bidirectional
rlabel metal4 s 275404 412960 276004 422320 6 vssd2
port 1190 nsew ground bidirectional
rlabel metal4 s 239404 412960 240004 422320 6 vssd2
port 1191 nsew ground bidirectional
rlabel metal4 s 203404 412960 204004 422320 6 vssd2
port 1192 nsew ground bidirectional
rlabel metal4 s 167404 412960 168004 422320 6 vssd2
port 1193 nsew ground bidirectional
rlabel metal4 s 131404 412960 132004 422320 6 vssd2
port 1194 nsew ground bidirectional
rlabel metal4 s 59404 412960 60004 422320 6 vssd2
port 1195 nsew ground bidirectional
rlabel metal4 s 23404 412960 24004 422320 6 vssd2
port 1196 nsew ground bidirectional
rlabel metal4 s 563404 343600 564004 352960 6 vssd2
port 1197 nsew ground bidirectional
rlabel metal4 s 527404 343600 528004 352960 6 vssd2
port 1198 nsew ground bidirectional
rlabel metal4 s 455404 343600 456004 352960 6 vssd2
port 1199 nsew ground bidirectional
rlabel metal4 s 419404 343600 420004 352960 6 vssd2
port 1200 nsew ground bidirectional
rlabel metal4 s 383404 343600 384004 352960 6 vssd2
port 1201 nsew ground bidirectional
rlabel metal4 s 347404 343600 348004 352960 6 vssd2
port 1202 nsew ground bidirectional
rlabel metal4 s 275404 343600 276004 352960 6 vssd2
port 1203 nsew ground bidirectional
rlabel metal4 s 239404 343600 240004 352960 6 vssd2
port 1204 nsew ground bidirectional
rlabel metal4 s 203404 343600 204004 352960 6 vssd2
port 1205 nsew ground bidirectional
rlabel metal4 s 167404 343600 168004 352960 6 vssd2
port 1206 nsew ground bidirectional
rlabel metal4 s 131404 343600 132004 352960 6 vssd2
port 1207 nsew ground bidirectional
rlabel metal4 s 59404 343600 60004 352960 6 vssd2
port 1208 nsew ground bidirectional
rlabel metal4 s 23404 343600 24004 352960 6 vssd2
port 1209 nsew ground bidirectional
rlabel metal4 s 563404 274240 564004 283600 6 vssd2
port 1210 nsew ground bidirectional
rlabel metal4 s 527404 274240 528004 283600 6 vssd2
port 1211 nsew ground bidirectional
rlabel metal4 s 455404 274240 456004 283600 6 vssd2
port 1212 nsew ground bidirectional
rlabel metal4 s 419404 274240 420004 283600 6 vssd2
port 1213 nsew ground bidirectional
rlabel metal4 s 383404 274240 384004 283600 6 vssd2
port 1214 nsew ground bidirectional
rlabel metal4 s 347404 274240 348004 283600 6 vssd2
port 1215 nsew ground bidirectional
rlabel metal4 s 275404 274240 276004 283600 6 vssd2
port 1216 nsew ground bidirectional
rlabel metal4 s 239404 274240 240004 283600 6 vssd2
port 1217 nsew ground bidirectional
rlabel metal4 s 203404 274240 204004 283600 6 vssd2
port 1218 nsew ground bidirectional
rlabel metal4 s 167404 274240 168004 283600 6 vssd2
port 1219 nsew ground bidirectional
rlabel metal4 s 131404 274240 132004 283600 6 vssd2
port 1220 nsew ground bidirectional
rlabel metal4 s 59404 274240 60004 283600 6 vssd2
port 1221 nsew ground bidirectional
rlabel metal4 s 23404 274240 24004 283600 6 vssd2
port 1222 nsew ground bidirectional
rlabel metal4 s 563404 204880 564004 214240 6 vssd2
port 1223 nsew ground bidirectional
rlabel metal4 s 527404 204880 528004 214240 6 vssd2
port 1224 nsew ground bidirectional
rlabel metal4 s 455404 204880 456004 214240 6 vssd2
port 1225 nsew ground bidirectional
rlabel metal4 s 419404 204880 420004 214240 6 vssd2
port 1226 nsew ground bidirectional
rlabel metal4 s 383404 204880 384004 214240 6 vssd2
port 1227 nsew ground bidirectional
rlabel metal4 s 347404 204880 348004 214240 6 vssd2
port 1228 nsew ground bidirectional
rlabel metal4 s 275404 204880 276004 214240 6 vssd2
port 1229 nsew ground bidirectional
rlabel metal4 s 239404 204880 240004 214240 6 vssd2
port 1230 nsew ground bidirectional
rlabel metal4 s 203404 204880 204004 214240 6 vssd2
port 1231 nsew ground bidirectional
rlabel metal4 s 167404 204880 168004 214240 6 vssd2
port 1232 nsew ground bidirectional
rlabel metal4 s 131404 204880 132004 214240 6 vssd2
port 1233 nsew ground bidirectional
rlabel metal4 s 59404 204880 60004 214240 6 vssd2
port 1234 nsew ground bidirectional
rlabel metal4 s 23404 204880 24004 214240 6 vssd2
port 1235 nsew ground bidirectional
rlabel metal4 s 563404 132200 564004 144880 6 vssd2
port 1236 nsew ground bidirectional
rlabel metal4 s 527404 132200 528004 144880 6 vssd2
port 1237 nsew ground bidirectional
rlabel metal4 s 455404 132200 456004 144880 6 vssd2
port 1238 nsew ground bidirectional
rlabel metal4 s 419404 132200 420004 144880 6 vssd2
port 1239 nsew ground bidirectional
rlabel metal4 s 383404 -3744 384004 144880 6 vssd2
port 1240 nsew ground bidirectional
rlabel metal4 s 347404 132200 348004 144880 6 vssd2
port 1241 nsew ground bidirectional
rlabel metal4 s 275404 132200 276004 144880 6 vssd2
port 1242 nsew ground bidirectional
rlabel metal4 s 239404 132200 240004 144880 6 vssd2
port 1243 nsew ground bidirectional
rlabel metal4 s 203404 132200 204004 144880 6 vssd2
port 1244 nsew ground bidirectional
rlabel metal4 s 167404 132200 168004 144880 6 vssd2
port 1245 nsew ground bidirectional
rlabel metal4 s 131404 132200 132004 144880 6 vssd2
port 1246 nsew ground bidirectional
rlabel metal4 s 59404 132200 60004 144880 6 vssd2
port 1247 nsew ground bidirectional
rlabel metal4 s 23404 -3744 24004 144880 6 vssd2
port 1248 nsew ground bidirectional
rlabel metal4 s 563404 -3744 564004 8200 6 vssd2
port 1249 nsew ground bidirectional
rlabel metal4 s 527404 -3744 528004 8200 6 vssd2
port 1250 nsew ground bidirectional
rlabel metal4 s 491404 -3744 492004 8200 6 vssd2
port 1251 nsew ground bidirectional
rlabel metal4 s 455404 -3744 456004 8200 6 vssd2
port 1252 nsew ground bidirectional
rlabel metal4 s 419404 -3744 420004 8200 6 vssd2
port 1253 nsew ground bidirectional
rlabel metal4 s 347404 -3744 348004 8200 6 vssd2
port 1254 nsew ground bidirectional
rlabel metal4 s 311404 -3744 312004 8200 6 vssd2
port 1255 nsew ground bidirectional
rlabel metal4 s 275404 -3744 276004 8200 6 vssd2
port 1256 nsew ground bidirectional
rlabel metal4 s 239404 -3744 240004 8200 6 vssd2
port 1257 nsew ground bidirectional
rlabel metal4 s 203404 -3744 204004 8200 6 vssd2
port 1258 nsew ground bidirectional
rlabel metal4 s 167404 -3744 168004 8200 6 vssd2
port 1259 nsew ground bidirectional
rlabel metal4 s 131404 -3744 132004 8200 6 vssd2
port 1260 nsew ground bidirectional
rlabel metal4 s 95404 -3744 96004 8200 6 vssd2
port 1261 nsew ground bidirectional
rlabel metal4 s 59404 -3744 60004 8200 6 vssd2
port 1262 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 1263 nsew ground bidirectional
rlabel metal5 s -4816 672476 588740 673076 6 vssd2
port 1264 nsew ground bidirectional
rlabel metal5 s -4816 636476 588740 637076 6 vssd2
port 1265 nsew ground bidirectional
rlabel metal5 s -4816 600476 588740 601076 6 vssd2
port 1266 nsew ground bidirectional
rlabel metal5 s -4816 564476 588740 565076 6 vssd2
port 1267 nsew ground bidirectional
rlabel metal5 s -4816 528476 588740 529076 6 vssd2
port 1268 nsew ground bidirectional
rlabel metal5 s -4816 492476 588740 493076 6 vssd2
port 1269 nsew ground bidirectional
rlabel metal5 s -4816 456476 588740 457076 6 vssd2
port 1270 nsew ground bidirectional
rlabel metal5 s -4816 420476 588740 421076 6 vssd2
port 1271 nsew ground bidirectional
rlabel metal5 s -4816 384476 588740 385076 6 vssd2
port 1272 nsew ground bidirectional
rlabel metal5 s -4816 348476 588740 349076 6 vssd2
port 1273 nsew ground bidirectional
rlabel metal5 s -4816 312476 588740 313076 6 vssd2
port 1274 nsew ground bidirectional
rlabel metal5 s -4816 276476 588740 277076 6 vssd2
port 1275 nsew ground bidirectional
rlabel metal5 s -4816 240476 588740 241076 6 vssd2
port 1276 nsew ground bidirectional
rlabel metal5 s -4816 204476 588740 205076 6 vssd2
port 1277 nsew ground bidirectional
rlabel metal5 s -4816 168476 588740 169076 6 vssd2
port 1278 nsew ground bidirectional
rlabel metal5 s -4816 132476 588740 133076 6 vssd2
port 1279 nsew ground bidirectional
rlabel metal5 s -4816 96476 588740 97076 6 vssd2
port 1280 nsew ground bidirectional
rlabel metal5 s -4816 60476 588740 61076 6 vssd2
port 1281 nsew ground bidirectional
rlabel metal5 s -4816 24476 588740 25076 6 vssd2
port 1282 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 1283 nsew ground bidirectional
rlabel metal4 s 549004 690400 549604 709560 6 vdda1
port 1284 nsew power bidirectional
rlabel metal4 s 513004 690400 513604 709560 6 vdda1
port 1285 nsew power bidirectional
rlabel metal4 s 477004 690400 477604 709560 6 vdda1
port 1286 nsew power bidirectional
rlabel metal4 s 441004 690400 441604 709560 6 vdda1
port 1287 nsew power bidirectional
rlabel metal4 s 405004 690400 405604 709560 6 vdda1
port 1288 nsew power bidirectional
rlabel metal4 s 369004 690400 369604 709560 6 vdda1
port 1289 nsew power bidirectional
rlabel metal4 s 333004 690400 333604 709560 6 vdda1
port 1290 nsew power bidirectional
rlabel metal4 s 297004 690400 297604 709560 6 vdda1
port 1291 nsew power bidirectional
rlabel metal4 s 261004 690400 261604 709560 6 vdda1
port 1292 nsew power bidirectional
rlabel metal4 s 225004 132200 225604 709560 6 vdda1
port 1293 nsew power bidirectional
rlabel metal4 s 189004 690400 189604 709560 6 vdda1
port 1294 nsew power bidirectional
rlabel metal4 s 153004 690400 153604 709560 6 vdda1
port 1295 nsew power bidirectional
rlabel metal4 s 117004 690400 117604 709560 6 vdda1
port 1296 nsew power bidirectional
rlabel metal4 s 81004 -5624 81604 709560 6 vdda1
port 1297 nsew power bidirectional
rlabel metal4 s 45004 690400 45604 709560 6 vdda1
port 1298 nsew power bidirectional
rlabel metal4 s 9004 -5624 9604 709560 6 vdda1
port 1299 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 1300 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 1301 nsew power bidirectional
rlabel metal4 s 549004 621040 549604 630400 6 vdda1
port 1302 nsew power bidirectional
rlabel metal4 s 513004 621040 513604 630400 6 vdda1
port 1303 nsew power bidirectional
rlabel metal4 s 477004 621040 477604 630400 6 vdda1
port 1304 nsew power bidirectional
rlabel metal4 s 441004 621040 441604 630400 6 vdda1
port 1305 nsew power bidirectional
rlabel metal4 s 405004 621040 405604 630400 6 vdda1
port 1306 nsew power bidirectional
rlabel metal4 s 369004 621040 369604 630400 6 vdda1
port 1307 nsew power bidirectional
rlabel metal4 s 333004 621040 333604 630400 6 vdda1
port 1308 nsew power bidirectional
rlabel metal4 s 297004 621040 297604 630400 6 vdda1
port 1309 nsew power bidirectional
rlabel metal4 s 261004 621040 261604 630400 6 vdda1
port 1310 nsew power bidirectional
rlabel metal4 s 189004 621040 189604 630400 6 vdda1
port 1311 nsew power bidirectional
rlabel metal4 s 153004 621040 153604 630400 6 vdda1
port 1312 nsew power bidirectional
rlabel metal4 s 117004 621040 117604 630400 6 vdda1
port 1313 nsew power bidirectional
rlabel metal4 s 45004 621040 45604 630400 6 vdda1
port 1314 nsew power bidirectional
rlabel metal4 s 549004 551680 549604 561040 6 vdda1
port 1315 nsew power bidirectional
rlabel metal4 s 513004 551680 513604 561040 6 vdda1
port 1316 nsew power bidirectional
rlabel metal4 s 477004 551680 477604 561040 6 vdda1
port 1317 nsew power bidirectional
rlabel metal4 s 441004 551680 441604 561040 6 vdda1
port 1318 nsew power bidirectional
rlabel metal4 s 405004 551680 405604 561040 6 vdda1
port 1319 nsew power bidirectional
rlabel metal4 s 369004 551680 369604 561040 6 vdda1
port 1320 nsew power bidirectional
rlabel metal4 s 333004 551680 333604 561040 6 vdda1
port 1321 nsew power bidirectional
rlabel metal4 s 297004 551680 297604 561040 6 vdda1
port 1322 nsew power bidirectional
rlabel metal4 s 261004 551680 261604 561040 6 vdda1
port 1323 nsew power bidirectional
rlabel metal4 s 189004 551680 189604 561040 6 vdda1
port 1324 nsew power bidirectional
rlabel metal4 s 153004 551680 153604 561040 6 vdda1
port 1325 nsew power bidirectional
rlabel metal4 s 117004 551680 117604 561040 6 vdda1
port 1326 nsew power bidirectional
rlabel metal4 s 45004 551680 45604 561040 6 vdda1
port 1327 nsew power bidirectional
rlabel metal4 s 549004 482320 549604 491680 6 vdda1
port 1328 nsew power bidirectional
rlabel metal4 s 513004 482320 513604 491680 6 vdda1
port 1329 nsew power bidirectional
rlabel metal4 s 477004 482320 477604 491680 6 vdda1
port 1330 nsew power bidirectional
rlabel metal4 s 441004 482320 441604 491680 6 vdda1
port 1331 nsew power bidirectional
rlabel metal4 s 405004 482320 405604 491680 6 vdda1
port 1332 nsew power bidirectional
rlabel metal4 s 369004 482320 369604 491680 6 vdda1
port 1333 nsew power bidirectional
rlabel metal4 s 333004 482320 333604 491680 6 vdda1
port 1334 nsew power bidirectional
rlabel metal4 s 297004 482320 297604 491680 6 vdda1
port 1335 nsew power bidirectional
rlabel metal4 s 261004 482320 261604 491680 6 vdda1
port 1336 nsew power bidirectional
rlabel metal4 s 189004 482320 189604 491680 6 vdda1
port 1337 nsew power bidirectional
rlabel metal4 s 153004 482320 153604 491680 6 vdda1
port 1338 nsew power bidirectional
rlabel metal4 s 117004 482320 117604 491680 6 vdda1
port 1339 nsew power bidirectional
rlabel metal4 s 45004 482320 45604 491680 6 vdda1
port 1340 nsew power bidirectional
rlabel metal4 s 549004 412960 549604 422320 6 vdda1
port 1341 nsew power bidirectional
rlabel metal4 s 513004 412960 513604 422320 6 vdda1
port 1342 nsew power bidirectional
rlabel metal4 s 477004 412960 477604 422320 6 vdda1
port 1343 nsew power bidirectional
rlabel metal4 s 441004 412960 441604 422320 6 vdda1
port 1344 nsew power bidirectional
rlabel metal4 s 405004 412960 405604 422320 6 vdda1
port 1345 nsew power bidirectional
rlabel metal4 s 369004 412960 369604 422320 6 vdda1
port 1346 nsew power bidirectional
rlabel metal4 s 333004 412960 333604 422320 6 vdda1
port 1347 nsew power bidirectional
rlabel metal4 s 297004 412960 297604 422320 6 vdda1
port 1348 nsew power bidirectional
rlabel metal4 s 261004 412960 261604 422320 6 vdda1
port 1349 nsew power bidirectional
rlabel metal4 s 189004 412960 189604 422320 6 vdda1
port 1350 nsew power bidirectional
rlabel metal4 s 153004 412960 153604 422320 6 vdda1
port 1351 nsew power bidirectional
rlabel metal4 s 117004 412960 117604 422320 6 vdda1
port 1352 nsew power bidirectional
rlabel metal4 s 45004 412960 45604 422320 6 vdda1
port 1353 nsew power bidirectional
rlabel metal4 s 549004 343600 549604 352960 6 vdda1
port 1354 nsew power bidirectional
rlabel metal4 s 513004 343600 513604 352960 6 vdda1
port 1355 nsew power bidirectional
rlabel metal4 s 477004 343600 477604 352960 6 vdda1
port 1356 nsew power bidirectional
rlabel metal4 s 441004 343600 441604 352960 6 vdda1
port 1357 nsew power bidirectional
rlabel metal4 s 405004 343600 405604 352960 6 vdda1
port 1358 nsew power bidirectional
rlabel metal4 s 369004 343600 369604 352960 6 vdda1
port 1359 nsew power bidirectional
rlabel metal4 s 333004 343600 333604 352960 6 vdda1
port 1360 nsew power bidirectional
rlabel metal4 s 297004 343600 297604 352960 6 vdda1
port 1361 nsew power bidirectional
rlabel metal4 s 261004 343600 261604 352960 6 vdda1
port 1362 nsew power bidirectional
rlabel metal4 s 189004 343600 189604 352960 6 vdda1
port 1363 nsew power bidirectional
rlabel metal4 s 153004 343600 153604 352960 6 vdda1
port 1364 nsew power bidirectional
rlabel metal4 s 117004 343600 117604 352960 6 vdda1
port 1365 nsew power bidirectional
rlabel metal4 s 45004 343600 45604 352960 6 vdda1
port 1366 nsew power bidirectional
rlabel metal4 s 549004 274240 549604 283600 6 vdda1
port 1367 nsew power bidirectional
rlabel metal4 s 513004 274240 513604 283600 6 vdda1
port 1368 nsew power bidirectional
rlabel metal4 s 477004 274240 477604 283600 6 vdda1
port 1369 nsew power bidirectional
rlabel metal4 s 441004 274240 441604 283600 6 vdda1
port 1370 nsew power bidirectional
rlabel metal4 s 405004 274240 405604 283600 6 vdda1
port 1371 nsew power bidirectional
rlabel metal4 s 369004 274240 369604 283600 6 vdda1
port 1372 nsew power bidirectional
rlabel metal4 s 333004 274240 333604 283600 6 vdda1
port 1373 nsew power bidirectional
rlabel metal4 s 297004 274240 297604 283600 6 vdda1
port 1374 nsew power bidirectional
rlabel metal4 s 261004 274240 261604 283600 6 vdda1
port 1375 nsew power bidirectional
rlabel metal4 s 189004 274240 189604 283600 6 vdda1
port 1376 nsew power bidirectional
rlabel metal4 s 153004 274240 153604 283600 6 vdda1
port 1377 nsew power bidirectional
rlabel metal4 s 117004 274240 117604 283600 6 vdda1
port 1378 nsew power bidirectional
rlabel metal4 s 45004 274240 45604 283600 6 vdda1
port 1379 nsew power bidirectional
rlabel metal4 s 549004 204880 549604 214240 6 vdda1
port 1380 nsew power bidirectional
rlabel metal4 s 513004 204880 513604 214240 6 vdda1
port 1381 nsew power bidirectional
rlabel metal4 s 477004 204880 477604 214240 6 vdda1
port 1382 nsew power bidirectional
rlabel metal4 s 441004 204880 441604 214240 6 vdda1
port 1383 nsew power bidirectional
rlabel metal4 s 405004 204880 405604 214240 6 vdda1
port 1384 nsew power bidirectional
rlabel metal4 s 369004 204880 369604 214240 6 vdda1
port 1385 nsew power bidirectional
rlabel metal4 s 333004 204880 333604 214240 6 vdda1
port 1386 nsew power bidirectional
rlabel metal4 s 297004 204880 297604 214240 6 vdda1
port 1387 nsew power bidirectional
rlabel metal4 s 261004 204880 261604 214240 6 vdda1
port 1388 nsew power bidirectional
rlabel metal4 s 189004 204880 189604 214240 6 vdda1
port 1389 nsew power bidirectional
rlabel metal4 s 153004 204880 153604 214240 6 vdda1
port 1390 nsew power bidirectional
rlabel metal4 s 117004 204880 117604 214240 6 vdda1
port 1391 nsew power bidirectional
rlabel metal4 s 45004 204880 45604 214240 6 vdda1
port 1392 nsew power bidirectional
rlabel metal4 s 549004 132200 549604 144880 6 vdda1
port 1393 nsew power bidirectional
rlabel metal4 s 513004 132200 513604 144880 6 vdda1
port 1394 nsew power bidirectional
rlabel metal4 s 477004 132200 477604 144880 6 vdda1
port 1395 nsew power bidirectional
rlabel metal4 s 441004 132200 441604 144880 6 vdda1
port 1396 nsew power bidirectional
rlabel metal4 s 405004 132200 405604 144880 6 vdda1
port 1397 nsew power bidirectional
rlabel metal4 s 369004 132200 369604 144880 6 vdda1
port 1398 nsew power bidirectional
rlabel metal4 s 333004 132200 333604 144880 6 vdda1
port 1399 nsew power bidirectional
rlabel metal4 s 297004 132200 297604 144880 6 vdda1
port 1400 nsew power bidirectional
rlabel metal4 s 261004 132200 261604 144880 6 vdda1
port 1401 nsew power bidirectional
rlabel metal4 s 189004 132200 189604 144880 6 vdda1
port 1402 nsew power bidirectional
rlabel metal4 s 153004 132200 153604 144880 6 vdda1
port 1403 nsew power bidirectional
rlabel metal4 s 117004 132200 117604 144880 6 vdda1
port 1404 nsew power bidirectional
rlabel metal4 s 45004 132200 45604 144880 6 vdda1
port 1405 nsew power bidirectional
rlabel metal4 s 549004 -5624 549604 8200 6 vdda1
port 1406 nsew power bidirectional
rlabel metal4 s 513004 -5624 513604 8200 6 vdda1
port 1407 nsew power bidirectional
rlabel metal4 s 477004 -5624 477604 8200 6 vdda1
port 1408 nsew power bidirectional
rlabel metal4 s 441004 -5624 441604 8200 6 vdda1
port 1409 nsew power bidirectional
rlabel metal4 s 405004 -5624 405604 8200 6 vdda1
port 1410 nsew power bidirectional
rlabel metal4 s 369004 -5624 369604 8200 6 vdda1
port 1411 nsew power bidirectional
rlabel metal4 s 333004 -5624 333604 8200 6 vdda1
port 1412 nsew power bidirectional
rlabel metal4 s 297004 -5624 297604 8200 6 vdda1
port 1413 nsew power bidirectional
rlabel metal4 s 261004 -5624 261604 8200 6 vdda1
port 1414 nsew power bidirectional
rlabel metal4 s 225004 -5624 225604 8200 6 vdda1
port 1415 nsew power bidirectional
rlabel metal4 s 189004 -5624 189604 8200 6 vdda1
port 1416 nsew power bidirectional
rlabel metal4 s 153004 -5624 153604 8200 6 vdda1
port 1417 nsew power bidirectional
rlabel metal4 s 117004 -5624 117604 8200 6 vdda1
port 1418 nsew power bidirectional
rlabel metal4 s 45004 -5624 45604 8200 6 vdda1
port 1419 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 1420 nsew power bidirectional
rlabel metal5 s -6696 694076 590620 694676 6 vdda1
port 1421 nsew power bidirectional
rlabel metal5 s -6696 658076 590620 658676 6 vdda1
port 1422 nsew power bidirectional
rlabel metal5 s -6696 622076 590620 622676 6 vdda1
port 1423 nsew power bidirectional
rlabel metal5 s -6696 586076 590620 586676 6 vdda1
port 1424 nsew power bidirectional
rlabel metal5 s -6696 550076 590620 550676 6 vdda1
port 1425 nsew power bidirectional
rlabel metal5 s -6696 514076 590620 514676 6 vdda1
port 1426 nsew power bidirectional
rlabel metal5 s -6696 478076 590620 478676 6 vdda1
port 1427 nsew power bidirectional
rlabel metal5 s -6696 442076 590620 442676 6 vdda1
port 1428 nsew power bidirectional
rlabel metal5 s -6696 406076 590620 406676 6 vdda1
port 1429 nsew power bidirectional
rlabel metal5 s -6696 370076 590620 370676 6 vdda1
port 1430 nsew power bidirectional
rlabel metal5 s -6696 334076 590620 334676 6 vdda1
port 1431 nsew power bidirectional
rlabel metal5 s -6696 298076 590620 298676 6 vdda1
port 1432 nsew power bidirectional
rlabel metal5 s -6696 262076 590620 262676 6 vdda1
port 1433 nsew power bidirectional
rlabel metal5 s -6696 226076 590620 226676 6 vdda1
port 1434 nsew power bidirectional
rlabel metal5 s -6696 190076 590620 190676 6 vdda1
port 1435 nsew power bidirectional
rlabel metal5 s -6696 154076 590620 154676 6 vdda1
port 1436 nsew power bidirectional
rlabel metal5 s -6696 118076 590620 118676 6 vdda1
port 1437 nsew power bidirectional
rlabel metal5 s -6696 82076 590620 82676 6 vdda1
port 1438 nsew power bidirectional
rlabel metal5 s -6696 46076 590620 46676 6 vdda1
port 1439 nsew power bidirectional
rlabel metal5 s -6696 10076 590620 10676 6 vdda1
port 1440 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 1441 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 1442 nsew ground bidirectional
rlabel metal4 s 567004 690400 567604 709560 6 vssa1
port 1443 nsew ground bidirectional
rlabel metal4 s 531004 690400 531604 709560 6 vssa1
port 1444 nsew ground bidirectional
rlabel metal4 s 495004 690400 495604 709560 6 vssa1
port 1445 nsew ground bidirectional
rlabel metal4 s 459004 690400 459604 709560 6 vssa1
port 1446 nsew ground bidirectional
rlabel metal4 s 423004 690400 423604 709560 6 vssa1
port 1447 nsew ground bidirectional
rlabel metal4 s 387004 690400 387604 709560 6 vssa1
port 1448 nsew ground bidirectional
rlabel metal4 s 351004 690400 351604 709560 6 vssa1
port 1449 nsew ground bidirectional
rlabel metal4 s 315004 132200 315604 709560 6 vssa1
port 1450 nsew ground bidirectional
rlabel metal4 s 279004 690400 279604 709560 6 vssa1
port 1451 nsew ground bidirectional
rlabel metal4 s 243004 690400 243604 709560 6 vssa1
port 1452 nsew ground bidirectional
rlabel metal4 s 207004 690400 207604 709560 6 vssa1
port 1453 nsew ground bidirectional
rlabel metal4 s 171004 690400 171604 709560 6 vssa1
port 1454 nsew ground bidirectional
rlabel metal4 s 135004 132200 135604 709560 6 vssa1
port 1455 nsew ground bidirectional
rlabel metal4 s 99004 690400 99604 709560 6 vssa1
port 1456 nsew ground bidirectional
rlabel metal4 s 63004 690400 63604 709560 6 vssa1
port 1457 nsew ground bidirectional
rlabel metal4 s 27004 690400 27604 709560 6 vssa1
port 1458 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 1459 nsew ground bidirectional
rlabel metal4 s 567004 621040 567604 630400 6 vssa1
port 1460 nsew ground bidirectional
rlabel metal4 s 531004 621040 531604 630400 6 vssa1
port 1461 nsew ground bidirectional
rlabel metal4 s 495004 621040 495604 630400 6 vssa1
port 1462 nsew ground bidirectional
rlabel metal4 s 459004 621040 459604 630400 6 vssa1
port 1463 nsew ground bidirectional
rlabel metal4 s 423004 621040 423604 630400 6 vssa1
port 1464 nsew ground bidirectional
rlabel metal4 s 387004 621040 387604 630400 6 vssa1
port 1465 nsew ground bidirectional
rlabel metal4 s 351004 621040 351604 630400 6 vssa1
port 1466 nsew ground bidirectional
rlabel metal4 s 279004 621040 279604 630400 6 vssa1
port 1467 nsew ground bidirectional
rlabel metal4 s 243004 621040 243604 630400 6 vssa1
port 1468 nsew ground bidirectional
rlabel metal4 s 207004 621040 207604 630400 6 vssa1
port 1469 nsew ground bidirectional
rlabel metal4 s 171004 621040 171604 630400 6 vssa1
port 1470 nsew ground bidirectional
rlabel metal4 s 99004 621040 99604 630400 6 vssa1
port 1471 nsew ground bidirectional
rlabel metal4 s 63004 621040 63604 630400 6 vssa1
port 1472 nsew ground bidirectional
rlabel metal4 s 27004 621040 27604 630400 6 vssa1
port 1473 nsew ground bidirectional
rlabel metal4 s 567004 551680 567604 561040 6 vssa1
port 1474 nsew ground bidirectional
rlabel metal4 s 531004 551680 531604 561040 6 vssa1
port 1475 nsew ground bidirectional
rlabel metal4 s 495004 551680 495604 561040 6 vssa1
port 1476 nsew ground bidirectional
rlabel metal4 s 459004 551680 459604 561040 6 vssa1
port 1477 nsew ground bidirectional
rlabel metal4 s 423004 551680 423604 561040 6 vssa1
port 1478 nsew ground bidirectional
rlabel metal4 s 387004 551680 387604 561040 6 vssa1
port 1479 nsew ground bidirectional
rlabel metal4 s 351004 551680 351604 561040 6 vssa1
port 1480 nsew ground bidirectional
rlabel metal4 s 279004 551680 279604 561040 6 vssa1
port 1481 nsew ground bidirectional
rlabel metal4 s 243004 551680 243604 561040 6 vssa1
port 1482 nsew ground bidirectional
rlabel metal4 s 207004 551680 207604 561040 6 vssa1
port 1483 nsew ground bidirectional
rlabel metal4 s 171004 551680 171604 561040 6 vssa1
port 1484 nsew ground bidirectional
rlabel metal4 s 99004 551680 99604 561040 6 vssa1
port 1485 nsew ground bidirectional
rlabel metal4 s 63004 551680 63604 561040 6 vssa1
port 1486 nsew ground bidirectional
rlabel metal4 s 27004 551680 27604 561040 6 vssa1
port 1487 nsew ground bidirectional
rlabel metal4 s 567004 482320 567604 491680 6 vssa1
port 1488 nsew ground bidirectional
rlabel metal4 s 531004 482320 531604 491680 6 vssa1
port 1489 nsew ground bidirectional
rlabel metal4 s 495004 482320 495604 491680 6 vssa1
port 1490 nsew ground bidirectional
rlabel metal4 s 459004 482320 459604 491680 6 vssa1
port 1491 nsew ground bidirectional
rlabel metal4 s 423004 482320 423604 491680 6 vssa1
port 1492 nsew ground bidirectional
rlabel metal4 s 387004 482320 387604 491680 6 vssa1
port 1493 nsew ground bidirectional
rlabel metal4 s 351004 482320 351604 491680 6 vssa1
port 1494 nsew ground bidirectional
rlabel metal4 s 279004 482320 279604 491680 6 vssa1
port 1495 nsew ground bidirectional
rlabel metal4 s 243004 482320 243604 491680 6 vssa1
port 1496 nsew ground bidirectional
rlabel metal4 s 207004 482320 207604 491680 6 vssa1
port 1497 nsew ground bidirectional
rlabel metal4 s 171004 482320 171604 491680 6 vssa1
port 1498 nsew ground bidirectional
rlabel metal4 s 99004 482320 99604 491680 6 vssa1
port 1499 nsew ground bidirectional
rlabel metal4 s 63004 482320 63604 491680 6 vssa1
port 1500 nsew ground bidirectional
rlabel metal4 s 27004 482320 27604 491680 6 vssa1
port 1501 nsew ground bidirectional
rlabel metal4 s 567004 412960 567604 422320 6 vssa1
port 1502 nsew ground bidirectional
rlabel metal4 s 531004 412960 531604 422320 6 vssa1
port 1503 nsew ground bidirectional
rlabel metal4 s 495004 412960 495604 422320 6 vssa1
port 1504 nsew ground bidirectional
rlabel metal4 s 459004 412960 459604 422320 6 vssa1
port 1505 nsew ground bidirectional
rlabel metal4 s 423004 412960 423604 422320 6 vssa1
port 1506 nsew ground bidirectional
rlabel metal4 s 387004 412960 387604 422320 6 vssa1
port 1507 nsew ground bidirectional
rlabel metal4 s 351004 412960 351604 422320 6 vssa1
port 1508 nsew ground bidirectional
rlabel metal4 s 279004 412960 279604 422320 6 vssa1
port 1509 nsew ground bidirectional
rlabel metal4 s 243004 412960 243604 422320 6 vssa1
port 1510 nsew ground bidirectional
rlabel metal4 s 207004 412960 207604 422320 6 vssa1
port 1511 nsew ground bidirectional
rlabel metal4 s 171004 412960 171604 422320 6 vssa1
port 1512 nsew ground bidirectional
rlabel metal4 s 99004 412960 99604 422320 6 vssa1
port 1513 nsew ground bidirectional
rlabel metal4 s 63004 412960 63604 422320 6 vssa1
port 1514 nsew ground bidirectional
rlabel metal4 s 27004 412960 27604 422320 6 vssa1
port 1515 nsew ground bidirectional
rlabel metal4 s 567004 343600 567604 352960 6 vssa1
port 1516 nsew ground bidirectional
rlabel metal4 s 531004 343600 531604 352960 6 vssa1
port 1517 nsew ground bidirectional
rlabel metal4 s 495004 343600 495604 352960 6 vssa1
port 1518 nsew ground bidirectional
rlabel metal4 s 459004 343600 459604 352960 6 vssa1
port 1519 nsew ground bidirectional
rlabel metal4 s 423004 343600 423604 352960 6 vssa1
port 1520 nsew ground bidirectional
rlabel metal4 s 387004 343600 387604 352960 6 vssa1
port 1521 nsew ground bidirectional
rlabel metal4 s 351004 343600 351604 352960 6 vssa1
port 1522 nsew ground bidirectional
rlabel metal4 s 279004 343600 279604 352960 6 vssa1
port 1523 nsew ground bidirectional
rlabel metal4 s 243004 343600 243604 352960 6 vssa1
port 1524 nsew ground bidirectional
rlabel metal4 s 207004 343600 207604 352960 6 vssa1
port 1525 nsew ground bidirectional
rlabel metal4 s 171004 343600 171604 352960 6 vssa1
port 1526 nsew ground bidirectional
rlabel metal4 s 99004 343600 99604 352960 6 vssa1
port 1527 nsew ground bidirectional
rlabel metal4 s 63004 343600 63604 352960 6 vssa1
port 1528 nsew ground bidirectional
rlabel metal4 s 27004 343600 27604 352960 6 vssa1
port 1529 nsew ground bidirectional
rlabel metal4 s 567004 274240 567604 283600 6 vssa1
port 1530 nsew ground bidirectional
rlabel metal4 s 531004 274240 531604 283600 6 vssa1
port 1531 nsew ground bidirectional
rlabel metal4 s 495004 274240 495604 283600 6 vssa1
port 1532 nsew ground bidirectional
rlabel metal4 s 459004 274240 459604 283600 6 vssa1
port 1533 nsew ground bidirectional
rlabel metal4 s 423004 274240 423604 283600 6 vssa1
port 1534 nsew ground bidirectional
rlabel metal4 s 387004 274240 387604 283600 6 vssa1
port 1535 nsew ground bidirectional
rlabel metal4 s 351004 274240 351604 283600 6 vssa1
port 1536 nsew ground bidirectional
rlabel metal4 s 279004 274240 279604 283600 6 vssa1
port 1537 nsew ground bidirectional
rlabel metal4 s 243004 274240 243604 283600 6 vssa1
port 1538 nsew ground bidirectional
rlabel metal4 s 207004 274240 207604 283600 6 vssa1
port 1539 nsew ground bidirectional
rlabel metal4 s 171004 274240 171604 283600 6 vssa1
port 1540 nsew ground bidirectional
rlabel metal4 s 99004 274240 99604 283600 6 vssa1
port 1541 nsew ground bidirectional
rlabel metal4 s 63004 274240 63604 283600 6 vssa1
port 1542 nsew ground bidirectional
rlabel metal4 s 27004 274240 27604 283600 6 vssa1
port 1543 nsew ground bidirectional
rlabel metal4 s 567004 204880 567604 214240 6 vssa1
port 1544 nsew ground bidirectional
rlabel metal4 s 531004 204880 531604 214240 6 vssa1
port 1545 nsew ground bidirectional
rlabel metal4 s 495004 204880 495604 214240 6 vssa1
port 1546 nsew ground bidirectional
rlabel metal4 s 459004 204880 459604 214240 6 vssa1
port 1547 nsew ground bidirectional
rlabel metal4 s 423004 204880 423604 214240 6 vssa1
port 1548 nsew ground bidirectional
rlabel metal4 s 387004 204880 387604 214240 6 vssa1
port 1549 nsew ground bidirectional
rlabel metal4 s 351004 204880 351604 214240 6 vssa1
port 1550 nsew ground bidirectional
rlabel metal4 s 279004 204880 279604 214240 6 vssa1
port 1551 nsew ground bidirectional
rlabel metal4 s 243004 204880 243604 214240 6 vssa1
port 1552 nsew ground bidirectional
rlabel metal4 s 207004 204880 207604 214240 6 vssa1
port 1553 nsew ground bidirectional
rlabel metal4 s 171004 204880 171604 214240 6 vssa1
port 1554 nsew ground bidirectional
rlabel metal4 s 99004 204880 99604 214240 6 vssa1
port 1555 nsew ground bidirectional
rlabel metal4 s 63004 204880 63604 214240 6 vssa1
port 1556 nsew ground bidirectional
rlabel metal4 s 27004 204880 27604 214240 6 vssa1
port 1557 nsew ground bidirectional
rlabel metal4 s 567004 132200 567604 144880 6 vssa1
port 1558 nsew ground bidirectional
rlabel metal4 s 531004 132200 531604 144880 6 vssa1
port 1559 nsew ground bidirectional
rlabel metal4 s 495004 132200 495604 144880 6 vssa1
port 1560 nsew ground bidirectional
rlabel metal4 s 459004 132200 459604 144880 6 vssa1
port 1561 nsew ground bidirectional
rlabel metal4 s 423004 132200 423604 144880 6 vssa1
port 1562 nsew ground bidirectional
rlabel metal4 s 387004 132200 387604 144880 6 vssa1
port 1563 nsew ground bidirectional
rlabel metal4 s 351004 132200 351604 144880 6 vssa1
port 1564 nsew ground bidirectional
rlabel metal4 s 279004 132200 279604 144880 6 vssa1
port 1565 nsew ground bidirectional
rlabel metal4 s 243004 132200 243604 144880 6 vssa1
port 1566 nsew ground bidirectional
rlabel metal4 s 207004 132200 207604 144880 6 vssa1
port 1567 nsew ground bidirectional
rlabel metal4 s 171004 132200 171604 144880 6 vssa1
port 1568 nsew ground bidirectional
rlabel metal4 s 99004 132200 99604 144880 6 vssa1
port 1569 nsew ground bidirectional
rlabel metal4 s 63004 132200 63604 144880 6 vssa1
port 1570 nsew ground bidirectional
rlabel metal4 s 27004 -5624 27604 144880 6 vssa1
port 1571 nsew ground bidirectional
rlabel metal4 s 567004 -5624 567604 8200 6 vssa1
port 1572 nsew ground bidirectional
rlabel metal4 s 531004 -5624 531604 8200 6 vssa1
port 1573 nsew ground bidirectional
rlabel metal4 s 495004 -5624 495604 8200 6 vssa1
port 1574 nsew ground bidirectional
rlabel metal4 s 459004 -5624 459604 8200 6 vssa1
port 1575 nsew ground bidirectional
rlabel metal4 s 423004 -5624 423604 8200 6 vssa1
port 1576 nsew ground bidirectional
rlabel metal4 s 387004 -5624 387604 8200 6 vssa1
port 1577 nsew ground bidirectional
rlabel metal4 s 351004 -5624 351604 8200 6 vssa1
port 1578 nsew ground bidirectional
rlabel metal4 s 315004 -5624 315604 8200 6 vssa1
port 1579 nsew ground bidirectional
rlabel metal4 s 279004 -5624 279604 8200 6 vssa1
port 1580 nsew ground bidirectional
rlabel metal4 s 243004 -5624 243604 8200 6 vssa1
port 1581 nsew ground bidirectional
rlabel metal4 s 207004 -5624 207604 8200 6 vssa1
port 1582 nsew ground bidirectional
rlabel metal4 s 171004 -5624 171604 8200 6 vssa1
port 1583 nsew ground bidirectional
rlabel metal4 s 135004 -5624 135604 8200 6 vssa1
port 1584 nsew ground bidirectional
rlabel metal4 s 99004 -5624 99604 8200 6 vssa1
port 1585 nsew ground bidirectional
rlabel metal4 s 63004 -5624 63604 8200 6 vssa1
port 1586 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 1587 nsew ground bidirectional
rlabel metal5 s -6696 676076 590620 676676 6 vssa1
port 1588 nsew ground bidirectional
rlabel metal5 s -6696 640076 590620 640676 6 vssa1
port 1589 nsew ground bidirectional
rlabel metal5 s -6696 604076 590620 604676 6 vssa1
port 1590 nsew ground bidirectional
rlabel metal5 s -6696 568076 590620 568676 6 vssa1
port 1591 nsew ground bidirectional
rlabel metal5 s -6696 532076 590620 532676 6 vssa1
port 1592 nsew ground bidirectional
rlabel metal5 s -6696 496076 590620 496676 6 vssa1
port 1593 nsew ground bidirectional
rlabel metal5 s -6696 460076 590620 460676 6 vssa1
port 1594 nsew ground bidirectional
rlabel metal5 s -6696 424076 590620 424676 6 vssa1
port 1595 nsew ground bidirectional
rlabel metal5 s -6696 388076 590620 388676 6 vssa1
port 1596 nsew ground bidirectional
rlabel metal5 s -6696 352076 590620 352676 6 vssa1
port 1597 nsew ground bidirectional
rlabel metal5 s -6696 316076 590620 316676 6 vssa1
port 1598 nsew ground bidirectional
rlabel metal5 s -6696 280076 590620 280676 6 vssa1
port 1599 nsew ground bidirectional
rlabel metal5 s -6696 244076 590620 244676 6 vssa1
port 1600 nsew ground bidirectional
rlabel metal5 s -6696 208076 590620 208676 6 vssa1
port 1601 nsew ground bidirectional
rlabel metal5 s -6696 172076 590620 172676 6 vssa1
port 1602 nsew ground bidirectional
rlabel metal5 s -6696 136076 590620 136676 6 vssa1
port 1603 nsew ground bidirectional
rlabel metal5 s -6696 100076 590620 100676 6 vssa1
port 1604 nsew ground bidirectional
rlabel metal5 s -6696 64076 590620 64676 6 vssa1
port 1605 nsew ground bidirectional
rlabel metal5 s -6696 28076 590620 28676 6 vssa1
port 1606 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 1607 nsew ground bidirectional
rlabel metal4 s 552604 690400 553204 711440 6 vdda2
port 1608 nsew power bidirectional
rlabel metal4 s 516604 690400 517204 711440 6 vdda2
port 1609 nsew power bidirectional
rlabel metal4 s 480604 690400 481204 711440 6 vdda2
port 1610 nsew power bidirectional
rlabel metal4 s 444604 132200 445204 711440 6 vdda2
port 1611 nsew power bidirectional
rlabel metal4 s 408604 690400 409204 711440 6 vdda2
port 1612 nsew power bidirectional
rlabel metal4 s 372604 690400 373204 711440 6 vdda2
port 1613 nsew power bidirectional
rlabel metal4 s 336604 690400 337204 711440 6 vdda2
port 1614 nsew power bidirectional
rlabel metal4 s 300604 690400 301204 711440 6 vdda2
port 1615 nsew power bidirectional
rlabel metal4 s 264604 690400 265204 711440 6 vdda2
port 1616 nsew power bidirectional
rlabel metal4 s 228604 690400 229204 711440 6 vdda2
port 1617 nsew power bidirectional
rlabel metal4 s 192604 690400 193204 711440 6 vdda2
port 1618 nsew power bidirectional
rlabel metal4 s 156604 690400 157204 711440 6 vdda2
port 1619 nsew power bidirectional
rlabel metal4 s 120604 690400 121204 711440 6 vdda2
port 1620 nsew power bidirectional
rlabel metal4 s 84604 -7504 85204 711440 6 vdda2
port 1621 nsew power bidirectional
rlabel metal4 s 48604 690400 49204 711440 6 vdda2
port 1622 nsew power bidirectional
rlabel metal4 s 12604 -7504 13204 711440 6 vdda2
port 1623 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 1624 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 1625 nsew power bidirectional
rlabel metal4 s 552604 621040 553204 630400 6 vdda2
port 1626 nsew power bidirectional
rlabel metal4 s 516604 621040 517204 630400 6 vdda2
port 1627 nsew power bidirectional
rlabel metal4 s 480604 621040 481204 630400 6 vdda2
port 1628 nsew power bidirectional
rlabel metal4 s 408604 621040 409204 630400 6 vdda2
port 1629 nsew power bidirectional
rlabel metal4 s 372604 621040 373204 630400 6 vdda2
port 1630 nsew power bidirectional
rlabel metal4 s 336604 621040 337204 630400 6 vdda2
port 1631 nsew power bidirectional
rlabel metal4 s 300604 621040 301204 630400 6 vdda2
port 1632 nsew power bidirectional
rlabel metal4 s 264604 621040 265204 630400 6 vdda2
port 1633 nsew power bidirectional
rlabel metal4 s 228604 621040 229204 630400 6 vdda2
port 1634 nsew power bidirectional
rlabel metal4 s 192604 621040 193204 630400 6 vdda2
port 1635 nsew power bidirectional
rlabel metal4 s 156604 621040 157204 630400 6 vdda2
port 1636 nsew power bidirectional
rlabel metal4 s 120604 621040 121204 630400 6 vdda2
port 1637 nsew power bidirectional
rlabel metal4 s 48604 621040 49204 630400 6 vdda2
port 1638 nsew power bidirectional
rlabel metal4 s 552604 551680 553204 561040 6 vdda2
port 1639 nsew power bidirectional
rlabel metal4 s 516604 551680 517204 561040 6 vdda2
port 1640 nsew power bidirectional
rlabel metal4 s 480604 551680 481204 561040 6 vdda2
port 1641 nsew power bidirectional
rlabel metal4 s 408604 551680 409204 561040 6 vdda2
port 1642 nsew power bidirectional
rlabel metal4 s 372604 551680 373204 561040 6 vdda2
port 1643 nsew power bidirectional
rlabel metal4 s 336604 551680 337204 561040 6 vdda2
port 1644 nsew power bidirectional
rlabel metal4 s 300604 551680 301204 561040 6 vdda2
port 1645 nsew power bidirectional
rlabel metal4 s 264604 551680 265204 561040 6 vdda2
port 1646 nsew power bidirectional
rlabel metal4 s 228604 551680 229204 561040 6 vdda2
port 1647 nsew power bidirectional
rlabel metal4 s 192604 551680 193204 561040 6 vdda2
port 1648 nsew power bidirectional
rlabel metal4 s 156604 551680 157204 561040 6 vdda2
port 1649 nsew power bidirectional
rlabel metal4 s 120604 551680 121204 561040 6 vdda2
port 1650 nsew power bidirectional
rlabel metal4 s 48604 551680 49204 561040 6 vdda2
port 1651 nsew power bidirectional
rlabel metal4 s 552604 482320 553204 491680 6 vdda2
port 1652 nsew power bidirectional
rlabel metal4 s 516604 482320 517204 491680 6 vdda2
port 1653 nsew power bidirectional
rlabel metal4 s 480604 482320 481204 491680 6 vdda2
port 1654 nsew power bidirectional
rlabel metal4 s 408604 482320 409204 491680 6 vdda2
port 1655 nsew power bidirectional
rlabel metal4 s 372604 482320 373204 491680 6 vdda2
port 1656 nsew power bidirectional
rlabel metal4 s 336604 482320 337204 491680 6 vdda2
port 1657 nsew power bidirectional
rlabel metal4 s 300604 482320 301204 491680 6 vdda2
port 1658 nsew power bidirectional
rlabel metal4 s 264604 482320 265204 491680 6 vdda2
port 1659 nsew power bidirectional
rlabel metal4 s 228604 482320 229204 491680 6 vdda2
port 1660 nsew power bidirectional
rlabel metal4 s 192604 482320 193204 491680 6 vdda2
port 1661 nsew power bidirectional
rlabel metal4 s 156604 482320 157204 491680 6 vdda2
port 1662 nsew power bidirectional
rlabel metal4 s 120604 482320 121204 491680 6 vdda2
port 1663 nsew power bidirectional
rlabel metal4 s 48604 482320 49204 491680 6 vdda2
port 1664 nsew power bidirectional
rlabel metal4 s 552604 412960 553204 422320 6 vdda2
port 1665 nsew power bidirectional
rlabel metal4 s 516604 412960 517204 422320 6 vdda2
port 1666 nsew power bidirectional
rlabel metal4 s 480604 412960 481204 422320 6 vdda2
port 1667 nsew power bidirectional
rlabel metal4 s 408604 412960 409204 422320 6 vdda2
port 1668 nsew power bidirectional
rlabel metal4 s 372604 412960 373204 422320 6 vdda2
port 1669 nsew power bidirectional
rlabel metal4 s 336604 412960 337204 422320 6 vdda2
port 1670 nsew power bidirectional
rlabel metal4 s 300604 412960 301204 422320 6 vdda2
port 1671 nsew power bidirectional
rlabel metal4 s 264604 412960 265204 422320 6 vdda2
port 1672 nsew power bidirectional
rlabel metal4 s 228604 412960 229204 422320 6 vdda2
port 1673 nsew power bidirectional
rlabel metal4 s 192604 412960 193204 422320 6 vdda2
port 1674 nsew power bidirectional
rlabel metal4 s 156604 412960 157204 422320 6 vdda2
port 1675 nsew power bidirectional
rlabel metal4 s 120604 412960 121204 422320 6 vdda2
port 1676 nsew power bidirectional
rlabel metal4 s 48604 412960 49204 422320 6 vdda2
port 1677 nsew power bidirectional
rlabel metal4 s 552604 343600 553204 352960 6 vdda2
port 1678 nsew power bidirectional
rlabel metal4 s 516604 343600 517204 352960 6 vdda2
port 1679 nsew power bidirectional
rlabel metal4 s 480604 343600 481204 352960 6 vdda2
port 1680 nsew power bidirectional
rlabel metal4 s 408604 343600 409204 352960 6 vdda2
port 1681 nsew power bidirectional
rlabel metal4 s 372604 343600 373204 352960 6 vdda2
port 1682 nsew power bidirectional
rlabel metal4 s 336604 343600 337204 352960 6 vdda2
port 1683 nsew power bidirectional
rlabel metal4 s 300604 343600 301204 352960 6 vdda2
port 1684 nsew power bidirectional
rlabel metal4 s 264604 343600 265204 352960 6 vdda2
port 1685 nsew power bidirectional
rlabel metal4 s 228604 343600 229204 352960 6 vdda2
port 1686 nsew power bidirectional
rlabel metal4 s 192604 343600 193204 352960 6 vdda2
port 1687 nsew power bidirectional
rlabel metal4 s 156604 343600 157204 352960 6 vdda2
port 1688 nsew power bidirectional
rlabel metal4 s 120604 343600 121204 352960 6 vdda2
port 1689 nsew power bidirectional
rlabel metal4 s 48604 343600 49204 352960 6 vdda2
port 1690 nsew power bidirectional
rlabel metal4 s 552604 274240 553204 283600 6 vdda2
port 1691 nsew power bidirectional
rlabel metal4 s 516604 274240 517204 283600 6 vdda2
port 1692 nsew power bidirectional
rlabel metal4 s 480604 274240 481204 283600 6 vdda2
port 1693 nsew power bidirectional
rlabel metal4 s 408604 274240 409204 283600 6 vdda2
port 1694 nsew power bidirectional
rlabel metal4 s 372604 274240 373204 283600 6 vdda2
port 1695 nsew power bidirectional
rlabel metal4 s 336604 274240 337204 283600 6 vdda2
port 1696 nsew power bidirectional
rlabel metal4 s 300604 274240 301204 283600 6 vdda2
port 1697 nsew power bidirectional
rlabel metal4 s 264604 274240 265204 283600 6 vdda2
port 1698 nsew power bidirectional
rlabel metal4 s 228604 274240 229204 283600 6 vdda2
port 1699 nsew power bidirectional
rlabel metal4 s 192604 274240 193204 283600 6 vdda2
port 1700 nsew power bidirectional
rlabel metal4 s 156604 274240 157204 283600 6 vdda2
port 1701 nsew power bidirectional
rlabel metal4 s 120604 274240 121204 283600 6 vdda2
port 1702 nsew power bidirectional
rlabel metal4 s 48604 274240 49204 283600 6 vdda2
port 1703 nsew power bidirectional
rlabel metal4 s 552604 204880 553204 214240 6 vdda2
port 1704 nsew power bidirectional
rlabel metal4 s 516604 204880 517204 214240 6 vdda2
port 1705 nsew power bidirectional
rlabel metal4 s 480604 204880 481204 214240 6 vdda2
port 1706 nsew power bidirectional
rlabel metal4 s 408604 204880 409204 214240 6 vdda2
port 1707 nsew power bidirectional
rlabel metal4 s 372604 204880 373204 214240 6 vdda2
port 1708 nsew power bidirectional
rlabel metal4 s 336604 204880 337204 214240 6 vdda2
port 1709 nsew power bidirectional
rlabel metal4 s 300604 204880 301204 214240 6 vdda2
port 1710 nsew power bidirectional
rlabel metal4 s 264604 204880 265204 214240 6 vdda2
port 1711 nsew power bidirectional
rlabel metal4 s 228604 204880 229204 214240 6 vdda2
port 1712 nsew power bidirectional
rlabel metal4 s 192604 204880 193204 214240 6 vdda2
port 1713 nsew power bidirectional
rlabel metal4 s 156604 204880 157204 214240 6 vdda2
port 1714 nsew power bidirectional
rlabel metal4 s 120604 204880 121204 214240 6 vdda2
port 1715 nsew power bidirectional
rlabel metal4 s 48604 204880 49204 214240 6 vdda2
port 1716 nsew power bidirectional
rlabel metal4 s 552604 132200 553204 144880 6 vdda2
port 1717 nsew power bidirectional
rlabel metal4 s 516604 132200 517204 144880 6 vdda2
port 1718 nsew power bidirectional
rlabel metal4 s 480604 132200 481204 144880 6 vdda2
port 1719 nsew power bidirectional
rlabel metal4 s 408604 132200 409204 144880 6 vdda2
port 1720 nsew power bidirectional
rlabel metal4 s 372604 132200 373204 144880 6 vdda2
port 1721 nsew power bidirectional
rlabel metal4 s 336604 132200 337204 144880 6 vdda2
port 1722 nsew power bidirectional
rlabel metal4 s 300604 132200 301204 144880 6 vdda2
port 1723 nsew power bidirectional
rlabel metal4 s 264604 132200 265204 144880 6 vdda2
port 1724 nsew power bidirectional
rlabel metal4 s 228604 132200 229204 144880 6 vdda2
port 1725 nsew power bidirectional
rlabel metal4 s 192604 132200 193204 144880 6 vdda2
port 1726 nsew power bidirectional
rlabel metal4 s 156604 132200 157204 144880 6 vdda2
port 1727 nsew power bidirectional
rlabel metal4 s 120604 132200 121204 144880 6 vdda2
port 1728 nsew power bidirectional
rlabel metal4 s 48604 132200 49204 144880 6 vdda2
port 1729 nsew power bidirectional
rlabel metal4 s 552604 -7504 553204 8200 6 vdda2
port 1730 nsew power bidirectional
rlabel metal4 s 516604 -7504 517204 8200 6 vdda2
port 1731 nsew power bidirectional
rlabel metal4 s 480604 -7504 481204 8200 6 vdda2
port 1732 nsew power bidirectional
rlabel metal4 s 444604 -7504 445204 8200 6 vdda2
port 1733 nsew power bidirectional
rlabel metal4 s 408604 -7504 409204 8200 6 vdda2
port 1734 nsew power bidirectional
rlabel metal4 s 372604 -7504 373204 8200 6 vdda2
port 1735 nsew power bidirectional
rlabel metal4 s 336604 -7504 337204 8200 6 vdda2
port 1736 nsew power bidirectional
rlabel metal4 s 300604 -7504 301204 8200 6 vdda2
port 1737 nsew power bidirectional
rlabel metal4 s 264604 -7504 265204 8200 6 vdda2
port 1738 nsew power bidirectional
rlabel metal4 s 228604 -7504 229204 8200 6 vdda2
port 1739 nsew power bidirectional
rlabel metal4 s 192604 -7504 193204 8200 6 vdda2
port 1740 nsew power bidirectional
rlabel metal4 s 156604 -7504 157204 8200 6 vdda2
port 1741 nsew power bidirectional
rlabel metal4 s 120604 -7504 121204 8200 6 vdda2
port 1742 nsew power bidirectional
rlabel metal4 s 48604 -7504 49204 8200 6 vdda2
port 1743 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1744 nsew power bidirectional
rlabel metal5 s -8576 697676 592500 698276 6 vdda2
port 1745 nsew power bidirectional
rlabel metal5 s -8576 661676 592500 662276 6 vdda2
port 1746 nsew power bidirectional
rlabel metal5 s -8576 625676 592500 626276 6 vdda2
port 1747 nsew power bidirectional
rlabel metal5 s -8576 589676 592500 590276 6 vdda2
port 1748 nsew power bidirectional
rlabel metal5 s -8576 553676 592500 554276 6 vdda2
port 1749 nsew power bidirectional
rlabel metal5 s -8576 517676 592500 518276 6 vdda2
port 1750 nsew power bidirectional
rlabel metal5 s -8576 481676 592500 482276 6 vdda2
port 1751 nsew power bidirectional
rlabel metal5 s -8576 445676 592500 446276 6 vdda2
port 1752 nsew power bidirectional
rlabel metal5 s -8576 409676 592500 410276 6 vdda2
port 1753 nsew power bidirectional
rlabel metal5 s -8576 373676 592500 374276 6 vdda2
port 1754 nsew power bidirectional
rlabel metal5 s -8576 337676 592500 338276 6 vdda2
port 1755 nsew power bidirectional
rlabel metal5 s -8576 301676 592500 302276 6 vdda2
port 1756 nsew power bidirectional
rlabel metal5 s -8576 265676 592500 266276 6 vdda2
port 1757 nsew power bidirectional
rlabel metal5 s -8576 229676 592500 230276 6 vdda2
port 1758 nsew power bidirectional
rlabel metal5 s -8576 193676 592500 194276 6 vdda2
port 1759 nsew power bidirectional
rlabel metal5 s -8576 157676 592500 158276 6 vdda2
port 1760 nsew power bidirectional
rlabel metal5 s -8576 121676 592500 122276 6 vdda2
port 1761 nsew power bidirectional
rlabel metal5 s -8576 85676 592500 86276 6 vdda2
port 1762 nsew power bidirectional
rlabel metal5 s -8576 49676 592500 50276 6 vdda2
port 1763 nsew power bidirectional
rlabel metal5 s -8576 13676 592500 14276 6 vdda2
port 1764 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1765 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1766 nsew ground bidirectional
rlabel metal4 s 570604 690400 571204 711440 6 vssa2
port 1767 nsew ground bidirectional
rlabel metal4 s 534604 132200 535204 711440 6 vssa2
port 1768 nsew ground bidirectional
rlabel metal4 s 498604 690400 499204 711440 6 vssa2
port 1769 nsew ground bidirectional
rlabel metal4 s 462604 690400 463204 711440 6 vssa2
port 1770 nsew ground bidirectional
rlabel metal4 s 426604 690400 427204 711440 6 vssa2
port 1771 nsew ground bidirectional
rlabel metal4 s 390604 690400 391204 711440 6 vssa2
port 1772 nsew ground bidirectional
rlabel metal4 s 354604 690400 355204 711440 6 vssa2
port 1773 nsew ground bidirectional
rlabel metal4 s 318604 690400 319204 711440 6 vssa2
port 1774 nsew ground bidirectional
rlabel metal4 s 282604 690400 283204 711440 6 vssa2
port 1775 nsew ground bidirectional
rlabel metal4 s 246604 690400 247204 711440 6 vssa2
port 1776 nsew ground bidirectional
rlabel metal4 s 210604 690400 211204 711440 6 vssa2
port 1777 nsew ground bidirectional
rlabel metal4 s 174604 690400 175204 711440 6 vssa2
port 1778 nsew ground bidirectional
rlabel metal4 s 138604 132200 139204 711440 6 vssa2
port 1779 nsew ground bidirectional
rlabel metal4 s 102604 690400 103204 711440 6 vssa2
port 1780 nsew ground bidirectional
rlabel metal4 s 66604 690400 67204 711440 6 vssa2
port 1781 nsew ground bidirectional
rlabel metal4 s 30604 690400 31204 711440 6 vssa2
port 1782 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1783 nsew ground bidirectional
rlabel metal4 s 570604 621040 571204 630400 6 vssa2
port 1784 nsew ground bidirectional
rlabel metal4 s 498604 621040 499204 630400 6 vssa2
port 1785 nsew ground bidirectional
rlabel metal4 s 462604 621040 463204 630400 6 vssa2
port 1786 nsew ground bidirectional
rlabel metal4 s 426604 621040 427204 630400 6 vssa2
port 1787 nsew ground bidirectional
rlabel metal4 s 390604 621040 391204 630400 6 vssa2
port 1788 nsew ground bidirectional
rlabel metal4 s 354604 621040 355204 630400 6 vssa2
port 1789 nsew ground bidirectional
rlabel metal4 s 318604 621040 319204 630400 6 vssa2
port 1790 nsew ground bidirectional
rlabel metal4 s 282604 621040 283204 630400 6 vssa2
port 1791 nsew ground bidirectional
rlabel metal4 s 246604 621040 247204 630400 6 vssa2
port 1792 nsew ground bidirectional
rlabel metal4 s 210604 621040 211204 630400 6 vssa2
port 1793 nsew ground bidirectional
rlabel metal4 s 174604 621040 175204 630400 6 vssa2
port 1794 nsew ground bidirectional
rlabel metal4 s 102604 621040 103204 630400 6 vssa2
port 1795 nsew ground bidirectional
rlabel metal4 s 66604 621040 67204 630400 6 vssa2
port 1796 nsew ground bidirectional
rlabel metal4 s 30604 621040 31204 630400 6 vssa2
port 1797 nsew ground bidirectional
rlabel metal4 s 570604 551680 571204 561040 6 vssa2
port 1798 nsew ground bidirectional
rlabel metal4 s 498604 551680 499204 561040 6 vssa2
port 1799 nsew ground bidirectional
rlabel metal4 s 462604 551680 463204 561040 6 vssa2
port 1800 nsew ground bidirectional
rlabel metal4 s 426604 551680 427204 561040 6 vssa2
port 1801 nsew ground bidirectional
rlabel metal4 s 390604 551680 391204 561040 6 vssa2
port 1802 nsew ground bidirectional
rlabel metal4 s 354604 551680 355204 561040 6 vssa2
port 1803 nsew ground bidirectional
rlabel metal4 s 318604 551680 319204 561040 6 vssa2
port 1804 nsew ground bidirectional
rlabel metal4 s 282604 551680 283204 561040 6 vssa2
port 1805 nsew ground bidirectional
rlabel metal4 s 246604 551680 247204 561040 6 vssa2
port 1806 nsew ground bidirectional
rlabel metal4 s 210604 551680 211204 561040 6 vssa2
port 1807 nsew ground bidirectional
rlabel metal4 s 174604 551680 175204 561040 6 vssa2
port 1808 nsew ground bidirectional
rlabel metal4 s 102604 551680 103204 561040 6 vssa2
port 1809 nsew ground bidirectional
rlabel metal4 s 66604 551680 67204 561040 6 vssa2
port 1810 nsew ground bidirectional
rlabel metal4 s 30604 551680 31204 561040 6 vssa2
port 1811 nsew ground bidirectional
rlabel metal4 s 570604 482320 571204 491680 6 vssa2
port 1812 nsew ground bidirectional
rlabel metal4 s 498604 482320 499204 491680 6 vssa2
port 1813 nsew ground bidirectional
rlabel metal4 s 462604 482320 463204 491680 6 vssa2
port 1814 nsew ground bidirectional
rlabel metal4 s 426604 482320 427204 491680 6 vssa2
port 1815 nsew ground bidirectional
rlabel metal4 s 390604 482320 391204 491680 6 vssa2
port 1816 nsew ground bidirectional
rlabel metal4 s 354604 482320 355204 491680 6 vssa2
port 1817 nsew ground bidirectional
rlabel metal4 s 318604 482320 319204 491680 6 vssa2
port 1818 nsew ground bidirectional
rlabel metal4 s 282604 482320 283204 491680 6 vssa2
port 1819 nsew ground bidirectional
rlabel metal4 s 246604 482320 247204 491680 6 vssa2
port 1820 nsew ground bidirectional
rlabel metal4 s 210604 482320 211204 491680 6 vssa2
port 1821 nsew ground bidirectional
rlabel metal4 s 174604 482320 175204 491680 6 vssa2
port 1822 nsew ground bidirectional
rlabel metal4 s 102604 482320 103204 491680 6 vssa2
port 1823 nsew ground bidirectional
rlabel metal4 s 66604 482320 67204 491680 6 vssa2
port 1824 nsew ground bidirectional
rlabel metal4 s 30604 482320 31204 491680 6 vssa2
port 1825 nsew ground bidirectional
rlabel metal4 s 570604 412960 571204 422320 6 vssa2
port 1826 nsew ground bidirectional
rlabel metal4 s 498604 412960 499204 422320 6 vssa2
port 1827 nsew ground bidirectional
rlabel metal4 s 462604 412960 463204 422320 6 vssa2
port 1828 nsew ground bidirectional
rlabel metal4 s 426604 412960 427204 422320 6 vssa2
port 1829 nsew ground bidirectional
rlabel metal4 s 390604 412960 391204 422320 6 vssa2
port 1830 nsew ground bidirectional
rlabel metal4 s 354604 412960 355204 422320 6 vssa2
port 1831 nsew ground bidirectional
rlabel metal4 s 318604 412960 319204 422320 6 vssa2
port 1832 nsew ground bidirectional
rlabel metal4 s 282604 412960 283204 422320 6 vssa2
port 1833 nsew ground bidirectional
rlabel metal4 s 246604 412960 247204 422320 6 vssa2
port 1834 nsew ground bidirectional
rlabel metal4 s 210604 412960 211204 422320 6 vssa2
port 1835 nsew ground bidirectional
rlabel metal4 s 174604 412960 175204 422320 6 vssa2
port 1836 nsew ground bidirectional
rlabel metal4 s 102604 412960 103204 422320 6 vssa2
port 1837 nsew ground bidirectional
rlabel metal4 s 66604 412960 67204 422320 6 vssa2
port 1838 nsew ground bidirectional
rlabel metal4 s 30604 412960 31204 422320 6 vssa2
port 1839 nsew ground bidirectional
rlabel metal4 s 570604 343600 571204 352960 6 vssa2
port 1840 nsew ground bidirectional
rlabel metal4 s 498604 343600 499204 352960 6 vssa2
port 1841 nsew ground bidirectional
rlabel metal4 s 462604 343600 463204 352960 6 vssa2
port 1842 nsew ground bidirectional
rlabel metal4 s 426604 343600 427204 352960 6 vssa2
port 1843 nsew ground bidirectional
rlabel metal4 s 390604 343600 391204 352960 6 vssa2
port 1844 nsew ground bidirectional
rlabel metal4 s 354604 343600 355204 352960 6 vssa2
port 1845 nsew ground bidirectional
rlabel metal4 s 318604 343600 319204 352960 6 vssa2
port 1846 nsew ground bidirectional
rlabel metal4 s 282604 343600 283204 352960 6 vssa2
port 1847 nsew ground bidirectional
rlabel metal4 s 246604 343600 247204 352960 6 vssa2
port 1848 nsew ground bidirectional
rlabel metal4 s 210604 343600 211204 352960 6 vssa2
port 1849 nsew ground bidirectional
rlabel metal4 s 174604 343600 175204 352960 6 vssa2
port 1850 nsew ground bidirectional
rlabel metal4 s 102604 343600 103204 352960 6 vssa2
port 1851 nsew ground bidirectional
rlabel metal4 s 66604 343600 67204 352960 6 vssa2
port 1852 nsew ground bidirectional
rlabel metal4 s 30604 343600 31204 352960 6 vssa2
port 1853 nsew ground bidirectional
rlabel metal4 s 570604 274240 571204 283600 6 vssa2
port 1854 nsew ground bidirectional
rlabel metal4 s 498604 274240 499204 283600 6 vssa2
port 1855 nsew ground bidirectional
rlabel metal4 s 462604 274240 463204 283600 6 vssa2
port 1856 nsew ground bidirectional
rlabel metal4 s 426604 274240 427204 283600 6 vssa2
port 1857 nsew ground bidirectional
rlabel metal4 s 390604 274240 391204 283600 6 vssa2
port 1858 nsew ground bidirectional
rlabel metal4 s 354604 274240 355204 283600 6 vssa2
port 1859 nsew ground bidirectional
rlabel metal4 s 318604 274240 319204 283600 6 vssa2
port 1860 nsew ground bidirectional
rlabel metal4 s 282604 274240 283204 283600 6 vssa2
port 1861 nsew ground bidirectional
rlabel metal4 s 246604 274240 247204 283600 6 vssa2
port 1862 nsew ground bidirectional
rlabel metal4 s 210604 274240 211204 283600 6 vssa2
port 1863 nsew ground bidirectional
rlabel metal4 s 174604 274240 175204 283600 6 vssa2
port 1864 nsew ground bidirectional
rlabel metal4 s 102604 274240 103204 283600 6 vssa2
port 1865 nsew ground bidirectional
rlabel metal4 s 66604 274240 67204 283600 6 vssa2
port 1866 nsew ground bidirectional
rlabel metal4 s 30604 274240 31204 283600 6 vssa2
port 1867 nsew ground bidirectional
rlabel metal4 s 570604 204880 571204 214240 6 vssa2
port 1868 nsew ground bidirectional
rlabel metal4 s 498604 204880 499204 214240 6 vssa2
port 1869 nsew ground bidirectional
rlabel metal4 s 462604 204880 463204 214240 6 vssa2
port 1870 nsew ground bidirectional
rlabel metal4 s 426604 204880 427204 214240 6 vssa2
port 1871 nsew ground bidirectional
rlabel metal4 s 390604 204880 391204 214240 6 vssa2
port 1872 nsew ground bidirectional
rlabel metal4 s 354604 204880 355204 214240 6 vssa2
port 1873 nsew ground bidirectional
rlabel metal4 s 318604 204880 319204 214240 6 vssa2
port 1874 nsew ground bidirectional
rlabel metal4 s 282604 204880 283204 214240 6 vssa2
port 1875 nsew ground bidirectional
rlabel metal4 s 246604 204880 247204 214240 6 vssa2
port 1876 nsew ground bidirectional
rlabel metal4 s 210604 204880 211204 214240 6 vssa2
port 1877 nsew ground bidirectional
rlabel metal4 s 174604 204880 175204 214240 6 vssa2
port 1878 nsew ground bidirectional
rlabel metal4 s 102604 204880 103204 214240 6 vssa2
port 1879 nsew ground bidirectional
rlabel metal4 s 66604 204880 67204 214240 6 vssa2
port 1880 nsew ground bidirectional
rlabel metal4 s 30604 204880 31204 214240 6 vssa2
port 1881 nsew ground bidirectional
rlabel metal4 s 570604 -7504 571204 144880 6 vssa2
port 1882 nsew ground bidirectional
rlabel metal4 s 498604 132200 499204 144880 6 vssa2
port 1883 nsew ground bidirectional
rlabel metal4 s 462604 132200 463204 144880 6 vssa2
port 1884 nsew ground bidirectional
rlabel metal4 s 426604 132200 427204 144880 6 vssa2
port 1885 nsew ground bidirectional
rlabel metal4 s 390604 132200 391204 144880 6 vssa2
port 1886 nsew ground bidirectional
rlabel metal4 s 354604 132200 355204 144880 6 vssa2
port 1887 nsew ground bidirectional
rlabel metal4 s 318604 132200 319204 144880 6 vssa2
port 1888 nsew ground bidirectional
rlabel metal4 s 282604 132200 283204 144880 6 vssa2
port 1889 nsew ground bidirectional
rlabel metal4 s 246604 132200 247204 144880 6 vssa2
port 1890 nsew ground bidirectional
rlabel metal4 s 210604 132200 211204 144880 6 vssa2
port 1891 nsew ground bidirectional
rlabel metal4 s 174604 132200 175204 144880 6 vssa2
port 1892 nsew ground bidirectional
rlabel metal4 s 102604 132200 103204 144880 6 vssa2
port 1893 nsew ground bidirectional
rlabel metal4 s 66604 132200 67204 144880 6 vssa2
port 1894 nsew ground bidirectional
rlabel metal4 s 30604 -7504 31204 144880 6 vssa2
port 1895 nsew ground bidirectional
rlabel metal4 s 534604 -7504 535204 8200 6 vssa2
port 1896 nsew ground bidirectional
rlabel metal4 s 498604 -7504 499204 8200 6 vssa2
port 1897 nsew ground bidirectional
rlabel metal4 s 462604 -7504 463204 8200 6 vssa2
port 1898 nsew ground bidirectional
rlabel metal4 s 426604 -7504 427204 8200 6 vssa2
port 1899 nsew ground bidirectional
rlabel metal4 s 390604 -7504 391204 8200 6 vssa2
port 1900 nsew ground bidirectional
rlabel metal4 s 354604 -7504 355204 8200 6 vssa2
port 1901 nsew ground bidirectional
rlabel metal4 s 318604 -7504 319204 8200 6 vssa2
port 1902 nsew ground bidirectional
rlabel metal4 s 282604 -7504 283204 8200 6 vssa2
port 1903 nsew ground bidirectional
rlabel metal4 s 246604 -7504 247204 8200 6 vssa2
port 1904 nsew ground bidirectional
rlabel metal4 s 210604 -7504 211204 8200 6 vssa2
port 1905 nsew ground bidirectional
rlabel metal4 s 174604 -7504 175204 8200 6 vssa2
port 1906 nsew ground bidirectional
rlabel metal4 s 138604 -7504 139204 8200 6 vssa2
port 1907 nsew ground bidirectional
rlabel metal4 s 102604 -7504 103204 8200 6 vssa2
port 1908 nsew ground bidirectional
rlabel metal4 s 66604 -7504 67204 8200 6 vssa2
port 1909 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1910 nsew ground bidirectional
rlabel metal5 s -8576 679676 592500 680276 6 vssa2
port 1911 nsew ground bidirectional
rlabel metal5 s -8576 643676 592500 644276 6 vssa2
port 1912 nsew ground bidirectional
rlabel metal5 s -8576 607676 592500 608276 6 vssa2
port 1913 nsew ground bidirectional
rlabel metal5 s -8576 571676 592500 572276 6 vssa2
port 1914 nsew ground bidirectional
rlabel metal5 s -8576 535676 592500 536276 6 vssa2
port 1915 nsew ground bidirectional
rlabel metal5 s -8576 499676 592500 500276 6 vssa2
port 1916 nsew ground bidirectional
rlabel metal5 s -8576 463676 592500 464276 6 vssa2
port 1917 nsew ground bidirectional
rlabel metal5 s -8576 427676 592500 428276 6 vssa2
port 1918 nsew ground bidirectional
rlabel metal5 s -8576 391676 592500 392276 6 vssa2
port 1919 nsew ground bidirectional
rlabel metal5 s -8576 355676 592500 356276 6 vssa2
port 1920 nsew ground bidirectional
rlabel metal5 s -8576 319676 592500 320276 6 vssa2
port 1921 nsew ground bidirectional
rlabel metal5 s -8576 283676 592500 284276 6 vssa2
port 1922 nsew ground bidirectional
rlabel metal5 s -8576 247676 592500 248276 6 vssa2
port 1923 nsew ground bidirectional
rlabel metal5 s -8576 211676 592500 212276 6 vssa2
port 1924 nsew ground bidirectional
rlabel metal5 s -8576 175676 592500 176276 6 vssa2
port 1925 nsew ground bidirectional
rlabel metal5 s -8576 139676 592500 140276 6 vssa2
port 1926 nsew ground bidirectional
rlabel metal5 s -8576 103676 592500 104276 6 vssa2
port 1927 nsew ground bidirectional
rlabel metal5 s -8576 67676 592500 68276 6 vssa2
port 1928 nsew ground bidirectional
rlabel metal5 s -8576 31676 592500 32276 6 vssa2
port 1929 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1930 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 584000 704000
string LEFview TRUE
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 104687420
string GDS_START 66671208
<< end >>

