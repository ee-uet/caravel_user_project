magic
tech sky130A
magscale 1 2
timestamp 1624054018
<< obsli1 >>
rect 1104 2159 38979 117521
<< obsm1 >>
rect 106 1436 39914 117972
<< metal2 >>
rect 110 119200 166 120800
rect 294 119200 350 120800
rect 478 119200 534 120800
rect 662 119200 718 120800
rect 938 119200 994 120800
rect 1122 119200 1178 120800
rect 1306 119200 1362 120800
rect 1582 119200 1638 120800
rect 1766 119200 1822 120800
rect 1950 119200 2006 120800
rect 2226 119200 2282 120800
rect 2410 119200 2466 120800
rect 2594 119200 2650 120800
rect 2778 119200 2834 120800
rect 3054 119200 3110 120800
rect 3238 119200 3294 120800
rect 3422 119200 3478 120800
rect 3698 119200 3754 120800
rect 3882 119200 3938 120800
rect 4066 119200 4122 120800
rect 4342 119200 4398 120800
rect 4526 119200 4582 120800
rect 4710 119200 4766 120800
rect 4894 119200 4950 120800
rect 5170 119200 5226 120800
rect 5354 119200 5410 120800
rect 5538 119200 5594 120800
rect 5814 119200 5870 120800
rect 5998 119200 6054 120800
rect 6182 119200 6238 120800
rect 6458 119200 6514 120800
rect 6642 119200 6698 120800
rect 6826 119200 6882 120800
rect 7010 119200 7066 120800
rect 7286 119200 7342 120800
rect 7470 119200 7526 120800
rect 7654 119200 7710 120800
rect 7930 119200 7986 120800
rect 8114 119200 8170 120800
rect 8298 119200 8354 120800
rect 8574 119200 8630 120800
rect 8758 119200 8814 120800
rect 8942 119200 8998 120800
rect 9126 119200 9182 120800
rect 9402 119200 9458 120800
rect 9586 119200 9642 120800
rect 9770 119200 9826 120800
rect 10046 119200 10102 120800
rect 10230 119200 10286 120800
rect 10414 119200 10470 120800
rect 10690 119200 10746 120800
rect 10874 119200 10930 120800
rect 11058 119200 11114 120800
rect 11242 119200 11298 120800
rect 11518 119200 11574 120800
rect 11702 119200 11758 120800
rect 11886 119200 11942 120800
rect 12162 119200 12218 120800
rect 12346 119200 12402 120800
rect 12530 119200 12586 120800
rect 12806 119200 12862 120800
rect 12990 119200 13046 120800
rect 13174 119200 13230 120800
rect 13450 119200 13506 120800
rect 13634 119200 13690 120800
rect 13818 119200 13874 120800
rect 14002 119200 14058 120800
rect 14278 119200 14334 120800
rect 14462 119200 14518 120800
rect 14646 119200 14702 120800
rect 14922 119200 14978 120800
rect 15106 119200 15162 120800
rect 15290 119200 15346 120800
rect 15566 119200 15622 120800
rect 15750 119200 15806 120800
rect 15934 119200 15990 120800
rect 16118 119200 16174 120800
rect 16394 119200 16450 120800
rect 16578 119200 16634 120800
rect 16762 119200 16818 120800
rect 17038 119200 17094 120800
rect 17222 119200 17278 120800
rect 17406 119200 17462 120800
rect 17682 119200 17738 120800
rect 17866 119200 17922 120800
rect 18050 119200 18106 120800
rect 18234 119200 18290 120800
rect 18510 119200 18566 120800
rect 18694 119200 18750 120800
rect 18878 119200 18934 120800
rect 19154 119200 19210 120800
rect 19338 119200 19394 120800
rect 19522 119200 19578 120800
rect 19798 119200 19854 120800
rect 19982 119200 20038 120800
rect 20166 119200 20222 120800
rect 20350 119200 20406 120800
rect 20626 119200 20682 120800
rect 20810 119200 20866 120800
rect 20994 119200 21050 120800
rect 21270 119200 21326 120800
rect 21454 119200 21510 120800
rect 21638 119200 21694 120800
rect 21914 119200 21970 120800
rect 22098 119200 22154 120800
rect 22282 119200 22338 120800
rect 22466 119200 22522 120800
rect 22742 119200 22798 120800
rect 22926 119200 22982 120800
rect 23110 119200 23166 120800
rect 23386 119200 23442 120800
rect 23570 119200 23626 120800
rect 23754 119200 23810 120800
rect 24030 119200 24086 120800
rect 24214 119200 24270 120800
rect 24398 119200 24454 120800
rect 24582 119200 24638 120800
rect 24858 119200 24914 120800
rect 25042 119200 25098 120800
rect 25226 119200 25282 120800
rect 25502 119200 25558 120800
rect 25686 119200 25742 120800
rect 25870 119200 25926 120800
rect 26146 119200 26202 120800
rect 26330 119200 26386 120800
rect 26514 119200 26570 120800
rect 26790 119200 26846 120800
rect 26974 119200 27030 120800
rect 27158 119200 27214 120800
rect 27342 119200 27398 120800
rect 27618 119200 27674 120800
rect 27802 119200 27858 120800
rect 27986 119200 28042 120800
rect 28262 119200 28318 120800
rect 28446 119200 28502 120800
rect 28630 119200 28686 120800
rect 28906 119200 28962 120800
rect 29090 119200 29146 120800
rect 29274 119200 29330 120800
rect 29458 119200 29514 120800
rect 29734 119200 29790 120800
rect 29918 119200 29974 120800
rect 30102 119200 30158 120800
rect 30378 119200 30434 120800
rect 30562 119200 30618 120800
rect 30746 119200 30802 120800
rect 31022 119200 31078 120800
rect 31206 119200 31262 120800
rect 31390 119200 31446 120800
rect 31574 119200 31630 120800
rect 31850 119200 31906 120800
rect 32034 119200 32090 120800
rect 32218 119200 32274 120800
rect 32494 119200 32550 120800
rect 32678 119200 32734 120800
rect 32862 119200 32918 120800
rect 33138 119200 33194 120800
rect 33322 119200 33378 120800
rect 33506 119200 33562 120800
rect 33690 119200 33746 120800
rect 33966 119200 34022 120800
rect 34150 119200 34206 120800
rect 34334 119200 34390 120800
rect 34610 119200 34666 120800
rect 34794 119200 34850 120800
rect 34978 119200 35034 120800
rect 35254 119200 35310 120800
rect 35438 119200 35494 120800
rect 35622 119200 35678 120800
rect 35806 119200 35862 120800
rect 36082 119200 36138 120800
rect 36266 119200 36322 120800
rect 36450 119200 36506 120800
rect 36726 119200 36782 120800
rect 36910 119200 36966 120800
rect 37094 119200 37150 120800
rect 37370 119200 37426 120800
rect 37554 119200 37610 120800
rect 37738 119200 37794 120800
rect 37922 119200 37978 120800
rect 38198 119200 38254 120800
rect 38382 119200 38438 120800
rect 38566 119200 38622 120800
rect 38842 119200 38898 120800
rect 39026 119200 39082 120800
rect 39210 119200 39266 120800
rect 39486 119200 39542 120800
rect 39670 119200 39726 120800
rect 39854 119200 39910 120800
rect 110 -800 166 800
rect 386 -800 442 800
rect 662 -800 718 800
rect 938 -800 994 800
rect 1214 -800 1270 800
rect 1490 -800 1546 800
rect 1858 -800 1914 800
rect 2134 -800 2190 800
rect 2410 -800 2466 800
rect 2686 -800 2742 800
rect 2962 -800 3018 800
rect 3238 -800 3294 800
rect 3606 -800 3662 800
rect 3882 -800 3938 800
rect 4158 -800 4214 800
rect 4434 -800 4490 800
rect 4710 -800 4766 800
rect 4986 -800 5042 800
rect 5354 -800 5410 800
rect 5630 -800 5686 800
rect 5906 -800 5962 800
rect 6182 -800 6238 800
rect 6458 -800 6514 800
rect 6826 -800 6882 800
rect 7102 -800 7158 800
rect 7378 -800 7434 800
rect 7654 -800 7710 800
rect 7930 -800 7986 800
rect 8206 -800 8262 800
rect 8574 -800 8630 800
rect 8850 -800 8906 800
rect 9126 -800 9182 800
rect 9402 -800 9458 800
rect 9678 -800 9734 800
rect 9954 -800 10010 800
rect 10322 -800 10378 800
rect 10598 -800 10654 800
rect 10874 -800 10930 800
rect 11150 -800 11206 800
rect 11426 -800 11482 800
rect 11794 -800 11850 800
rect 12070 -800 12126 800
rect 12346 -800 12402 800
rect 12622 -800 12678 800
rect 12898 -800 12954 800
rect 13174 -800 13230 800
rect 13542 -800 13598 800
rect 13818 -800 13874 800
rect 14094 -800 14150 800
rect 14370 -800 14426 800
rect 14646 -800 14702 800
rect 14922 -800 14978 800
rect 15290 -800 15346 800
rect 15566 -800 15622 800
rect 15842 -800 15898 800
rect 16118 -800 16174 800
rect 16394 -800 16450 800
rect 16670 -800 16726 800
rect 17038 -800 17094 800
rect 17314 -800 17370 800
rect 17590 -800 17646 800
rect 17866 -800 17922 800
rect 18142 -800 18198 800
rect 18510 -800 18566 800
rect 18786 -800 18842 800
rect 19062 -800 19118 800
rect 19338 -800 19394 800
rect 19614 -800 19670 800
rect 19890 -800 19946 800
rect 20258 -800 20314 800
rect 20534 -800 20590 800
rect 20810 -800 20866 800
rect 21086 -800 21142 800
rect 21362 -800 21418 800
rect 21638 -800 21694 800
rect 22006 -800 22062 800
rect 22282 -800 22338 800
rect 22558 -800 22614 800
rect 22834 -800 22890 800
rect 23110 -800 23166 800
rect 23478 -800 23534 800
rect 23754 -800 23810 800
rect 24030 -800 24086 800
rect 24306 -800 24362 800
rect 24582 -800 24638 800
rect 24858 -800 24914 800
rect 25226 -800 25282 800
rect 25502 -800 25558 800
rect 25778 -800 25834 800
rect 26054 -800 26110 800
rect 26330 -800 26386 800
rect 26606 -800 26662 800
rect 26974 -800 27030 800
rect 27250 -800 27306 800
rect 27526 -800 27582 800
rect 27802 -800 27858 800
rect 28078 -800 28134 800
rect 28354 -800 28410 800
rect 28722 -800 28778 800
rect 28998 -800 29054 800
rect 29274 -800 29330 800
rect 29550 -800 29606 800
rect 29826 -800 29882 800
rect 30194 -800 30250 800
rect 30470 -800 30526 800
rect 30746 -800 30802 800
rect 31022 -800 31078 800
rect 31298 -800 31354 800
rect 31574 -800 31630 800
rect 31942 -800 31998 800
rect 32218 -800 32274 800
rect 32494 -800 32550 800
rect 32770 -800 32826 800
rect 33046 -800 33102 800
rect 33322 -800 33378 800
rect 33690 -800 33746 800
rect 33966 -800 34022 800
rect 34242 -800 34298 800
rect 34518 -800 34574 800
rect 34794 -800 34850 800
rect 35162 -800 35218 800
rect 35438 -800 35494 800
rect 35714 -800 35770 800
rect 35990 -800 36046 800
rect 36266 -800 36322 800
rect 36542 -800 36598 800
rect 36910 -800 36966 800
rect 37186 -800 37242 800
rect 37462 -800 37518 800
rect 37738 -800 37794 800
rect 38014 -800 38070 800
rect 38290 -800 38346 800
rect 38658 -800 38714 800
rect 38934 -800 38990 800
rect 39210 -800 39266 800
rect 39486 -800 39542 800
rect 39762 -800 39818 800
<< obsm2 >>
rect 222 119144 238 119649
rect 406 119144 422 119649
rect 590 119144 606 119649
rect 774 119144 882 119649
rect 1050 119144 1066 119649
rect 1234 119144 1250 119649
rect 1418 119144 1526 119649
rect 1694 119144 1710 119649
rect 1878 119144 1894 119649
rect 2062 119144 2170 119649
rect 2338 119144 2354 119649
rect 2522 119144 2538 119649
rect 2706 119144 2722 119649
rect 2890 119144 2998 119649
rect 3166 119144 3182 119649
rect 3350 119144 3366 119649
rect 3534 119144 3642 119649
rect 3810 119144 3826 119649
rect 3994 119144 4010 119649
rect 4178 119144 4286 119649
rect 4454 119144 4470 119649
rect 4638 119144 4654 119649
rect 4822 119144 4838 119649
rect 5006 119144 5114 119649
rect 5282 119144 5298 119649
rect 5466 119144 5482 119649
rect 5650 119144 5758 119649
rect 5926 119144 5942 119649
rect 6110 119144 6126 119649
rect 6294 119144 6402 119649
rect 6570 119144 6586 119649
rect 6754 119144 6770 119649
rect 6938 119144 6954 119649
rect 7122 119144 7230 119649
rect 7398 119144 7414 119649
rect 7582 119144 7598 119649
rect 7766 119144 7874 119649
rect 8042 119144 8058 119649
rect 8226 119144 8242 119649
rect 8410 119144 8518 119649
rect 8686 119144 8702 119649
rect 8870 119144 8886 119649
rect 9054 119144 9070 119649
rect 9238 119144 9346 119649
rect 9514 119144 9530 119649
rect 9698 119144 9714 119649
rect 9882 119144 9990 119649
rect 10158 119144 10174 119649
rect 10342 119144 10358 119649
rect 10526 119144 10634 119649
rect 10802 119144 10818 119649
rect 10986 119144 11002 119649
rect 11170 119144 11186 119649
rect 11354 119144 11462 119649
rect 11630 119144 11646 119649
rect 11814 119144 11830 119649
rect 11998 119144 12106 119649
rect 12274 119144 12290 119649
rect 12458 119144 12474 119649
rect 12642 119144 12750 119649
rect 12918 119144 12934 119649
rect 13102 119144 13118 119649
rect 13286 119144 13394 119649
rect 13562 119144 13578 119649
rect 13746 119144 13762 119649
rect 13930 119144 13946 119649
rect 14114 119144 14222 119649
rect 14390 119144 14406 119649
rect 14574 119144 14590 119649
rect 14758 119144 14866 119649
rect 15034 119144 15050 119649
rect 15218 119144 15234 119649
rect 15402 119144 15510 119649
rect 15678 119144 15694 119649
rect 15862 119144 15878 119649
rect 16046 119144 16062 119649
rect 16230 119144 16338 119649
rect 16506 119144 16522 119649
rect 16690 119144 16706 119649
rect 16874 119144 16982 119649
rect 17150 119144 17166 119649
rect 17334 119144 17350 119649
rect 17518 119144 17626 119649
rect 17794 119144 17810 119649
rect 17978 119144 17994 119649
rect 18162 119144 18178 119649
rect 18346 119144 18454 119649
rect 18622 119144 18638 119649
rect 18806 119144 18822 119649
rect 18990 119144 19098 119649
rect 19266 119144 19282 119649
rect 19450 119144 19466 119649
rect 19634 119144 19742 119649
rect 19910 119144 19926 119649
rect 20094 119144 20110 119649
rect 20278 119144 20294 119649
rect 20462 119144 20570 119649
rect 20738 119144 20754 119649
rect 20922 119144 20938 119649
rect 21106 119144 21214 119649
rect 21382 119144 21398 119649
rect 21566 119144 21582 119649
rect 21750 119144 21858 119649
rect 22026 119144 22042 119649
rect 22210 119144 22226 119649
rect 22394 119144 22410 119649
rect 22578 119144 22686 119649
rect 22854 119144 22870 119649
rect 23038 119144 23054 119649
rect 23222 119144 23330 119649
rect 23498 119144 23514 119649
rect 23682 119144 23698 119649
rect 23866 119144 23974 119649
rect 24142 119144 24158 119649
rect 24326 119144 24342 119649
rect 24510 119144 24526 119649
rect 24694 119144 24802 119649
rect 24970 119144 24986 119649
rect 25154 119144 25170 119649
rect 25338 119144 25446 119649
rect 25614 119144 25630 119649
rect 25798 119144 25814 119649
rect 25982 119144 26090 119649
rect 26258 119144 26274 119649
rect 26442 119144 26458 119649
rect 26626 119144 26734 119649
rect 26902 119144 26918 119649
rect 27086 119144 27102 119649
rect 27270 119144 27286 119649
rect 27454 119144 27562 119649
rect 27730 119144 27746 119649
rect 27914 119144 27930 119649
rect 28098 119144 28206 119649
rect 28374 119144 28390 119649
rect 28558 119144 28574 119649
rect 28742 119144 28850 119649
rect 29018 119144 29034 119649
rect 29202 119144 29218 119649
rect 29386 119144 29402 119649
rect 29570 119144 29678 119649
rect 29846 119144 29862 119649
rect 30030 119144 30046 119649
rect 30214 119144 30322 119649
rect 30490 119144 30506 119649
rect 30674 119144 30690 119649
rect 30858 119144 30966 119649
rect 31134 119144 31150 119649
rect 31318 119144 31334 119649
rect 31502 119144 31518 119649
rect 31686 119144 31794 119649
rect 31962 119144 31978 119649
rect 32146 119144 32162 119649
rect 32330 119144 32438 119649
rect 32606 119144 32622 119649
rect 32790 119144 32806 119649
rect 32974 119144 33082 119649
rect 33250 119144 33266 119649
rect 33434 119144 33450 119649
rect 33618 119144 33634 119649
rect 33802 119144 33910 119649
rect 34078 119144 34094 119649
rect 34262 119144 34278 119649
rect 34446 119144 34554 119649
rect 34722 119144 34738 119649
rect 34906 119144 34922 119649
rect 35090 119144 35198 119649
rect 35366 119144 35382 119649
rect 35550 119144 35566 119649
rect 35734 119144 35750 119649
rect 35918 119144 36026 119649
rect 36194 119144 36210 119649
rect 36378 119144 36394 119649
rect 36562 119144 36670 119649
rect 36838 119144 36854 119649
rect 37022 119144 37038 119649
rect 37206 119144 37314 119649
rect 37482 119144 37498 119649
rect 37666 119144 37682 119649
rect 37850 119144 37866 119649
rect 38034 119144 38142 119649
rect 38310 119144 38326 119649
rect 38494 119144 38510 119649
rect 38678 119144 38786 119649
rect 38954 119144 38970 119649
rect 39138 119144 39154 119649
rect 39322 119144 39430 119649
rect 39598 119144 39614 119649
rect 39782 119144 39798 119649
rect 112 856 39908 119144
rect 222 167 330 856
rect 498 167 606 856
rect 774 167 882 856
rect 1050 167 1158 856
rect 1326 167 1434 856
rect 1602 167 1802 856
rect 1970 167 2078 856
rect 2246 167 2354 856
rect 2522 167 2630 856
rect 2798 167 2906 856
rect 3074 167 3182 856
rect 3350 167 3550 856
rect 3718 167 3826 856
rect 3994 167 4102 856
rect 4270 167 4378 856
rect 4546 167 4654 856
rect 4822 167 4930 856
rect 5098 167 5298 856
rect 5466 167 5574 856
rect 5742 167 5850 856
rect 6018 167 6126 856
rect 6294 167 6402 856
rect 6570 167 6770 856
rect 6938 167 7046 856
rect 7214 167 7322 856
rect 7490 167 7598 856
rect 7766 167 7874 856
rect 8042 167 8150 856
rect 8318 167 8518 856
rect 8686 167 8794 856
rect 8962 167 9070 856
rect 9238 167 9346 856
rect 9514 167 9622 856
rect 9790 167 9898 856
rect 10066 167 10266 856
rect 10434 167 10542 856
rect 10710 167 10818 856
rect 10986 167 11094 856
rect 11262 167 11370 856
rect 11538 167 11738 856
rect 11906 167 12014 856
rect 12182 167 12290 856
rect 12458 167 12566 856
rect 12734 167 12842 856
rect 13010 167 13118 856
rect 13286 167 13486 856
rect 13654 167 13762 856
rect 13930 167 14038 856
rect 14206 167 14314 856
rect 14482 167 14590 856
rect 14758 167 14866 856
rect 15034 167 15234 856
rect 15402 167 15510 856
rect 15678 167 15786 856
rect 15954 167 16062 856
rect 16230 167 16338 856
rect 16506 167 16614 856
rect 16782 167 16982 856
rect 17150 167 17258 856
rect 17426 167 17534 856
rect 17702 167 17810 856
rect 17978 167 18086 856
rect 18254 167 18454 856
rect 18622 167 18730 856
rect 18898 167 19006 856
rect 19174 167 19282 856
rect 19450 167 19558 856
rect 19726 167 19834 856
rect 20002 167 20202 856
rect 20370 167 20478 856
rect 20646 167 20754 856
rect 20922 167 21030 856
rect 21198 167 21306 856
rect 21474 167 21582 856
rect 21750 167 21950 856
rect 22118 167 22226 856
rect 22394 167 22502 856
rect 22670 167 22778 856
rect 22946 167 23054 856
rect 23222 167 23422 856
rect 23590 167 23698 856
rect 23866 167 23974 856
rect 24142 167 24250 856
rect 24418 167 24526 856
rect 24694 167 24802 856
rect 24970 167 25170 856
rect 25338 167 25446 856
rect 25614 167 25722 856
rect 25890 167 25998 856
rect 26166 167 26274 856
rect 26442 167 26550 856
rect 26718 167 26918 856
rect 27086 167 27194 856
rect 27362 167 27470 856
rect 27638 167 27746 856
rect 27914 167 28022 856
rect 28190 167 28298 856
rect 28466 167 28666 856
rect 28834 167 28942 856
rect 29110 167 29218 856
rect 29386 167 29494 856
rect 29662 167 29770 856
rect 29938 167 30138 856
rect 30306 167 30414 856
rect 30582 167 30690 856
rect 30858 167 30966 856
rect 31134 167 31242 856
rect 31410 167 31518 856
rect 31686 167 31886 856
rect 32054 167 32162 856
rect 32330 167 32438 856
rect 32606 167 32714 856
rect 32882 167 32990 856
rect 33158 167 33266 856
rect 33434 167 33634 856
rect 33802 167 33910 856
rect 34078 167 34186 856
rect 34354 167 34462 856
rect 34630 167 34738 856
rect 34906 167 35106 856
rect 35274 167 35382 856
rect 35550 167 35658 856
rect 35826 167 35934 856
rect 36102 167 36210 856
rect 36378 167 36486 856
rect 36654 167 36854 856
rect 37022 167 37130 856
rect 37298 167 37406 856
rect 37574 167 37682 856
rect 37850 167 37958 856
rect 38126 167 38234 856
rect 38402 167 38602 856
rect 38770 167 38878 856
rect 39046 167 39154 856
rect 39322 167 39430 856
rect 39598 167 39706 856
rect 39874 167 39908 856
<< metal3 >>
rect -800 119416 800 119536
rect 39200 119552 40800 119672
rect 39200 119144 40800 119264
rect -800 118600 800 118720
rect 39200 118736 40800 118856
rect 39200 118328 40800 118448
rect -800 117784 800 117904
rect 39200 117920 40800 118040
rect 39200 117376 40800 117496
rect -800 116968 800 117088
rect 39200 116968 40800 117088
rect 39200 116560 40800 116680
rect -800 116152 800 116272
rect 39200 116152 40800 116272
rect 39200 115744 40800 115864
rect -800 115336 800 115456
rect 39200 115336 40800 115456
rect 39200 114792 40800 114912
rect -800 114520 800 114640
rect 39200 114384 40800 114504
rect 39200 113976 40800 114096
rect -800 113704 800 113824
rect 39200 113568 40800 113688
rect 39200 113160 40800 113280
rect -800 112888 800 113008
rect 39200 112752 40800 112872
rect -800 112072 800 112192
rect 39200 112208 40800 112328
rect 39200 111800 40800 111920
rect -800 111256 800 111376
rect 39200 111392 40800 111512
rect 39200 110984 40800 111104
rect -800 110440 800 110560
rect 39200 110576 40800 110696
rect 39200 110168 40800 110288
rect -800 109488 800 109608
rect 39200 109624 40800 109744
rect 39200 109216 40800 109336
rect -800 108672 800 108792
rect 39200 108808 40800 108928
rect 39200 108400 40800 108520
rect -800 107856 800 107976
rect 39200 107992 40800 108112
rect 39200 107448 40800 107568
rect -800 107040 800 107160
rect 39200 107040 40800 107160
rect 39200 106632 40800 106752
rect -800 106224 800 106344
rect 39200 106224 40800 106344
rect 39200 105816 40800 105936
rect -800 105408 800 105528
rect 39200 105408 40800 105528
rect 39200 104864 40800 104984
rect -800 104592 800 104712
rect 39200 104456 40800 104576
rect 39200 104048 40800 104168
rect -800 103776 800 103896
rect 39200 103640 40800 103760
rect 39200 103232 40800 103352
rect -800 102960 800 103080
rect 39200 102824 40800 102944
rect -800 102144 800 102264
rect 39200 102280 40800 102400
rect 39200 101872 40800 101992
rect -800 101328 800 101448
rect 39200 101464 40800 101584
rect 39200 101056 40800 101176
rect -800 100512 800 100632
rect 39200 100648 40800 100768
rect 39200 100240 40800 100360
rect -800 99560 800 99680
rect 39200 99696 40800 99816
rect 39200 99288 40800 99408
rect -800 98744 800 98864
rect 39200 98880 40800 99000
rect 39200 98472 40800 98592
rect -800 97928 800 98048
rect 39200 98064 40800 98184
rect 39200 97656 40800 97776
rect -800 97112 800 97232
rect 39200 97112 40800 97232
rect 39200 96704 40800 96824
rect -800 96296 800 96416
rect 39200 96296 40800 96416
rect 39200 95888 40800 96008
rect -800 95480 800 95600
rect 39200 95480 40800 95600
rect 39200 94936 40800 95056
rect -800 94664 800 94784
rect 39200 94528 40800 94648
rect 39200 94120 40800 94240
rect -800 93848 800 93968
rect 39200 93712 40800 93832
rect 39200 93304 40800 93424
rect -800 93032 800 93152
rect 39200 92896 40800 93016
rect -800 92216 800 92336
rect 39200 92352 40800 92472
rect 39200 91944 40800 92064
rect -800 91400 800 91520
rect 39200 91536 40800 91656
rect 39200 91128 40800 91248
rect -800 90584 800 90704
rect 39200 90720 40800 90840
rect 39200 90312 40800 90432
rect -800 89632 800 89752
rect 39200 89768 40800 89888
rect 39200 89360 40800 89480
rect -800 88816 800 88936
rect 39200 88952 40800 89072
rect 39200 88544 40800 88664
rect -800 88000 800 88120
rect 39200 88136 40800 88256
rect 39200 87728 40800 87848
rect -800 87184 800 87304
rect 39200 87184 40800 87304
rect 39200 86776 40800 86896
rect -800 86368 800 86488
rect 39200 86368 40800 86488
rect 39200 85960 40800 86080
rect -800 85552 800 85672
rect 39200 85552 40800 85672
rect 39200 85144 40800 85264
rect -800 84736 800 84856
rect 39200 84600 40800 84720
rect 39200 84192 40800 84312
rect -800 83920 800 84040
rect 39200 83784 40800 83904
rect 39200 83376 40800 83496
rect -800 83104 800 83224
rect 39200 82968 40800 83088
rect -800 82288 800 82408
rect 39200 82424 40800 82544
rect 39200 82016 40800 82136
rect -800 81472 800 81592
rect 39200 81608 40800 81728
rect 39200 81200 40800 81320
rect -800 80656 800 80776
rect 39200 80792 40800 80912
rect 39200 80384 40800 80504
rect -800 79704 800 79824
rect 39200 79840 40800 79960
rect 39200 79432 40800 79552
rect -800 78888 800 79008
rect 39200 79024 40800 79144
rect 39200 78616 40800 78736
rect -800 78072 800 78192
rect 39200 78208 40800 78328
rect 39200 77800 40800 77920
rect -800 77256 800 77376
rect 39200 77256 40800 77376
rect 39200 76848 40800 76968
rect -800 76440 800 76560
rect 39200 76440 40800 76560
rect 39200 76032 40800 76152
rect -800 75624 800 75744
rect 39200 75624 40800 75744
rect 39200 75216 40800 75336
rect -800 74808 800 74928
rect 39200 74672 40800 74792
rect 39200 74264 40800 74384
rect -800 73992 800 74112
rect 39200 73856 40800 73976
rect 39200 73448 40800 73568
rect -800 73176 800 73296
rect 39200 73040 40800 73160
rect 39200 72632 40800 72752
rect -800 72360 800 72480
rect 39200 72088 40800 72208
rect -800 71544 800 71664
rect 39200 71680 40800 71800
rect 39200 71272 40800 71392
rect -800 70728 800 70848
rect 39200 70864 40800 70984
rect 39200 70456 40800 70576
rect -800 69776 800 69896
rect 39200 69912 40800 70032
rect 39200 69504 40800 69624
rect -800 68960 800 69080
rect 39200 69096 40800 69216
rect 39200 68688 40800 68808
rect -800 68144 800 68264
rect 39200 68280 40800 68400
rect 39200 67872 40800 67992
rect -800 67328 800 67448
rect 39200 67328 40800 67448
rect 39200 66920 40800 67040
rect -800 66512 800 66632
rect 39200 66512 40800 66632
rect 39200 66104 40800 66224
rect -800 65696 800 65816
rect 39200 65696 40800 65816
rect 39200 65288 40800 65408
rect -800 64880 800 65000
rect 39200 64744 40800 64864
rect 39200 64336 40800 64456
rect -800 64064 800 64184
rect 39200 63928 40800 64048
rect 39200 63520 40800 63640
rect -800 63248 800 63368
rect 39200 63112 40800 63232
rect 39200 62704 40800 62824
rect -800 62432 800 62552
rect 39200 62160 40800 62280
rect -800 61616 800 61736
rect 39200 61752 40800 61872
rect 39200 61344 40800 61464
rect -800 60800 800 60920
rect 39200 60936 40800 61056
rect 39200 60528 40800 60648
rect 39200 60120 40800 60240
rect -800 59848 800 59968
rect 39200 59576 40800 59696
rect -800 59032 800 59152
rect 39200 59168 40800 59288
rect 39200 58760 40800 58880
rect -800 58216 800 58336
rect 39200 58352 40800 58472
rect 39200 57944 40800 58064
rect -800 57400 800 57520
rect 39200 57400 40800 57520
rect 39200 56992 40800 57112
rect -800 56584 800 56704
rect 39200 56584 40800 56704
rect 39200 56176 40800 56296
rect -800 55768 800 55888
rect 39200 55768 40800 55888
rect 39200 55360 40800 55480
rect -800 54952 800 55072
rect 39200 54816 40800 54936
rect 39200 54408 40800 54528
rect -800 54136 800 54256
rect 39200 54000 40800 54120
rect 39200 53592 40800 53712
rect -800 53320 800 53440
rect 39200 53184 40800 53304
rect 39200 52776 40800 52896
rect -800 52504 800 52624
rect 39200 52232 40800 52352
rect -800 51688 800 51808
rect 39200 51824 40800 51944
rect 39200 51416 40800 51536
rect -800 50872 800 50992
rect 39200 51008 40800 51128
rect 39200 50600 40800 50720
rect 39200 50192 40800 50312
rect -800 49920 800 50040
rect 39200 49648 40800 49768
rect -800 49104 800 49224
rect 39200 49240 40800 49360
rect 39200 48832 40800 48952
rect -800 48288 800 48408
rect 39200 48424 40800 48544
rect 39200 48016 40800 48136
rect -800 47472 800 47592
rect 39200 47472 40800 47592
rect 39200 47064 40800 47184
rect -800 46656 800 46776
rect 39200 46656 40800 46776
rect 39200 46248 40800 46368
rect -800 45840 800 45960
rect 39200 45840 40800 45960
rect 39200 45432 40800 45552
rect -800 45024 800 45144
rect 39200 44888 40800 45008
rect 39200 44480 40800 44600
rect -800 44208 800 44328
rect 39200 44072 40800 44192
rect 39200 43664 40800 43784
rect -800 43392 800 43512
rect 39200 43256 40800 43376
rect 39200 42848 40800 42968
rect -800 42576 800 42696
rect 39200 42304 40800 42424
rect -800 41760 800 41880
rect 39200 41896 40800 42016
rect 39200 41488 40800 41608
rect -800 40944 800 41064
rect 39200 41080 40800 41200
rect 39200 40672 40800 40792
rect 39200 40264 40800 40384
rect -800 39992 800 40112
rect 39200 39720 40800 39840
rect -800 39176 800 39296
rect 39200 39312 40800 39432
rect 39200 38904 40800 39024
rect -800 38360 800 38480
rect 39200 38496 40800 38616
rect 39200 38088 40800 38208
rect -800 37544 800 37664
rect 39200 37680 40800 37800
rect 39200 37136 40800 37256
rect -800 36728 800 36848
rect 39200 36728 40800 36848
rect 39200 36320 40800 36440
rect -800 35912 800 36032
rect 39200 35912 40800 36032
rect 39200 35504 40800 35624
rect -800 35096 800 35216
rect 39200 34960 40800 35080
rect 39200 34552 40800 34672
rect -800 34280 800 34400
rect 39200 34144 40800 34264
rect 39200 33736 40800 33856
rect -800 33464 800 33584
rect 39200 33328 40800 33448
rect 39200 32920 40800 33040
rect -800 32648 800 32768
rect 39200 32376 40800 32496
rect -800 31832 800 31952
rect 39200 31968 40800 32088
rect 39200 31560 40800 31680
rect -800 31016 800 31136
rect 39200 31152 40800 31272
rect 39200 30744 40800 30864
rect 39200 30336 40800 30456
rect -800 30064 800 30184
rect 39200 29792 40800 29912
rect -800 29248 800 29368
rect 39200 29384 40800 29504
rect 39200 28976 40800 29096
rect -800 28432 800 28552
rect 39200 28568 40800 28688
rect 39200 28160 40800 28280
rect -800 27616 800 27736
rect 39200 27752 40800 27872
rect 39200 27208 40800 27328
rect -800 26800 800 26920
rect 39200 26800 40800 26920
rect 39200 26392 40800 26512
rect -800 25984 800 26104
rect 39200 25984 40800 26104
rect 39200 25576 40800 25696
rect -800 25168 800 25288
rect 39200 25168 40800 25288
rect 39200 24624 40800 24744
rect -800 24352 800 24472
rect 39200 24216 40800 24336
rect 39200 23808 40800 23928
rect -800 23536 800 23656
rect 39200 23400 40800 23520
rect 39200 22992 40800 23112
rect -800 22720 800 22840
rect 39200 22448 40800 22568
rect -800 21904 800 22024
rect 39200 22040 40800 22160
rect 39200 21632 40800 21752
rect -800 21088 800 21208
rect 39200 21224 40800 21344
rect 39200 20816 40800 20936
rect 39200 20408 40800 20528
rect -800 20136 800 20256
rect 39200 19864 40800 19984
rect -800 19320 800 19440
rect 39200 19456 40800 19576
rect 39200 19048 40800 19168
rect -800 18504 800 18624
rect 39200 18640 40800 18760
rect 39200 18232 40800 18352
rect -800 17688 800 17808
rect 39200 17824 40800 17944
rect 39200 17280 40800 17400
rect -800 16872 800 16992
rect 39200 16872 40800 16992
rect 39200 16464 40800 16584
rect -800 16056 800 16176
rect 39200 16056 40800 16176
rect 39200 15648 40800 15768
rect -800 15240 800 15360
rect 39200 15240 40800 15360
rect 39200 14696 40800 14816
rect -800 14424 800 14544
rect 39200 14288 40800 14408
rect 39200 13880 40800 14000
rect -800 13608 800 13728
rect 39200 13472 40800 13592
rect 39200 13064 40800 13184
rect -800 12792 800 12912
rect 39200 12656 40800 12776
rect -800 11976 800 12096
rect 39200 12112 40800 12232
rect 39200 11704 40800 11824
rect -800 11160 800 11280
rect 39200 11296 40800 11416
rect 39200 10888 40800 11008
rect 39200 10480 40800 10600
rect -800 10208 800 10328
rect 39200 9936 40800 10056
rect -800 9392 800 9512
rect 39200 9528 40800 9648
rect 39200 9120 40800 9240
rect -800 8576 800 8696
rect 39200 8712 40800 8832
rect 39200 8304 40800 8424
rect -800 7760 800 7880
rect 39200 7896 40800 8016
rect 39200 7352 40800 7472
rect -800 6944 800 7064
rect 39200 6944 40800 7064
rect 39200 6536 40800 6656
rect -800 6128 800 6248
rect 39200 6128 40800 6248
rect 39200 5720 40800 5840
rect -800 5312 800 5432
rect 39200 5312 40800 5432
rect 39200 4768 40800 4888
rect -800 4496 800 4616
rect 39200 4360 40800 4480
rect 39200 3952 40800 4072
rect -800 3680 800 3800
rect 39200 3544 40800 3664
rect 39200 3136 40800 3256
rect -800 2864 800 2984
rect 39200 2728 40800 2848
rect -800 2048 800 2168
rect 39200 2184 40800 2304
rect 39200 1776 40800 1896
rect -800 1232 800 1352
rect 39200 1368 40800 1488
rect 39200 960 40800 1080
rect -800 416 800 536
rect 39200 552 40800 672
rect 39200 144 40800 264
<< obsm3 >>
rect 800 119616 39120 119645
rect 880 119472 39120 119616
rect 880 119344 39200 119472
rect 880 119336 39120 119344
rect 800 119064 39120 119336
rect 800 118936 39200 119064
rect 800 118800 39120 118936
rect 880 118656 39120 118800
rect 880 118528 39200 118656
rect 880 118520 39120 118528
rect 800 118248 39120 118520
rect 800 118120 39200 118248
rect 800 117984 39120 118120
rect 880 117840 39120 117984
rect 880 117704 39200 117840
rect 800 117576 39200 117704
rect 800 117296 39120 117576
rect 800 117168 39200 117296
rect 880 116888 39120 117168
rect 800 116760 39200 116888
rect 800 116480 39120 116760
rect 800 116352 39200 116480
rect 880 116072 39120 116352
rect 800 115944 39200 116072
rect 800 115664 39120 115944
rect 800 115536 39200 115664
rect 880 115256 39120 115536
rect 800 114992 39200 115256
rect 800 114720 39120 114992
rect 880 114712 39120 114720
rect 880 114584 39200 114712
rect 880 114440 39120 114584
rect 800 114304 39120 114440
rect 800 114176 39200 114304
rect 800 113904 39120 114176
rect 880 113896 39120 113904
rect 880 113768 39200 113896
rect 880 113624 39120 113768
rect 800 113488 39120 113624
rect 800 113360 39200 113488
rect 800 113088 39120 113360
rect 880 113080 39120 113088
rect 880 112952 39200 113080
rect 880 112808 39120 112952
rect 800 112672 39120 112808
rect 800 112408 39200 112672
rect 800 112272 39120 112408
rect 880 112128 39120 112272
rect 880 112000 39200 112128
rect 880 111992 39120 112000
rect 800 111720 39120 111992
rect 800 111592 39200 111720
rect 800 111456 39120 111592
rect 880 111312 39120 111456
rect 880 111184 39200 111312
rect 880 111176 39120 111184
rect 800 110904 39120 111176
rect 800 110776 39200 110904
rect 800 110640 39120 110776
rect 880 110496 39120 110640
rect 880 110368 39200 110496
rect 880 110360 39120 110368
rect 800 110088 39120 110360
rect 800 109824 39200 110088
rect 800 109688 39120 109824
rect 880 109544 39120 109688
rect 880 109416 39200 109544
rect 880 109408 39120 109416
rect 800 109136 39120 109408
rect 800 109008 39200 109136
rect 800 108872 39120 109008
rect 880 108728 39120 108872
rect 880 108600 39200 108728
rect 880 108592 39120 108600
rect 800 108320 39120 108592
rect 800 108192 39200 108320
rect 800 108056 39120 108192
rect 880 107912 39120 108056
rect 880 107776 39200 107912
rect 800 107648 39200 107776
rect 800 107368 39120 107648
rect 800 107240 39200 107368
rect 880 106960 39120 107240
rect 800 106832 39200 106960
rect 800 106552 39120 106832
rect 800 106424 39200 106552
rect 880 106144 39120 106424
rect 800 106016 39200 106144
rect 800 105736 39120 106016
rect 800 105608 39200 105736
rect 880 105328 39120 105608
rect 800 105064 39200 105328
rect 800 104792 39120 105064
rect 880 104784 39120 104792
rect 880 104656 39200 104784
rect 880 104512 39120 104656
rect 800 104376 39120 104512
rect 800 104248 39200 104376
rect 800 103976 39120 104248
rect 880 103968 39120 103976
rect 880 103840 39200 103968
rect 880 103696 39120 103840
rect 800 103560 39120 103696
rect 800 103432 39200 103560
rect 800 103160 39120 103432
rect 880 103152 39120 103160
rect 880 103024 39200 103152
rect 880 102880 39120 103024
rect 800 102744 39120 102880
rect 800 102480 39200 102744
rect 800 102344 39120 102480
rect 880 102200 39120 102344
rect 880 102072 39200 102200
rect 880 102064 39120 102072
rect 800 101792 39120 102064
rect 800 101664 39200 101792
rect 800 101528 39120 101664
rect 880 101384 39120 101528
rect 880 101256 39200 101384
rect 880 101248 39120 101256
rect 800 100976 39120 101248
rect 800 100848 39200 100976
rect 800 100712 39120 100848
rect 880 100568 39120 100712
rect 880 100440 39200 100568
rect 880 100432 39120 100440
rect 800 100160 39120 100432
rect 800 99896 39200 100160
rect 800 99760 39120 99896
rect 880 99616 39120 99760
rect 880 99488 39200 99616
rect 880 99480 39120 99488
rect 800 99208 39120 99480
rect 800 99080 39200 99208
rect 800 98944 39120 99080
rect 880 98800 39120 98944
rect 880 98672 39200 98800
rect 880 98664 39120 98672
rect 800 98392 39120 98664
rect 800 98264 39200 98392
rect 800 98128 39120 98264
rect 880 97984 39120 98128
rect 880 97856 39200 97984
rect 880 97848 39120 97856
rect 800 97576 39120 97848
rect 800 97312 39200 97576
rect 880 97032 39120 97312
rect 800 96904 39200 97032
rect 800 96624 39120 96904
rect 800 96496 39200 96624
rect 880 96216 39120 96496
rect 800 96088 39200 96216
rect 800 95808 39120 96088
rect 800 95680 39200 95808
rect 880 95400 39120 95680
rect 800 95136 39200 95400
rect 800 94864 39120 95136
rect 880 94856 39120 94864
rect 880 94728 39200 94856
rect 880 94584 39120 94728
rect 800 94448 39120 94584
rect 800 94320 39200 94448
rect 800 94048 39120 94320
rect 880 94040 39120 94048
rect 880 93912 39200 94040
rect 880 93768 39120 93912
rect 800 93632 39120 93768
rect 800 93504 39200 93632
rect 800 93232 39120 93504
rect 880 93224 39120 93232
rect 880 93096 39200 93224
rect 880 92952 39120 93096
rect 800 92816 39120 92952
rect 800 92552 39200 92816
rect 800 92416 39120 92552
rect 880 92272 39120 92416
rect 880 92144 39200 92272
rect 880 92136 39120 92144
rect 800 91864 39120 92136
rect 800 91736 39200 91864
rect 800 91600 39120 91736
rect 880 91456 39120 91600
rect 880 91328 39200 91456
rect 880 91320 39120 91328
rect 800 91048 39120 91320
rect 800 90920 39200 91048
rect 800 90784 39120 90920
rect 880 90640 39120 90784
rect 880 90512 39200 90640
rect 880 90504 39120 90512
rect 800 90232 39120 90504
rect 800 89968 39200 90232
rect 800 89832 39120 89968
rect 880 89688 39120 89832
rect 880 89560 39200 89688
rect 880 89552 39120 89560
rect 800 89280 39120 89552
rect 800 89152 39200 89280
rect 800 89016 39120 89152
rect 880 88872 39120 89016
rect 880 88744 39200 88872
rect 880 88736 39120 88744
rect 800 88464 39120 88736
rect 800 88336 39200 88464
rect 800 88200 39120 88336
rect 880 88056 39120 88200
rect 880 87928 39200 88056
rect 880 87920 39120 87928
rect 800 87648 39120 87920
rect 800 87384 39200 87648
rect 880 87104 39120 87384
rect 800 86976 39200 87104
rect 800 86696 39120 86976
rect 800 86568 39200 86696
rect 880 86288 39120 86568
rect 800 86160 39200 86288
rect 800 85880 39120 86160
rect 800 85752 39200 85880
rect 880 85472 39120 85752
rect 800 85344 39200 85472
rect 800 85064 39120 85344
rect 800 84936 39200 85064
rect 880 84800 39200 84936
rect 880 84656 39120 84800
rect 800 84520 39120 84656
rect 800 84392 39200 84520
rect 800 84120 39120 84392
rect 880 84112 39120 84120
rect 880 83984 39200 84112
rect 880 83840 39120 83984
rect 800 83704 39120 83840
rect 800 83576 39200 83704
rect 800 83304 39120 83576
rect 880 83296 39120 83304
rect 880 83168 39200 83296
rect 880 83024 39120 83168
rect 800 82888 39120 83024
rect 800 82624 39200 82888
rect 800 82488 39120 82624
rect 880 82344 39120 82488
rect 880 82216 39200 82344
rect 880 82208 39120 82216
rect 800 81936 39120 82208
rect 800 81808 39200 81936
rect 800 81672 39120 81808
rect 880 81528 39120 81672
rect 880 81400 39200 81528
rect 880 81392 39120 81400
rect 800 81120 39120 81392
rect 800 80992 39200 81120
rect 800 80856 39120 80992
rect 880 80712 39120 80856
rect 880 80584 39200 80712
rect 880 80576 39120 80584
rect 800 80304 39120 80576
rect 800 80040 39200 80304
rect 800 79904 39120 80040
rect 880 79760 39120 79904
rect 880 79632 39200 79760
rect 880 79624 39120 79632
rect 800 79352 39120 79624
rect 800 79224 39200 79352
rect 800 79088 39120 79224
rect 880 78944 39120 79088
rect 880 78816 39200 78944
rect 880 78808 39120 78816
rect 800 78536 39120 78808
rect 800 78408 39200 78536
rect 800 78272 39120 78408
rect 880 78128 39120 78272
rect 880 78000 39200 78128
rect 880 77992 39120 78000
rect 800 77720 39120 77992
rect 800 77456 39200 77720
rect 880 77176 39120 77456
rect 800 77048 39200 77176
rect 800 76768 39120 77048
rect 800 76640 39200 76768
rect 880 76360 39120 76640
rect 800 76232 39200 76360
rect 800 75952 39120 76232
rect 800 75824 39200 75952
rect 880 75544 39120 75824
rect 800 75416 39200 75544
rect 800 75136 39120 75416
rect 800 75008 39200 75136
rect 880 74872 39200 75008
rect 880 74728 39120 74872
rect 800 74592 39120 74728
rect 800 74464 39200 74592
rect 800 74192 39120 74464
rect 880 74184 39120 74192
rect 880 74056 39200 74184
rect 880 73912 39120 74056
rect 800 73776 39120 73912
rect 800 73648 39200 73776
rect 800 73376 39120 73648
rect 880 73368 39120 73376
rect 880 73240 39200 73368
rect 880 73096 39120 73240
rect 800 72960 39120 73096
rect 800 72832 39200 72960
rect 800 72560 39120 72832
rect 880 72552 39120 72560
rect 880 72288 39200 72552
rect 880 72280 39120 72288
rect 800 72008 39120 72280
rect 800 71880 39200 72008
rect 800 71744 39120 71880
rect 880 71600 39120 71744
rect 880 71472 39200 71600
rect 880 71464 39120 71472
rect 800 71192 39120 71464
rect 800 71064 39200 71192
rect 800 70928 39120 71064
rect 880 70784 39120 70928
rect 880 70656 39200 70784
rect 880 70648 39120 70656
rect 800 70376 39120 70648
rect 800 70112 39200 70376
rect 800 69976 39120 70112
rect 880 69832 39120 69976
rect 880 69704 39200 69832
rect 880 69696 39120 69704
rect 800 69424 39120 69696
rect 800 69296 39200 69424
rect 800 69160 39120 69296
rect 880 69016 39120 69160
rect 880 68888 39200 69016
rect 880 68880 39120 68888
rect 800 68608 39120 68880
rect 800 68480 39200 68608
rect 800 68344 39120 68480
rect 880 68200 39120 68344
rect 880 68072 39200 68200
rect 880 68064 39120 68072
rect 800 67792 39120 68064
rect 800 67528 39200 67792
rect 880 67248 39120 67528
rect 800 67120 39200 67248
rect 800 66840 39120 67120
rect 800 66712 39200 66840
rect 880 66432 39120 66712
rect 800 66304 39200 66432
rect 800 66024 39120 66304
rect 800 65896 39200 66024
rect 880 65616 39120 65896
rect 800 65488 39200 65616
rect 800 65208 39120 65488
rect 800 65080 39200 65208
rect 880 64944 39200 65080
rect 880 64800 39120 64944
rect 800 64664 39120 64800
rect 800 64536 39200 64664
rect 800 64264 39120 64536
rect 880 64256 39120 64264
rect 880 64128 39200 64256
rect 880 63984 39120 64128
rect 800 63848 39120 63984
rect 800 63720 39200 63848
rect 800 63448 39120 63720
rect 880 63440 39120 63448
rect 880 63312 39200 63440
rect 880 63168 39120 63312
rect 800 63032 39120 63168
rect 800 62904 39200 63032
rect 800 62632 39120 62904
rect 880 62624 39120 62632
rect 880 62360 39200 62624
rect 880 62352 39120 62360
rect 800 62080 39120 62352
rect 800 61952 39200 62080
rect 800 61816 39120 61952
rect 880 61672 39120 61816
rect 880 61544 39200 61672
rect 880 61536 39120 61544
rect 800 61264 39120 61536
rect 800 61136 39200 61264
rect 800 61000 39120 61136
rect 880 60856 39120 61000
rect 880 60728 39200 60856
rect 880 60720 39120 60728
rect 800 60448 39120 60720
rect 800 60320 39200 60448
rect 800 60048 39120 60320
rect 880 60040 39120 60048
rect 880 59776 39200 60040
rect 880 59768 39120 59776
rect 800 59496 39120 59768
rect 800 59368 39200 59496
rect 800 59232 39120 59368
rect 880 59088 39120 59232
rect 880 58960 39200 59088
rect 880 58952 39120 58960
rect 800 58680 39120 58952
rect 800 58552 39200 58680
rect 800 58416 39120 58552
rect 880 58272 39120 58416
rect 880 58144 39200 58272
rect 880 58136 39120 58144
rect 800 57864 39120 58136
rect 800 57600 39200 57864
rect 880 57320 39120 57600
rect 800 57192 39200 57320
rect 800 56912 39120 57192
rect 800 56784 39200 56912
rect 880 56504 39120 56784
rect 800 56376 39200 56504
rect 800 56096 39120 56376
rect 800 55968 39200 56096
rect 880 55688 39120 55968
rect 800 55560 39200 55688
rect 800 55280 39120 55560
rect 800 55152 39200 55280
rect 880 55016 39200 55152
rect 880 54872 39120 55016
rect 800 54736 39120 54872
rect 800 54608 39200 54736
rect 800 54336 39120 54608
rect 880 54328 39120 54336
rect 880 54200 39200 54328
rect 880 54056 39120 54200
rect 800 53920 39120 54056
rect 800 53792 39200 53920
rect 800 53520 39120 53792
rect 880 53512 39120 53520
rect 880 53384 39200 53512
rect 880 53240 39120 53384
rect 800 53104 39120 53240
rect 800 52976 39200 53104
rect 800 52704 39120 52976
rect 880 52696 39120 52704
rect 880 52432 39200 52696
rect 880 52424 39120 52432
rect 800 52152 39120 52424
rect 800 52024 39200 52152
rect 800 51888 39120 52024
rect 880 51744 39120 51888
rect 880 51616 39200 51744
rect 880 51608 39120 51616
rect 800 51336 39120 51608
rect 800 51208 39200 51336
rect 800 51072 39120 51208
rect 880 50928 39120 51072
rect 880 50800 39200 50928
rect 880 50792 39120 50800
rect 800 50520 39120 50792
rect 800 50392 39200 50520
rect 800 50120 39120 50392
rect 880 50112 39120 50120
rect 880 49848 39200 50112
rect 880 49840 39120 49848
rect 800 49568 39120 49840
rect 800 49440 39200 49568
rect 800 49304 39120 49440
rect 880 49160 39120 49304
rect 880 49032 39200 49160
rect 880 49024 39120 49032
rect 800 48752 39120 49024
rect 800 48624 39200 48752
rect 800 48488 39120 48624
rect 880 48344 39120 48488
rect 880 48216 39200 48344
rect 880 48208 39120 48216
rect 800 47936 39120 48208
rect 800 47672 39200 47936
rect 880 47392 39120 47672
rect 800 47264 39200 47392
rect 800 46984 39120 47264
rect 800 46856 39200 46984
rect 880 46576 39120 46856
rect 800 46448 39200 46576
rect 800 46168 39120 46448
rect 800 46040 39200 46168
rect 880 45760 39120 46040
rect 800 45632 39200 45760
rect 800 45352 39120 45632
rect 800 45224 39200 45352
rect 880 45088 39200 45224
rect 880 44944 39120 45088
rect 800 44808 39120 44944
rect 800 44680 39200 44808
rect 800 44408 39120 44680
rect 880 44400 39120 44408
rect 880 44272 39200 44400
rect 880 44128 39120 44272
rect 800 43992 39120 44128
rect 800 43864 39200 43992
rect 800 43592 39120 43864
rect 880 43584 39120 43592
rect 880 43456 39200 43584
rect 880 43312 39120 43456
rect 800 43176 39120 43312
rect 800 43048 39200 43176
rect 800 42776 39120 43048
rect 880 42768 39120 42776
rect 880 42504 39200 42768
rect 880 42496 39120 42504
rect 800 42224 39120 42496
rect 800 42096 39200 42224
rect 800 41960 39120 42096
rect 880 41816 39120 41960
rect 880 41688 39200 41816
rect 880 41680 39120 41688
rect 800 41408 39120 41680
rect 800 41280 39200 41408
rect 800 41144 39120 41280
rect 880 41000 39120 41144
rect 880 40872 39200 41000
rect 880 40864 39120 40872
rect 800 40592 39120 40864
rect 800 40464 39200 40592
rect 800 40192 39120 40464
rect 880 40184 39120 40192
rect 880 39920 39200 40184
rect 880 39912 39120 39920
rect 800 39640 39120 39912
rect 800 39512 39200 39640
rect 800 39376 39120 39512
rect 880 39232 39120 39376
rect 880 39104 39200 39232
rect 880 39096 39120 39104
rect 800 38824 39120 39096
rect 800 38696 39200 38824
rect 800 38560 39120 38696
rect 880 38416 39120 38560
rect 880 38288 39200 38416
rect 880 38280 39120 38288
rect 800 38008 39120 38280
rect 800 37880 39200 38008
rect 800 37744 39120 37880
rect 880 37600 39120 37744
rect 880 37464 39200 37600
rect 800 37336 39200 37464
rect 800 37056 39120 37336
rect 800 36928 39200 37056
rect 880 36648 39120 36928
rect 800 36520 39200 36648
rect 800 36240 39120 36520
rect 800 36112 39200 36240
rect 880 35832 39120 36112
rect 800 35704 39200 35832
rect 800 35424 39120 35704
rect 800 35296 39200 35424
rect 880 35160 39200 35296
rect 880 35016 39120 35160
rect 800 34880 39120 35016
rect 800 34752 39200 34880
rect 800 34480 39120 34752
rect 880 34472 39120 34480
rect 880 34344 39200 34472
rect 880 34200 39120 34344
rect 800 34064 39120 34200
rect 800 33936 39200 34064
rect 800 33664 39120 33936
rect 880 33656 39120 33664
rect 880 33528 39200 33656
rect 880 33384 39120 33528
rect 800 33248 39120 33384
rect 800 33120 39200 33248
rect 800 32848 39120 33120
rect 880 32840 39120 32848
rect 880 32576 39200 32840
rect 880 32568 39120 32576
rect 800 32296 39120 32568
rect 800 32168 39200 32296
rect 800 32032 39120 32168
rect 880 31888 39120 32032
rect 880 31760 39200 31888
rect 880 31752 39120 31760
rect 800 31480 39120 31752
rect 800 31352 39200 31480
rect 800 31216 39120 31352
rect 880 31072 39120 31216
rect 880 30944 39200 31072
rect 880 30936 39120 30944
rect 800 30664 39120 30936
rect 800 30536 39200 30664
rect 800 30264 39120 30536
rect 880 30256 39120 30264
rect 880 29992 39200 30256
rect 880 29984 39120 29992
rect 800 29712 39120 29984
rect 800 29584 39200 29712
rect 800 29448 39120 29584
rect 880 29304 39120 29448
rect 880 29176 39200 29304
rect 880 29168 39120 29176
rect 800 28896 39120 29168
rect 800 28768 39200 28896
rect 800 28632 39120 28768
rect 880 28488 39120 28632
rect 880 28360 39200 28488
rect 880 28352 39120 28360
rect 800 28080 39120 28352
rect 800 27952 39200 28080
rect 800 27816 39120 27952
rect 880 27672 39120 27816
rect 880 27536 39200 27672
rect 800 27408 39200 27536
rect 800 27128 39120 27408
rect 800 27000 39200 27128
rect 880 26720 39120 27000
rect 800 26592 39200 26720
rect 800 26312 39120 26592
rect 800 26184 39200 26312
rect 880 25904 39120 26184
rect 800 25776 39200 25904
rect 800 25496 39120 25776
rect 800 25368 39200 25496
rect 880 25088 39120 25368
rect 800 24824 39200 25088
rect 800 24552 39120 24824
rect 880 24544 39120 24552
rect 880 24416 39200 24544
rect 880 24272 39120 24416
rect 800 24136 39120 24272
rect 800 24008 39200 24136
rect 800 23736 39120 24008
rect 880 23728 39120 23736
rect 880 23600 39200 23728
rect 880 23456 39120 23600
rect 800 23320 39120 23456
rect 800 23192 39200 23320
rect 800 22920 39120 23192
rect 880 22912 39120 22920
rect 880 22648 39200 22912
rect 880 22640 39120 22648
rect 800 22368 39120 22640
rect 800 22240 39200 22368
rect 800 22104 39120 22240
rect 880 21960 39120 22104
rect 880 21832 39200 21960
rect 880 21824 39120 21832
rect 800 21552 39120 21824
rect 800 21424 39200 21552
rect 800 21288 39120 21424
rect 880 21144 39120 21288
rect 880 21016 39200 21144
rect 880 21008 39120 21016
rect 800 20736 39120 21008
rect 800 20608 39200 20736
rect 800 20336 39120 20608
rect 880 20328 39120 20336
rect 880 20064 39200 20328
rect 880 20056 39120 20064
rect 800 19784 39120 20056
rect 800 19656 39200 19784
rect 800 19520 39120 19656
rect 880 19376 39120 19520
rect 880 19248 39200 19376
rect 880 19240 39120 19248
rect 800 18968 39120 19240
rect 800 18840 39200 18968
rect 800 18704 39120 18840
rect 880 18560 39120 18704
rect 880 18432 39200 18560
rect 880 18424 39120 18432
rect 800 18152 39120 18424
rect 800 18024 39200 18152
rect 800 17888 39120 18024
rect 880 17744 39120 17888
rect 880 17608 39200 17744
rect 800 17480 39200 17608
rect 800 17200 39120 17480
rect 800 17072 39200 17200
rect 880 16792 39120 17072
rect 800 16664 39200 16792
rect 800 16384 39120 16664
rect 800 16256 39200 16384
rect 880 15976 39120 16256
rect 800 15848 39200 15976
rect 800 15568 39120 15848
rect 800 15440 39200 15568
rect 880 15160 39120 15440
rect 800 14896 39200 15160
rect 800 14624 39120 14896
rect 880 14616 39120 14624
rect 880 14488 39200 14616
rect 880 14344 39120 14488
rect 800 14208 39120 14344
rect 800 14080 39200 14208
rect 800 13808 39120 14080
rect 880 13800 39120 13808
rect 880 13672 39200 13800
rect 880 13528 39120 13672
rect 800 13392 39120 13528
rect 800 13264 39200 13392
rect 800 12992 39120 13264
rect 880 12984 39120 12992
rect 880 12856 39200 12984
rect 880 12712 39120 12856
rect 800 12576 39120 12712
rect 800 12312 39200 12576
rect 800 12176 39120 12312
rect 880 12032 39120 12176
rect 880 11904 39200 12032
rect 880 11896 39120 11904
rect 800 11624 39120 11896
rect 800 11496 39200 11624
rect 800 11360 39120 11496
rect 880 11216 39120 11360
rect 880 11088 39200 11216
rect 880 11080 39120 11088
rect 800 10808 39120 11080
rect 800 10680 39200 10808
rect 800 10408 39120 10680
rect 880 10400 39120 10408
rect 880 10136 39200 10400
rect 880 10128 39120 10136
rect 800 9856 39120 10128
rect 800 9728 39200 9856
rect 800 9592 39120 9728
rect 880 9448 39120 9592
rect 880 9320 39200 9448
rect 880 9312 39120 9320
rect 800 9040 39120 9312
rect 800 8912 39200 9040
rect 800 8776 39120 8912
rect 880 8632 39120 8776
rect 880 8504 39200 8632
rect 880 8496 39120 8504
rect 800 8224 39120 8496
rect 800 8096 39200 8224
rect 800 7960 39120 8096
rect 880 7816 39120 7960
rect 880 7680 39200 7816
rect 800 7552 39200 7680
rect 800 7272 39120 7552
rect 800 7144 39200 7272
rect 880 6864 39120 7144
rect 800 6736 39200 6864
rect 800 6456 39120 6736
rect 800 6328 39200 6456
rect 880 6048 39120 6328
rect 800 5920 39200 6048
rect 800 5640 39120 5920
rect 800 5512 39200 5640
rect 880 5232 39120 5512
rect 800 4968 39200 5232
rect 800 4696 39120 4968
rect 880 4688 39120 4696
rect 880 4560 39200 4688
rect 880 4416 39120 4560
rect 800 4280 39120 4416
rect 800 4152 39200 4280
rect 800 3880 39120 4152
rect 880 3872 39120 3880
rect 880 3744 39200 3872
rect 880 3600 39120 3744
rect 800 3464 39120 3600
rect 800 3336 39200 3464
rect 800 3064 39120 3336
rect 880 3056 39120 3064
rect 880 2928 39200 3056
rect 880 2784 39120 2928
rect 800 2648 39120 2784
rect 800 2384 39200 2648
rect 800 2248 39120 2384
rect 880 2104 39120 2248
rect 880 1976 39200 2104
rect 880 1968 39120 1976
rect 800 1696 39120 1968
rect 800 1568 39200 1696
rect 800 1432 39120 1568
rect 880 1288 39120 1432
rect 880 1160 39200 1288
rect 880 1152 39120 1160
rect 800 880 39120 1152
rect 800 752 39200 880
rect 800 616 39120 752
rect 880 472 39120 616
rect 880 344 39200 472
rect 880 336 39120 344
rect 800 171 39120 336
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
<< labels >>
rlabel metal2 s 110 119200 166 120800 6 dsi[0]
port 1 nsew signal output
rlabel metal2 s 294 119200 350 120800 6 dsi[1]
port 2 nsew signal output
rlabel metal2 s 478 119200 534 120800 6 dsi[2]
port 3 nsew signal output
rlabel metal2 s 662 119200 718 120800 6 dsi[3]
port 4 nsew signal output
rlabel metal2 s 938 119200 994 120800 6 dsi[4]
port 5 nsew signal output
rlabel metal2 s 1122 119200 1178 120800 6 dsi[5]
port 6 nsew signal output
rlabel metal2 s 1306 119200 1362 120800 6 dsi[6]
port 7 nsew signal output
rlabel metal2 s 1582 119200 1638 120800 6 dsi[7]
port 8 nsew signal output
rlabel metal2 s 1766 119200 1822 120800 6 io_in[0]
port 9 nsew signal input
rlabel metal2 s 8114 119200 8170 120800 6 io_in[10]
port 10 nsew signal input
rlabel metal2 s 8758 119200 8814 120800 6 io_in[11]
port 11 nsew signal input
rlabel metal2 s 9402 119200 9458 120800 6 io_in[12]
port 12 nsew signal input
rlabel metal2 s 10046 119200 10102 120800 6 io_in[13]
port 13 nsew signal input
rlabel metal2 s 10690 119200 10746 120800 6 io_in[14]
port 14 nsew signal input
rlabel metal2 s 11242 119200 11298 120800 6 io_in[15]
port 15 nsew signal input
rlabel metal2 s 11886 119200 11942 120800 6 io_in[16]
port 16 nsew signal input
rlabel metal2 s 12530 119200 12586 120800 6 io_in[17]
port 17 nsew signal input
rlabel metal2 s 13174 119200 13230 120800 6 io_in[18]
port 18 nsew signal input
rlabel metal2 s 13818 119200 13874 120800 6 io_in[19]
port 19 nsew signal input
rlabel metal2 s 2410 119200 2466 120800 6 io_in[1]
port 20 nsew signal input
rlabel metal2 s 14462 119200 14518 120800 6 io_in[20]
port 21 nsew signal input
rlabel metal2 s 15106 119200 15162 120800 6 io_in[21]
port 22 nsew signal input
rlabel metal2 s 15750 119200 15806 120800 6 io_in[22]
port 23 nsew signal input
rlabel metal2 s 16394 119200 16450 120800 6 io_in[23]
port 24 nsew signal input
rlabel metal2 s 17038 119200 17094 120800 6 io_in[24]
port 25 nsew signal input
rlabel metal2 s 17682 119200 17738 120800 6 io_in[25]
port 26 nsew signal input
rlabel metal2 s 18234 119200 18290 120800 6 io_in[26]
port 27 nsew signal input
rlabel metal2 s 18878 119200 18934 120800 6 io_in[27]
port 28 nsew signal input
rlabel metal2 s 19522 119200 19578 120800 6 io_in[28]
port 29 nsew signal input
rlabel metal2 s 20166 119200 20222 120800 6 io_in[29]
port 30 nsew signal input
rlabel metal2 s 3054 119200 3110 120800 6 io_in[2]
port 31 nsew signal input
rlabel metal2 s 20810 119200 20866 120800 6 io_in[30]
port 32 nsew signal input
rlabel metal2 s 21454 119200 21510 120800 6 io_in[31]
port 33 nsew signal input
rlabel metal2 s 22098 119200 22154 120800 6 io_in[32]
port 34 nsew signal input
rlabel metal2 s 22742 119200 22798 120800 6 io_in[33]
port 35 nsew signal input
rlabel metal2 s 23386 119200 23442 120800 6 io_in[34]
port 36 nsew signal input
rlabel metal2 s 24030 119200 24086 120800 6 io_in[35]
port 37 nsew signal input
rlabel metal2 s 24582 119200 24638 120800 6 io_in[36]
port 38 nsew signal input
rlabel metal2 s 25226 119200 25282 120800 6 io_in[37]
port 39 nsew signal input
rlabel metal2 s 3698 119200 3754 120800 6 io_in[3]
port 40 nsew signal input
rlabel metal2 s 4342 119200 4398 120800 6 io_in[4]
port 41 nsew signal input
rlabel metal2 s 4894 119200 4950 120800 6 io_in[5]
port 42 nsew signal input
rlabel metal2 s 5538 119200 5594 120800 6 io_in[6]
port 43 nsew signal input
rlabel metal2 s 6182 119200 6238 120800 6 io_in[7]
port 44 nsew signal input
rlabel metal2 s 6826 119200 6882 120800 6 io_in[8]
port 45 nsew signal input
rlabel metal2 s 7470 119200 7526 120800 6 io_in[9]
port 46 nsew signal input
rlabel metal2 s 1950 119200 2006 120800 6 io_oeb[0]
port 47 nsew signal output
rlabel metal2 s 8298 119200 8354 120800 6 io_oeb[10]
port 48 nsew signal output
rlabel metal2 s 8942 119200 8998 120800 6 io_oeb[11]
port 49 nsew signal output
rlabel metal2 s 9586 119200 9642 120800 6 io_oeb[12]
port 50 nsew signal output
rlabel metal2 s 10230 119200 10286 120800 6 io_oeb[13]
port 51 nsew signal output
rlabel metal2 s 10874 119200 10930 120800 6 io_oeb[14]
port 52 nsew signal output
rlabel metal2 s 11518 119200 11574 120800 6 io_oeb[15]
port 53 nsew signal output
rlabel metal2 s 12162 119200 12218 120800 6 io_oeb[16]
port 54 nsew signal output
rlabel metal2 s 12806 119200 12862 120800 6 io_oeb[17]
port 55 nsew signal output
rlabel metal2 s 13450 119200 13506 120800 6 io_oeb[18]
port 56 nsew signal output
rlabel metal2 s 14002 119200 14058 120800 6 io_oeb[19]
port 57 nsew signal output
rlabel metal2 s 2594 119200 2650 120800 6 io_oeb[1]
port 58 nsew signal output
rlabel metal2 s 14646 119200 14702 120800 6 io_oeb[20]
port 59 nsew signal output
rlabel metal2 s 15290 119200 15346 120800 6 io_oeb[21]
port 60 nsew signal output
rlabel metal2 s 15934 119200 15990 120800 6 io_oeb[22]
port 61 nsew signal output
rlabel metal2 s 16578 119200 16634 120800 6 io_oeb[23]
port 62 nsew signal output
rlabel metal2 s 17222 119200 17278 120800 6 io_oeb[24]
port 63 nsew signal output
rlabel metal2 s 17866 119200 17922 120800 6 io_oeb[25]
port 64 nsew signal output
rlabel metal2 s 18510 119200 18566 120800 6 io_oeb[26]
port 65 nsew signal output
rlabel metal2 s 19154 119200 19210 120800 6 io_oeb[27]
port 66 nsew signal output
rlabel metal2 s 19798 119200 19854 120800 6 io_oeb[28]
port 67 nsew signal output
rlabel metal2 s 20350 119200 20406 120800 6 io_oeb[29]
port 68 nsew signal output
rlabel metal2 s 3238 119200 3294 120800 6 io_oeb[2]
port 69 nsew signal output
rlabel metal2 s 20994 119200 21050 120800 6 io_oeb[30]
port 70 nsew signal output
rlabel metal2 s 21638 119200 21694 120800 6 io_oeb[31]
port 71 nsew signal output
rlabel metal2 s 22282 119200 22338 120800 6 io_oeb[32]
port 72 nsew signal output
rlabel metal2 s 22926 119200 22982 120800 6 io_oeb[33]
port 73 nsew signal output
rlabel metal2 s 23570 119200 23626 120800 6 io_oeb[34]
port 74 nsew signal output
rlabel metal2 s 24214 119200 24270 120800 6 io_oeb[35]
port 75 nsew signal output
rlabel metal2 s 24858 119200 24914 120800 6 io_oeb[36]
port 76 nsew signal output
rlabel metal2 s 25502 119200 25558 120800 6 io_oeb[37]
port 77 nsew signal output
rlabel metal2 s 3882 119200 3938 120800 6 io_oeb[3]
port 78 nsew signal output
rlabel metal2 s 4526 119200 4582 120800 6 io_oeb[4]
port 79 nsew signal output
rlabel metal2 s 5170 119200 5226 120800 6 io_oeb[5]
port 80 nsew signal output
rlabel metal2 s 5814 119200 5870 120800 6 io_oeb[6]
port 81 nsew signal output
rlabel metal2 s 6458 119200 6514 120800 6 io_oeb[7]
port 82 nsew signal output
rlabel metal2 s 7010 119200 7066 120800 6 io_oeb[8]
port 83 nsew signal output
rlabel metal2 s 7654 119200 7710 120800 6 io_oeb[9]
port 84 nsew signal output
rlabel metal2 s 2226 119200 2282 120800 6 io_out[0]
port 85 nsew signal output
rlabel metal2 s 8574 119200 8630 120800 6 io_out[10]
port 86 nsew signal output
rlabel metal2 s 9126 119200 9182 120800 6 io_out[11]
port 87 nsew signal output
rlabel metal2 s 9770 119200 9826 120800 6 io_out[12]
port 88 nsew signal output
rlabel metal2 s 10414 119200 10470 120800 6 io_out[13]
port 89 nsew signal output
rlabel metal2 s 11058 119200 11114 120800 6 io_out[14]
port 90 nsew signal output
rlabel metal2 s 11702 119200 11758 120800 6 io_out[15]
port 91 nsew signal output
rlabel metal2 s 12346 119200 12402 120800 6 io_out[16]
port 92 nsew signal output
rlabel metal2 s 12990 119200 13046 120800 6 io_out[17]
port 93 nsew signal output
rlabel metal2 s 13634 119200 13690 120800 6 io_out[18]
port 94 nsew signal output
rlabel metal2 s 14278 119200 14334 120800 6 io_out[19]
port 95 nsew signal output
rlabel metal2 s 2778 119200 2834 120800 6 io_out[1]
port 96 nsew signal output
rlabel metal2 s 14922 119200 14978 120800 6 io_out[20]
port 97 nsew signal output
rlabel metal2 s 15566 119200 15622 120800 6 io_out[21]
port 98 nsew signal output
rlabel metal2 s 16118 119200 16174 120800 6 io_out[22]
port 99 nsew signal output
rlabel metal2 s 16762 119200 16818 120800 6 io_out[23]
port 100 nsew signal output
rlabel metal2 s 17406 119200 17462 120800 6 io_out[24]
port 101 nsew signal output
rlabel metal2 s 18050 119200 18106 120800 6 io_out[25]
port 102 nsew signal output
rlabel metal2 s 18694 119200 18750 120800 6 io_out[26]
port 103 nsew signal output
rlabel metal2 s 19338 119200 19394 120800 6 io_out[27]
port 104 nsew signal output
rlabel metal2 s 19982 119200 20038 120800 6 io_out[28]
port 105 nsew signal output
rlabel metal2 s 20626 119200 20682 120800 6 io_out[29]
port 106 nsew signal output
rlabel metal2 s 3422 119200 3478 120800 6 io_out[2]
port 107 nsew signal output
rlabel metal2 s 21270 119200 21326 120800 6 io_out[30]
port 108 nsew signal output
rlabel metal2 s 21914 119200 21970 120800 6 io_out[31]
port 109 nsew signal output
rlabel metal2 s 22466 119200 22522 120800 6 io_out[32]
port 110 nsew signal output
rlabel metal2 s 23110 119200 23166 120800 6 io_out[33]
port 111 nsew signal output
rlabel metal2 s 23754 119200 23810 120800 6 io_out[34]
port 112 nsew signal output
rlabel metal2 s 24398 119200 24454 120800 6 io_out[35]
port 113 nsew signal output
rlabel metal2 s 25042 119200 25098 120800 6 io_out[36]
port 114 nsew signal output
rlabel metal2 s 25686 119200 25742 120800 6 io_out[37]
port 115 nsew signal output
rlabel metal2 s 4066 119200 4122 120800 6 io_out[3]
port 116 nsew signal output
rlabel metal2 s 4710 119200 4766 120800 6 io_out[4]
port 117 nsew signal output
rlabel metal2 s 5354 119200 5410 120800 6 io_out[5]
port 118 nsew signal output
rlabel metal2 s 5998 119200 6054 120800 6 io_out[6]
port 119 nsew signal output
rlabel metal2 s 6642 119200 6698 120800 6 io_out[7]
port 120 nsew signal output
rlabel metal2 s 7286 119200 7342 120800 6 io_out[8]
port 121 nsew signal output
rlabel metal2 s 7930 119200 7986 120800 6 io_out[9]
port 122 nsew signal output
rlabel metal2 s 662 -800 718 800 8 irq[0]
port 123 nsew signal output
rlabel metal2 s 938 -800 994 800 8 irq[1]
port 124 nsew signal output
rlabel metal2 s 1214 -800 1270 800 8 irq[2]
port 125 nsew signal output
rlabel metal2 s 31942 -800 31998 800 8 la_reset[0]
port 126 nsew signal input
rlabel metal2 s 34794 -800 34850 800 8 la_reset[10]
port 127 nsew signal input
rlabel metal2 s 35162 -800 35218 800 8 la_reset[11]
port 128 nsew signal input
rlabel metal2 s 32218 -800 32274 800 8 la_reset[1]
port 129 nsew signal input
rlabel metal2 s 32494 -800 32550 800 8 la_reset[2]
port 130 nsew signal input
rlabel metal2 s 32770 -800 32826 800 8 la_reset[3]
port 131 nsew signal input
rlabel metal2 s 33046 -800 33102 800 8 la_reset[4]
port 132 nsew signal input
rlabel metal2 s 33322 -800 33378 800 8 la_reset[5]
port 133 nsew signal input
rlabel metal2 s 33690 -800 33746 800 8 la_reset[6]
port 134 nsew signal input
rlabel metal2 s 33966 -800 34022 800 8 la_reset[7]
port 135 nsew signal input
rlabel metal2 s 34242 -800 34298 800 8 la_reset[8]
port 136 nsew signal input
rlabel metal2 s 34518 -800 34574 800 8 la_reset[9]
port 137 nsew signal input
rlabel metal2 s 31574 119200 31630 120800 6 m_irqs[0]
port 138 nsew signal input
rlabel metal2 s 33690 119200 33746 120800 6 m_irqs[10]
port 139 nsew signal input
rlabel metal2 s 33966 119200 34022 120800 6 m_irqs[11]
port 140 nsew signal input
rlabel metal2 s 31850 119200 31906 120800 6 m_irqs[1]
port 141 nsew signal input
rlabel metal2 s 32034 119200 32090 120800 6 m_irqs[2]
port 142 nsew signal input
rlabel metal2 s 32218 119200 32274 120800 6 m_irqs[3]
port 143 nsew signal input
rlabel metal2 s 32494 119200 32550 120800 6 m_irqs[4]
port 144 nsew signal input
rlabel metal2 s 32678 119200 32734 120800 6 m_irqs[5]
port 145 nsew signal input
rlabel metal2 s 32862 119200 32918 120800 6 m_irqs[6]
port 146 nsew signal input
rlabel metal2 s 33138 119200 33194 120800 6 m_irqs[7]
port 147 nsew signal input
rlabel metal2 s 33322 119200 33378 120800 6 m_irqs[8]
port 148 nsew signal input
rlabel metal2 s 33506 119200 33562 120800 6 m_irqs[9]
port 149 nsew signal input
rlabel metal2 s 34150 119200 34206 120800 6 m_la_reset[0]
port 150 nsew signal output
rlabel metal2 s 36266 119200 36322 120800 6 m_la_reset[10]
port 151 nsew signal output
rlabel metal2 s 36450 119200 36506 120800 6 m_la_reset[11]
port 152 nsew signal output
rlabel metal2 s 34334 119200 34390 120800 6 m_la_reset[1]
port 153 nsew signal output
rlabel metal2 s 34610 119200 34666 120800 6 m_la_reset[2]
port 154 nsew signal output
rlabel metal2 s 34794 119200 34850 120800 6 m_la_reset[3]
port 155 nsew signal output
rlabel metal2 s 34978 119200 35034 120800 6 m_la_reset[4]
port 156 nsew signal output
rlabel metal2 s 35254 119200 35310 120800 6 m_la_reset[5]
port 157 nsew signal output
rlabel metal2 s 35438 119200 35494 120800 6 m_la_reset[6]
port 158 nsew signal output
rlabel metal2 s 35622 119200 35678 120800 6 m_la_reset[7]
port 159 nsew signal output
rlabel metal2 s 35806 119200 35862 120800 6 m_la_reset[8]
port 160 nsew signal output
rlabel metal2 s 36082 119200 36138 120800 6 m_la_reset[9]
port 161 nsew signal output
rlabel metal2 s 35438 -800 35494 800 8 m_wb_clk_i
port 162 nsew signal output
rlabel metal3 s -800 106224 800 106344 4 m_wb_rst_i
port 163 nsew signal output
rlabel metal3 s 39200 110576 40800 110696 6 m_wbs_ack_o[0]
port 164 nsew signal input
rlabel metal2 s 38290 -800 38346 800 8 m_wbs_ack_o[10]
port 165 nsew signal input
rlabel metal3 s 39200 116560 40800 116680 6 m_wbs_ack_o[11]
port 166 nsew signal input
rlabel metal3 s 39200 111800 40800 111920 6 m_wbs_ack_o[1]
port 167 nsew signal input
rlabel metal2 s 35714 -800 35770 800 8 m_wbs_ack_o[2]
port 168 nsew signal input
rlabel metal2 s 37094 119200 37150 120800 6 m_wbs_ack_o[3]
port 169 nsew signal input
rlabel metal2 s 36542 -800 36598 800 8 m_wbs_ack_o[4]
port 170 nsew signal input
rlabel metal3 s 39200 114384 40800 114504 6 m_wbs_ack_o[5]
port 171 nsew signal input
rlabel metal2 s 37738 119200 37794 120800 6 m_wbs_ack_o[6]
port 172 nsew signal input
rlabel metal3 s 39200 115336 40800 115456 6 m_wbs_ack_o[7]
port 173 nsew signal input
rlabel metal3 s -800 111256 800 111376 4 m_wbs_ack_o[8]
port 174 nsew signal input
rlabel metal3 s -800 112888 800 113008 4 m_wbs_ack_o[9]
port 175 nsew signal input
rlabel metal3 s 39200 110984 40800 111104 6 m_wbs_adr_i[0]
port 176 nsew signal output
rlabel metal3 s -800 114520 800 114640 4 m_wbs_adr_i[10]
port 177 nsew signal output
rlabel metal3 s 39200 116968 40800 117088 6 m_wbs_adr_i[11]
port 178 nsew signal output
rlabel metal3 s 39200 112208 40800 112328 6 m_wbs_adr_i[1]
port 179 nsew signal output
rlabel metal2 s 35990 -800 36046 800 8 m_wbs_adr_i[2]
port 180 nsew signal output
rlabel metal3 s 39200 112752 40800 112872 6 m_wbs_adr_i[3]
port 181 nsew signal output
rlabel metal2 s 36910 -800 36966 800 8 m_wbs_adr_i[4]
port 182 nsew signal output
rlabel metal2 s 37186 -800 37242 800 8 m_wbs_adr_i[5]
port 183 nsew signal output
rlabel metal2 s 37922 119200 37978 120800 6 m_wbs_adr_i[6]
port 184 nsew signal output
rlabel metal3 s 39200 115744 40800 115864 6 m_wbs_adr_i[7]
port 185 nsew signal output
rlabel metal2 s 38198 119200 38254 120800 6 m_wbs_adr_i[8]
port 186 nsew signal output
rlabel metal3 s -800 113704 800 113824 4 m_wbs_adr_i[9]
port 187 nsew signal output
rlabel metal3 s -800 107040 800 107160 4 m_wbs_cs_i[0]
port 188 nsew signal output
rlabel metal3 s -800 115336 800 115456 4 m_wbs_cs_i[10]
port 189 nsew signal output
rlabel metal2 s 38658 -800 38714 800 8 m_wbs_cs_i[11]
port 190 nsew signal output
rlabel metal3 s -800 107856 800 107976 4 m_wbs_cs_i[1]
port 191 nsew signal output
rlabel metal3 s -800 108672 800 108792 4 m_wbs_cs_i[2]
port 192 nsew signal output
rlabel metal3 s 39200 113160 40800 113280 6 m_wbs_cs_i[3]
port 193 nsew signal output
rlabel metal3 s 39200 113976 40800 114096 6 m_wbs_cs_i[4]
port 194 nsew signal output
rlabel metal3 s -800 109488 800 109608 4 m_wbs_cs_i[5]
port 195 nsew signal output
rlabel metal3 s 39200 114792 40800 114912 6 m_wbs_cs_i[6]
port 196 nsew signal output
rlabel metal2 s 37738 -800 37794 800 8 m_wbs_cs_i[7]
port 197 nsew signal output
rlabel metal3 s -800 112072 800 112192 4 m_wbs_cs_i[8]
port 198 nsew signal output
rlabel metal2 s 38014 -800 38070 800 8 m_wbs_cs_i[9]
port 199 nsew signal output
rlabel metal3 s 39200 111392 40800 111512 6 m_wbs_dat_i[0]
port 200 nsew signal output
rlabel metal3 s 39200 116152 40800 116272 6 m_wbs_dat_i[10]
port 201 nsew signal output
rlabel metal3 s -800 116152 800 116272 4 m_wbs_dat_i[11]
port 202 nsew signal output
rlabel metal2 s 38934 -800 38990 800 8 m_wbs_dat_i[12]
port 203 nsew signal output
rlabel metal3 s -800 116968 800 117088 4 m_wbs_dat_i[13]
port 204 nsew signal output
rlabel metal2 s 38842 119200 38898 120800 6 m_wbs_dat_i[14]
port 205 nsew signal output
rlabel metal3 s -800 117784 800 117904 4 m_wbs_dat_i[15]
port 206 nsew signal output
rlabel metal2 s 39026 119200 39082 120800 6 m_wbs_dat_i[16]
port 207 nsew signal output
rlabel metal3 s 39200 117376 40800 117496 6 m_wbs_dat_i[17]
port 208 nsew signal output
rlabel metal2 s 39210 119200 39266 120800 6 m_wbs_dat_i[18]
port 209 nsew signal output
rlabel metal2 s 39486 119200 39542 120800 6 m_wbs_dat_i[19]
port 210 nsew signal output
rlabel metal2 s 36910 119200 36966 120800 6 m_wbs_dat_i[1]
port 211 nsew signal output
rlabel metal3 s -800 118600 800 118720 4 m_wbs_dat_i[20]
port 212 nsew signal output
rlabel metal2 s 39210 -800 39266 800 8 m_wbs_dat_i[21]
port 213 nsew signal output
rlabel metal3 s 39200 117920 40800 118040 6 m_wbs_dat_i[22]
port 214 nsew signal output
rlabel metal3 s 39200 118328 40800 118448 6 m_wbs_dat_i[23]
port 215 nsew signal output
rlabel metal2 s 39486 -800 39542 800 8 m_wbs_dat_i[24]
port 216 nsew signal output
rlabel metal2 s 39670 119200 39726 120800 6 m_wbs_dat_i[25]
port 217 nsew signal output
rlabel metal3 s 39200 118736 40800 118856 6 m_wbs_dat_i[26]
port 218 nsew signal output
rlabel metal3 s 39200 119144 40800 119264 6 m_wbs_dat_i[27]
port 219 nsew signal output
rlabel metal3 s 39200 119552 40800 119672 6 m_wbs_dat_i[28]
port 220 nsew signal output
rlabel metal2 s 39854 119200 39910 120800 6 m_wbs_dat_i[29]
port 221 nsew signal output
rlabel metal2 s 36266 -800 36322 800 8 m_wbs_dat_i[2]
port 222 nsew signal output
rlabel metal3 s -800 119416 800 119536 4 m_wbs_dat_i[30]
port 223 nsew signal output
rlabel metal2 s 39762 -800 39818 800 8 m_wbs_dat_i[31]
port 224 nsew signal output
rlabel metal3 s 39200 113568 40800 113688 6 m_wbs_dat_i[3]
port 225 nsew signal output
rlabel metal2 s 37370 119200 37426 120800 6 m_wbs_dat_i[4]
port 226 nsew signal output
rlabel metal2 s 37554 119200 37610 120800 6 m_wbs_dat_i[5]
port 227 nsew signal output
rlabel metal2 s 37462 -800 37518 800 8 m_wbs_dat_i[6]
port 228 nsew signal output
rlabel metal3 s -800 110440 800 110560 4 m_wbs_dat_i[7]
port 229 nsew signal output
rlabel metal2 s 38382 119200 38438 120800 6 m_wbs_dat_i[8]
port 230 nsew signal output
rlabel metal2 s 38566 119200 38622 120800 6 m_wbs_dat_i[9]
port 231 nsew signal output
rlabel metal3 s 39200 144 40800 264 6 m_wbs_dat_o_0[0]
port 232 nsew signal input
rlabel metal3 s 39200 4360 40800 4480 6 m_wbs_dat_o_0[10]
port 233 nsew signal input
rlabel metal3 s 39200 4768 40800 4888 6 m_wbs_dat_o_0[11]
port 234 nsew signal input
rlabel metal3 s 39200 5312 40800 5432 6 m_wbs_dat_o_0[12]
port 235 nsew signal input
rlabel metal3 s 39200 5720 40800 5840 6 m_wbs_dat_o_0[13]
port 236 nsew signal input
rlabel metal3 s 39200 6128 40800 6248 6 m_wbs_dat_o_0[14]
port 237 nsew signal input
rlabel metal3 s 39200 6536 40800 6656 6 m_wbs_dat_o_0[15]
port 238 nsew signal input
rlabel metal3 s 39200 6944 40800 7064 6 m_wbs_dat_o_0[16]
port 239 nsew signal input
rlabel metal3 s 39200 7352 40800 7472 6 m_wbs_dat_o_0[17]
port 240 nsew signal input
rlabel metal3 s 39200 7896 40800 8016 6 m_wbs_dat_o_0[18]
port 241 nsew signal input
rlabel metal3 s 39200 8304 40800 8424 6 m_wbs_dat_o_0[19]
port 242 nsew signal input
rlabel metal3 s 39200 552 40800 672 6 m_wbs_dat_o_0[1]
port 243 nsew signal input
rlabel metal3 s 39200 8712 40800 8832 6 m_wbs_dat_o_0[20]
port 244 nsew signal input
rlabel metal3 s 39200 9120 40800 9240 6 m_wbs_dat_o_0[21]
port 245 nsew signal input
rlabel metal3 s 39200 9528 40800 9648 6 m_wbs_dat_o_0[22]
port 246 nsew signal input
rlabel metal3 s 39200 9936 40800 10056 6 m_wbs_dat_o_0[23]
port 247 nsew signal input
rlabel metal3 s 39200 10480 40800 10600 6 m_wbs_dat_o_0[24]
port 248 nsew signal input
rlabel metal3 s 39200 10888 40800 11008 6 m_wbs_dat_o_0[25]
port 249 nsew signal input
rlabel metal3 s 39200 11296 40800 11416 6 m_wbs_dat_o_0[26]
port 250 nsew signal input
rlabel metal3 s 39200 11704 40800 11824 6 m_wbs_dat_o_0[27]
port 251 nsew signal input
rlabel metal3 s 39200 12112 40800 12232 6 m_wbs_dat_o_0[28]
port 252 nsew signal input
rlabel metal3 s 39200 12656 40800 12776 6 m_wbs_dat_o_0[29]
port 253 nsew signal input
rlabel metal3 s 39200 960 40800 1080 6 m_wbs_dat_o_0[2]
port 254 nsew signal input
rlabel metal3 s 39200 13064 40800 13184 6 m_wbs_dat_o_0[30]
port 255 nsew signal input
rlabel metal3 s 39200 13472 40800 13592 6 m_wbs_dat_o_0[31]
port 256 nsew signal input
rlabel metal3 s 39200 1368 40800 1488 6 m_wbs_dat_o_0[3]
port 257 nsew signal input
rlabel metal3 s 39200 1776 40800 1896 6 m_wbs_dat_o_0[4]
port 258 nsew signal input
rlabel metal3 s 39200 2184 40800 2304 6 m_wbs_dat_o_0[5]
port 259 nsew signal input
rlabel metal3 s 39200 2728 40800 2848 6 m_wbs_dat_o_0[6]
port 260 nsew signal input
rlabel metal3 s 39200 3136 40800 3256 6 m_wbs_dat_o_0[7]
port 261 nsew signal input
rlabel metal3 s 39200 3544 40800 3664 6 m_wbs_dat_o_0[8]
port 262 nsew signal input
rlabel metal3 s 39200 3952 40800 4072 6 m_wbs_dat_o_0[9]
port 263 nsew signal input
rlabel metal3 s 39200 14288 40800 14408 6 m_wbs_dat_o_10[0]
port 264 nsew signal input
rlabel metal3 s 39200 27208 40800 27328 6 m_wbs_dat_o_10[10]
port 265 nsew signal input
rlabel metal3 s 39200 28568 40800 28688 6 m_wbs_dat_o_10[11]
port 266 nsew signal input
rlabel metal3 s 39200 29792 40800 29912 6 m_wbs_dat_o_10[12]
port 267 nsew signal input
rlabel metal3 s 39200 31152 40800 31272 6 m_wbs_dat_o_10[13]
port 268 nsew signal input
rlabel metal3 s 39200 32376 40800 32496 6 m_wbs_dat_o_10[14]
port 269 nsew signal input
rlabel metal3 s 39200 33736 40800 33856 6 m_wbs_dat_o_10[15]
port 270 nsew signal input
rlabel metal3 s 39200 34960 40800 35080 6 m_wbs_dat_o_10[16]
port 271 nsew signal input
rlabel metal3 s 39200 36320 40800 36440 6 m_wbs_dat_o_10[17]
port 272 nsew signal input
rlabel metal3 s 39200 37680 40800 37800 6 m_wbs_dat_o_10[18]
port 273 nsew signal input
rlabel metal3 s 39200 38904 40800 39024 6 m_wbs_dat_o_10[19]
port 274 nsew signal input
rlabel metal3 s 39200 15648 40800 15768 6 m_wbs_dat_o_10[1]
port 275 nsew signal input
rlabel metal3 s 39200 40264 40800 40384 6 m_wbs_dat_o_10[20]
port 276 nsew signal input
rlabel metal3 s 39200 41488 40800 41608 6 m_wbs_dat_o_10[21]
port 277 nsew signal input
rlabel metal3 s 39200 42848 40800 42968 6 m_wbs_dat_o_10[22]
port 278 nsew signal input
rlabel metal3 s 39200 44072 40800 44192 6 m_wbs_dat_o_10[23]
port 279 nsew signal input
rlabel metal3 s 39200 45432 40800 45552 6 m_wbs_dat_o_10[24]
port 280 nsew signal input
rlabel metal3 s 39200 46656 40800 46776 6 m_wbs_dat_o_10[25]
port 281 nsew signal input
rlabel metal3 s 39200 48016 40800 48136 6 m_wbs_dat_o_10[26]
port 282 nsew signal input
rlabel metal3 s 39200 49240 40800 49360 6 m_wbs_dat_o_10[27]
port 283 nsew signal input
rlabel metal3 s 39200 50600 40800 50720 6 m_wbs_dat_o_10[28]
port 284 nsew signal input
rlabel metal3 s 39200 51824 40800 51944 6 m_wbs_dat_o_10[29]
port 285 nsew signal input
rlabel metal3 s 39200 16872 40800 16992 6 m_wbs_dat_o_10[2]
port 286 nsew signal input
rlabel metal3 s 39200 53184 40800 53304 6 m_wbs_dat_o_10[30]
port 287 nsew signal input
rlabel metal3 s 39200 54408 40800 54528 6 m_wbs_dat_o_10[31]
port 288 nsew signal input
rlabel metal3 s 39200 18232 40800 18352 6 m_wbs_dat_o_10[3]
port 289 nsew signal input
rlabel metal3 s 39200 19456 40800 19576 6 m_wbs_dat_o_10[4]
port 290 nsew signal input
rlabel metal3 s 39200 20816 40800 20936 6 m_wbs_dat_o_10[5]
port 291 nsew signal input
rlabel metal3 s 39200 22040 40800 22160 6 m_wbs_dat_o_10[6]
port 292 nsew signal input
rlabel metal3 s 39200 23400 40800 23520 6 m_wbs_dat_o_10[7]
port 293 nsew signal input
rlabel metal3 s 39200 24624 40800 24744 6 m_wbs_dat_o_10[8]
port 294 nsew signal input
rlabel metal3 s 39200 25984 40800 26104 6 m_wbs_dat_o_10[9]
port 295 nsew signal input
rlabel metal3 s 39200 14696 40800 14816 6 m_wbs_dat_o_11[0]
port 296 nsew signal input
rlabel metal3 s 39200 27752 40800 27872 6 m_wbs_dat_o_11[10]
port 297 nsew signal input
rlabel metal3 s 39200 28976 40800 29096 6 m_wbs_dat_o_11[11]
port 298 nsew signal input
rlabel metal3 s 39200 30336 40800 30456 6 m_wbs_dat_o_11[12]
port 299 nsew signal input
rlabel metal3 s 39200 31560 40800 31680 6 m_wbs_dat_o_11[13]
port 300 nsew signal input
rlabel metal3 s 39200 32920 40800 33040 6 m_wbs_dat_o_11[14]
port 301 nsew signal input
rlabel metal3 s 39200 34144 40800 34264 6 m_wbs_dat_o_11[15]
port 302 nsew signal input
rlabel metal3 s 39200 35504 40800 35624 6 m_wbs_dat_o_11[16]
port 303 nsew signal input
rlabel metal3 s 39200 36728 40800 36848 6 m_wbs_dat_o_11[17]
port 304 nsew signal input
rlabel metal3 s 39200 38088 40800 38208 6 m_wbs_dat_o_11[18]
port 305 nsew signal input
rlabel metal3 s 39200 39312 40800 39432 6 m_wbs_dat_o_11[19]
port 306 nsew signal input
rlabel metal3 s 39200 16056 40800 16176 6 m_wbs_dat_o_11[1]
port 307 nsew signal input
rlabel metal3 s 39200 40672 40800 40792 6 m_wbs_dat_o_11[20]
port 308 nsew signal input
rlabel metal3 s 39200 41896 40800 42016 6 m_wbs_dat_o_11[21]
port 309 nsew signal input
rlabel metal3 s 39200 43256 40800 43376 6 m_wbs_dat_o_11[22]
port 310 nsew signal input
rlabel metal3 s 39200 44480 40800 44600 6 m_wbs_dat_o_11[23]
port 311 nsew signal input
rlabel metal3 s 39200 45840 40800 45960 6 m_wbs_dat_o_11[24]
port 312 nsew signal input
rlabel metal3 s 39200 47064 40800 47184 6 m_wbs_dat_o_11[25]
port 313 nsew signal input
rlabel metal3 s 39200 48424 40800 48544 6 m_wbs_dat_o_11[26]
port 314 nsew signal input
rlabel metal3 s 39200 49648 40800 49768 6 m_wbs_dat_o_11[27]
port 315 nsew signal input
rlabel metal3 s 39200 51008 40800 51128 6 m_wbs_dat_o_11[28]
port 316 nsew signal input
rlabel metal3 s 39200 52232 40800 52352 6 m_wbs_dat_o_11[29]
port 317 nsew signal input
rlabel metal3 s 39200 17280 40800 17400 6 m_wbs_dat_o_11[2]
port 318 nsew signal input
rlabel metal3 s 39200 53592 40800 53712 6 m_wbs_dat_o_11[30]
port 319 nsew signal input
rlabel metal3 s 39200 54816 40800 54936 6 m_wbs_dat_o_11[31]
port 320 nsew signal input
rlabel metal3 s 39200 18640 40800 18760 6 m_wbs_dat_o_11[3]
port 321 nsew signal input
rlabel metal3 s 39200 19864 40800 19984 6 m_wbs_dat_o_11[4]
port 322 nsew signal input
rlabel metal3 s 39200 21224 40800 21344 6 m_wbs_dat_o_11[5]
port 323 nsew signal input
rlabel metal3 s 39200 22448 40800 22568 6 m_wbs_dat_o_11[6]
port 324 nsew signal input
rlabel metal3 s 39200 23808 40800 23928 6 m_wbs_dat_o_11[7]
port 325 nsew signal input
rlabel metal3 s 39200 25168 40800 25288 6 m_wbs_dat_o_11[8]
port 326 nsew signal input
rlabel metal3 s 39200 26392 40800 26512 6 m_wbs_dat_o_11[9]
port 327 nsew signal input
rlabel metal3 s 39200 13880 40800 14000 6 m_wbs_dat_o_1[0]
port 328 nsew signal input
rlabel metal3 s 39200 26800 40800 26920 6 m_wbs_dat_o_1[10]
port 329 nsew signal input
rlabel metal3 s 39200 28160 40800 28280 6 m_wbs_dat_o_1[11]
port 330 nsew signal input
rlabel metal3 s 39200 29384 40800 29504 6 m_wbs_dat_o_1[12]
port 331 nsew signal input
rlabel metal3 s 39200 30744 40800 30864 6 m_wbs_dat_o_1[13]
port 332 nsew signal input
rlabel metal3 s 39200 31968 40800 32088 6 m_wbs_dat_o_1[14]
port 333 nsew signal input
rlabel metal3 s 39200 33328 40800 33448 6 m_wbs_dat_o_1[15]
port 334 nsew signal input
rlabel metal3 s 39200 34552 40800 34672 6 m_wbs_dat_o_1[16]
port 335 nsew signal input
rlabel metal3 s 39200 35912 40800 36032 6 m_wbs_dat_o_1[17]
port 336 nsew signal input
rlabel metal3 s 39200 37136 40800 37256 6 m_wbs_dat_o_1[18]
port 337 nsew signal input
rlabel metal3 s 39200 38496 40800 38616 6 m_wbs_dat_o_1[19]
port 338 nsew signal input
rlabel metal3 s 39200 15240 40800 15360 6 m_wbs_dat_o_1[1]
port 339 nsew signal input
rlabel metal3 s 39200 39720 40800 39840 6 m_wbs_dat_o_1[20]
port 340 nsew signal input
rlabel metal3 s 39200 41080 40800 41200 6 m_wbs_dat_o_1[21]
port 341 nsew signal input
rlabel metal3 s 39200 42304 40800 42424 6 m_wbs_dat_o_1[22]
port 342 nsew signal input
rlabel metal3 s 39200 43664 40800 43784 6 m_wbs_dat_o_1[23]
port 343 nsew signal input
rlabel metal3 s 39200 44888 40800 45008 6 m_wbs_dat_o_1[24]
port 344 nsew signal input
rlabel metal3 s 39200 46248 40800 46368 6 m_wbs_dat_o_1[25]
port 345 nsew signal input
rlabel metal3 s 39200 47472 40800 47592 6 m_wbs_dat_o_1[26]
port 346 nsew signal input
rlabel metal3 s 39200 48832 40800 48952 6 m_wbs_dat_o_1[27]
port 347 nsew signal input
rlabel metal3 s 39200 50192 40800 50312 6 m_wbs_dat_o_1[28]
port 348 nsew signal input
rlabel metal3 s 39200 51416 40800 51536 6 m_wbs_dat_o_1[29]
port 349 nsew signal input
rlabel metal3 s 39200 16464 40800 16584 6 m_wbs_dat_o_1[2]
port 350 nsew signal input
rlabel metal3 s 39200 52776 40800 52896 6 m_wbs_dat_o_1[30]
port 351 nsew signal input
rlabel metal3 s 39200 54000 40800 54120 6 m_wbs_dat_o_1[31]
port 352 nsew signal input
rlabel metal3 s 39200 17824 40800 17944 6 m_wbs_dat_o_1[3]
port 353 nsew signal input
rlabel metal3 s 39200 19048 40800 19168 6 m_wbs_dat_o_1[4]
port 354 nsew signal input
rlabel metal3 s 39200 20408 40800 20528 6 m_wbs_dat_o_1[5]
port 355 nsew signal input
rlabel metal3 s 39200 21632 40800 21752 6 m_wbs_dat_o_1[6]
port 356 nsew signal input
rlabel metal3 s 39200 22992 40800 23112 6 m_wbs_dat_o_1[7]
port 357 nsew signal input
rlabel metal3 s 39200 24216 40800 24336 6 m_wbs_dat_o_1[8]
port 358 nsew signal input
rlabel metal3 s 39200 25576 40800 25696 6 m_wbs_dat_o_1[9]
port 359 nsew signal input
rlabel metal3 s 39200 55360 40800 55480 6 m_wbs_dat_o_2[0]
port 360 nsew signal input
rlabel metal3 s 39200 59576 40800 59696 6 m_wbs_dat_o_2[10]
port 361 nsew signal input
rlabel metal3 s 39200 60120 40800 60240 6 m_wbs_dat_o_2[11]
port 362 nsew signal input
rlabel metal3 s 39200 60528 40800 60648 6 m_wbs_dat_o_2[12]
port 363 nsew signal input
rlabel metal3 s 39200 60936 40800 61056 6 m_wbs_dat_o_2[13]
port 364 nsew signal input
rlabel metal3 s 39200 61344 40800 61464 6 m_wbs_dat_o_2[14]
port 365 nsew signal input
rlabel metal3 s 39200 61752 40800 61872 6 m_wbs_dat_o_2[15]
port 366 nsew signal input
rlabel metal3 s 39200 62160 40800 62280 6 m_wbs_dat_o_2[16]
port 367 nsew signal input
rlabel metal3 s 39200 62704 40800 62824 6 m_wbs_dat_o_2[17]
port 368 nsew signal input
rlabel metal3 s 39200 63112 40800 63232 6 m_wbs_dat_o_2[18]
port 369 nsew signal input
rlabel metal3 s 39200 63520 40800 63640 6 m_wbs_dat_o_2[19]
port 370 nsew signal input
rlabel metal3 s 39200 55768 40800 55888 6 m_wbs_dat_o_2[1]
port 371 nsew signal input
rlabel metal3 s 39200 63928 40800 64048 6 m_wbs_dat_o_2[20]
port 372 nsew signal input
rlabel metal3 s 39200 64336 40800 64456 6 m_wbs_dat_o_2[21]
port 373 nsew signal input
rlabel metal3 s 39200 64744 40800 64864 6 m_wbs_dat_o_2[22]
port 374 nsew signal input
rlabel metal3 s 39200 65288 40800 65408 6 m_wbs_dat_o_2[23]
port 375 nsew signal input
rlabel metal3 s 39200 65696 40800 65816 6 m_wbs_dat_o_2[24]
port 376 nsew signal input
rlabel metal3 s 39200 66104 40800 66224 6 m_wbs_dat_o_2[25]
port 377 nsew signal input
rlabel metal3 s 39200 66512 40800 66632 6 m_wbs_dat_o_2[26]
port 378 nsew signal input
rlabel metal3 s 39200 66920 40800 67040 6 m_wbs_dat_o_2[27]
port 379 nsew signal input
rlabel metal3 s 39200 67328 40800 67448 6 m_wbs_dat_o_2[28]
port 380 nsew signal input
rlabel metal3 s 39200 67872 40800 67992 6 m_wbs_dat_o_2[29]
port 381 nsew signal input
rlabel metal3 s 39200 56176 40800 56296 6 m_wbs_dat_o_2[2]
port 382 nsew signal input
rlabel metal3 s 39200 68280 40800 68400 6 m_wbs_dat_o_2[30]
port 383 nsew signal input
rlabel metal3 s 39200 68688 40800 68808 6 m_wbs_dat_o_2[31]
port 384 nsew signal input
rlabel metal3 s 39200 56584 40800 56704 6 m_wbs_dat_o_2[3]
port 385 nsew signal input
rlabel metal3 s 39200 56992 40800 57112 6 m_wbs_dat_o_2[4]
port 386 nsew signal input
rlabel metal3 s 39200 57400 40800 57520 6 m_wbs_dat_o_2[5]
port 387 nsew signal input
rlabel metal3 s 39200 57944 40800 58064 6 m_wbs_dat_o_2[6]
port 388 nsew signal input
rlabel metal3 s 39200 58352 40800 58472 6 m_wbs_dat_o_2[7]
port 389 nsew signal input
rlabel metal3 s 39200 58760 40800 58880 6 m_wbs_dat_o_2[8]
port 390 nsew signal input
rlabel metal3 s 39200 59168 40800 59288 6 m_wbs_dat_o_2[9]
port 391 nsew signal input
rlabel metal3 s 39200 69096 40800 69216 6 m_wbs_dat_o_3[0]
port 392 nsew signal input
rlabel metal3 s 39200 73448 40800 73568 6 m_wbs_dat_o_3[10]
port 393 nsew signal input
rlabel metal3 s 39200 73856 40800 73976 6 m_wbs_dat_o_3[11]
port 394 nsew signal input
rlabel metal3 s 39200 74264 40800 74384 6 m_wbs_dat_o_3[12]
port 395 nsew signal input
rlabel metal3 s 39200 74672 40800 74792 6 m_wbs_dat_o_3[13]
port 396 nsew signal input
rlabel metal3 s 39200 75216 40800 75336 6 m_wbs_dat_o_3[14]
port 397 nsew signal input
rlabel metal3 s 39200 75624 40800 75744 6 m_wbs_dat_o_3[15]
port 398 nsew signal input
rlabel metal3 s 39200 76032 40800 76152 6 m_wbs_dat_o_3[16]
port 399 nsew signal input
rlabel metal3 s 39200 76440 40800 76560 6 m_wbs_dat_o_3[17]
port 400 nsew signal input
rlabel metal3 s 39200 76848 40800 76968 6 m_wbs_dat_o_3[18]
port 401 nsew signal input
rlabel metal3 s 39200 77256 40800 77376 6 m_wbs_dat_o_3[19]
port 402 nsew signal input
rlabel metal3 s 39200 69504 40800 69624 6 m_wbs_dat_o_3[1]
port 403 nsew signal input
rlabel metal3 s 39200 77800 40800 77920 6 m_wbs_dat_o_3[20]
port 404 nsew signal input
rlabel metal3 s 39200 78208 40800 78328 6 m_wbs_dat_o_3[21]
port 405 nsew signal input
rlabel metal3 s 39200 78616 40800 78736 6 m_wbs_dat_o_3[22]
port 406 nsew signal input
rlabel metal3 s 39200 79024 40800 79144 6 m_wbs_dat_o_3[23]
port 407 nsew signal input
rlabel metal3 s 39200 79432 40800 79552 6 m_wbs_dat_o_3[24]
port 408 nsew signal input
rlabel metal3 s 39200 79840 40800 79960 6 m_wbs_dat_o_3[25]
port 409 nsew signal input
rlabel metal3 s 39200 80384 40800 80504 6 m_wbs_dat_o_3[26]
port 410 nsew signal input
rlabel metal3 s 39200 80792 40800 80912 6 m_wbs_dat_o_3[27]
port 411 nsew signal input
rlabel metal3 s 39200 81200 40800 81320 6 m_wbs_dat_o_3[28]
port 412 nsew signal input
rlabel metal3 s 39200 81608 40800 81728 6 m_wbs_dat_o_3[29]
port 413 nsew signal input
rlabel metal3 s 39200 69912 40800 70032 6 m_wbs_dat_o_3[2]
port 414 nsew signal input
rlabel metal3 s 39200 82016 40800 82136 6 m_wbs_dat_o_3[30]
port 415 nsew signal input
rlabel metal3 s 39200 82424 40800 82544 6 m_wbs_dat_o_3[31]
port 416 nsew signal input
rlabel metal3 s 39200 70456 40800 70576 6 m_wbs_dat_o_3[3]
port 417 nsew signal input
rlabel metal3 s 39200 70864 40800 70984 6 m_wbs_dat_o_3[4]
port 418 nsew signal input
rlabel metal3 s 39200 71272 40800 71392 6 m_wbs_dat_o_3[5]
port 419 nsew signal input
rlabel metal3 s 39200 71680 40800 71800 6 m_wbs_dat_o_3[6]
port 420 nsew signal input
rlabel metal3 s 39200 72088 40800 72208 6 m_wbs_dat_o_3[7]
port 421 nsew signal input
rlabel metal3 s 39200 72632 40800 72752 6 m_wbs_dat_o_3[8]
port 422 nsew signal input
rlabel metal3 s 39200 73040 40800 73160 6 m_wbs_dat_o_3[9]
port 423 nsew signal input
rlabel metal3 s 39200 82968 40800 83088 6 m_wbs_dat_o_4[0]
port 424 nsew signal input
rlabel metal3 s 39200 87184 40800 87304 6 m_wbs_dat_o_4[10]
port 425 nsew signal input
rlabel metal3 s 39200 87728 40800 87848 6 m_wbs_dat_o_4[11]
port 426 nsew signal input
rlabel metal3 s 39200 88136 40800 88256 6 m_wbs_dat_o_4[12]
port 427 nsew signal input
rlabel metal3 s 39200 88544 40800 88664 6 m_wbs_dat_o_4[13]
port 428 nsew signal input
rlabel metal3 s 39200 88952 40800 89072 6 m_wbs_dat_o_4[14]
port 429 nsew signal input
rlabel metal3 s 39200 89360 40800 89480 6 m_wbs_dat_o_4[15]
port 430 nsew signal input
rlabel metal3 s 39200 89768 40800 89888 6 m_wbs_dat_o_4[16]
port 431 nsew signal input
rlabel metal3 s 39200 90312 40800 90432 6 m_wbs_dat_o_4[17]
port 432 nsew signal input
rlabel metal3 s 39200 90720 40800 90840 6 m_wbs_dat_o_4[18]
port 433 nsew signal input
rlabel metal3 s 39200 91128 40800 91248 6 m_wbs_dat_o_4[19]
port 434 nsew signal input
rlabel metal3 s 39200 83376 40800 83496 6 m_wbs_dat_o_4[1]
port 435 nsew signal input
rlabel metal3 s 39200 91536 40800 91656 6 m_wbs_dat_o_4[20]
port 436 nsew signal input
rlabel metal3 s 39200 91944 40800 92064 6 m_wbs_dat_o_4[21]
port 437 nsew signal input
rlabel metal3 s 39200 92352 40800 92472 6 m_wbs_dat_o_4[22]
port 438 nsew signal input
rlabel metal3 s 39200 92896 40800 93016 6 m_wbs_dat_o_4[23]
port 439 nsew signal input
rlabel metal3 s 39200 93304 40800 93424 6 m_wbs_dat_o_4[24]
port 440 nsew signal input
rlabel metal3 s 39200 93712 40800 93832 6 m_wbs_dat_o_4[25]
port 441 nsew signal input
rlabel metal3 s 39200 94120 40800 94240 6 m_wbs_dat_o_4[26]
port 442 nsew signal input
rlabel metal3 s 39200 94528 40800 94648 6 m_wbs_dat_o_4[27]
port 443 nsew signal input
rlabel metal3 s 39200 94936 40800 95056 6 m_wbs_dat_o_4[28]
port 444 nsew signal input
rlabel metal3 s 39200 95480 40800 95600 6 m_wbs_dat_o_4[29]
port 445 nsew signal input
rlabel metal3 s 39200 83784 40800 83904 6 m_wbs_dat_o_4[2]
port 446 nsew signal input
rlabel metal3 s 39200 95888 40800 96008 6 m_wbs_dat_o_4[30]
port 447 nsew signal input
rlabel metal3 s 39200 96296 40800 96416 6 m_wbs_dat_o_4[31]
port 448 nsew signal input
rlabel metal3 s 39200 84192 40800 84312 6 m_wbs_dat_o_4[3]
port 449 nsew signal input
rlabel metal3 s 39200 84600 40800 84720 6 m_wbs_dat_o_4[4]
port 450 nsew signal input
rlabel metal3 s 39200 85144 40800 85264 6 m_wbs_dat_o_4[5]
port 451 nsew signal input
rlabel metal3 s 39200 85552 40800 85672 6 m_wbs_dat_o_4[6]
port 452 nsew signal input
rlabel metal3 s 39200 85960 40800 86080 6 m_wbs_dat_o_4[7]
port 453 nsew signal input
rlabel metal3 s 39200 86368 40800 86488 6 m_wbs_dat_o_4[8]
port 454 nsew signal input
rlabel metal3 s 39200 86776 40800 86896 6 m_wbs_dat_o_4[9]
port 455 nsew signal input
rlabel metal3 s 39200 96704 40800 96824 6 m_wbs_dat_o_5[0]
port 456 nsew signal input
rlabel metal3 s 39200 101056 40800 101176 6 m_wbs_dat_o_5[10]
port 457 nsew signal input
rlabel metal3 s 39200 101464 40800 101584 6 m_wbs_dat_o_5[11]
port 458 nsew signal input
rlabel metal3 s 39200 101872 40800 101992 6 m_wbs_dat_o_5[12]
port 459 nsew signal input
rlabel metal3 s 39200 102280 40800 102400 6 m_wbs_dat_o_5[13]
port 460 nsew signal input
rlabel metal3 s 39200 102824 40800 102944 6 m_wbs_dat_o_5[14]
port 461 nsew signal input
rlabel metal3 s 39200 103232 40800 103352 6 m_wbs_dat_o_5[15]
port 462 nsew signal input
rlabel metal3 s 39200 103640 40800 103760 6 m_wbs_dat_o_5[16]
port 463 nsew signal input
rlabel metal3 s 39200 104048 40800 104168 6 m_wbs_dat_o_5[17]
port 464 nsew signal input
rlabel metal3 s 39200 104456 40800 104576 6 m_wbs_dat_o_5[18]
port 465 nsew signal input
rlabel metal3 s 39200 104864 40800 104984 6 m_wbs_dat_o_5[19]
port 466 nsew signal input
rlabel metal3 s 39200 97112 40800 97232 6 m_wbs_dat_o_5[1]
port 467 nsew signal input
rlabel metal3 s 39200 105408 40800 105528 6 m_wbs_dat_o_5[20]
port 468 nsew signal input
rlabel metal3 s 39200 105816 40800 105936 6 m_wbs_dat_o_5[21]
port 469 nsew signal input
rlabel metal3 s 39200 106224 40800 106344 6 m_wbs_dat_o_5[22]
port 470 nsew signal input
rlabel metal3 s 39200 106632 40800 106752 6 m_wbs_dat_o_5[23]
port 471 nsew signal input
rlabel metal3 s 39200 107040 40800 107160 6 m_wbs_dat_o_5[24]
port 472 nsew signal input
rlabel metal3 s 39200 107448 40800 107568 6 m_wbs_dat_o_5[25]
port 473 nsew signal input
rlabel metal3 s 39200 107992 40800 108112 6 m_wbs_dat_o_5[26]
port 474 nsew signal input
rlabel metal3 s 39200 108400 40800 108520 6 m_wbs_dat_o_5[27]
port 475 nsew signal input
rlabel metal3 s 39200 108808 40800 108928 6 m_wbs_dat_o_5[28]
port 476 nsew signal input
rlabel metal3 s 39200 109216 40800 109336 6 m_wbs_dat_o_5[29]
port 477 nsew signal input
rlabel metal3 s 39200 97656 40800 97776 6 m_wbs_dat_o_5[2]
port 478 nsew signal input
rlabel metal3 s 39200 109624 40800 109744 6 m_wbs_dat_o_5[30]
port 479 nsew signal input
rlabel metal3 s 39200 110168 40800 110288 6 m_wbs_dat_o_5[31]
port 480 nsew signal input
rlabel metal3 s 39200 98064 40800 98184 6 m_wbs_dat_o_5[3]
port 481 nsew signal input
rlabel metal3 s 39200 98472 40800 98592 6 m_wbs_dat_o_5[4]
port 482 nsew signal input
rlabel metal3 s 39200 98880 40800 99000 6 m_wbs_dat_o_5[5]
port 483 nsew signal input
rlabel metal3 s 39200 99288 40800 99408 6 m_wbs_dat_o_5[6]
port 484 nsew signal input
rlabel metal3 s 39200 99696 40800 99816 6 m_wbs_dat_o_5[7]
port 485 nsew signal input
rlabel metal3 s 39200 100240 40800 100360 6 m_wbs_dat_o_5[8]
port 486 nsew signal input
rlabel metal3 s 39200 100648 40800 100768 6 m_wbs_dat_o_5[9]
port 487 nsew signal input
rlabel metal3 s -800 416 800 536 4 m_wbs_dat_o_6[0]
port 488 nsew signal input
rlabel metal3 s -800 8576 800 8696 4 m_wbs_dat_o_6[10]
port 489 nsew signal input
rlabel metal3 s -800 9392 800 9512 4 m_wbs_dat_o_6[11]
port 490 nsew signal input
rlabel metal3 s -800 10208 800 10328 4 m_wbs_dat_o_6[12]
port 491 nsew signal input
rlabel metal3 s -800 11160 800 11280 4 m_wbs_dat_o_6[13]
port 492 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 m_wbs_dat_o_6[14]
port 493 nsew signal input
rlabel metal3 s -800 12792 800 12912 4 m_wbs_dat_o_6[15]
port 494 nsew signal input
rlabel metal3 s -800 13608 800 13728 4 m_wbs_dat_o_6[16]
port 495 nsew signal input
rlabel metal3 s -800 14424 800 14544 4 m_wbs_dat_o_6[17]
port 496 nsew signal input
rlabel metal3 s -800 15240 800 15360 4 m_wbs_dat_o_6[18]
port 497 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 m_wbs_dat_o_6[19]
port 498 nsew signal input
rlabel metal3 s -800 1232 800 1352 4 m_wbs_dat_o_6[1]
port 499 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 m_wbs_dat_o_6[20]
port 500 nsew signal input
rlabel metal3 s -800 17688 800 17808 4 m_wbs_dat_o_6[21]
port 501 nsew signal input
rlabel metal3 s -800 18504 800 18624 4 m_wbs_dat_o_6[22]
port 502 nsew signal input
rlabel metal3 s -800 19320 800 19440 4 m_wbs_dat_o_6[23]
port 503 nsew signal input
rlabel metal3 s -800 20136 800 20256 4 m_wbs_dat_o_6[24]
port 504 nsew signal input
rlabel metal3 s -800 21088 800 21208 4 m_wbs_dat_o_6[25]
port 505 nsew signal input
rlabel metal3 s -800 21904 800 22024 4 m_wbs_dat_o_6[26]
port 506 nsew signal input
rlabel metal3 s -800 22720 800 22840 4 m_wbs_dat_o_6[27]
port 507 nsew signal input
rlabel metal3 s -800 23536 800 23656 4 m_wbs_dat_o_6[28]
port 508 nsew signal input
rlabel metal3 s -800 24352 800 24472 4 m_wbs_dat_o_6[29]
port 509 nsew signal input
rlabel metal3 s -800 2048 800 2168 4 m_wbs_dat_o_6[2]
port 510 nsew signal input
rlabel metal3 s -800 25168 800 25288 4 m_wbs_dat_o_6[30]
port 511 nsew signal input
rlabel metal3 s -800 25984 800 26104 4 m_wbs_dat_o_6[31]
port 512 nsew signal input
rlabel metal3 s -800 2864 800 2984 4 m_wbs_dat_o_6[3]
port 513 nsew signal input
rlabel metal3 s -800 3680 800 3800 4 m_wbs_dat_o_6[4]
port 514 nsew signal input
rlabel metal3 s -800 4496 800 4616 4 m_wbs_dat_o_6[5]
port 515 nsew signal input
rlabel metal3 s -800 5312 800 5432 4 m_wbs_dat_o_6[6]
port 516 nsew signal input
rlabel metal3 s -800 6128 800 6248 4 m_wbs_dat_o_6[7]
port 517 nsew signal input
rlabel metal3 s -800 6944 800 7064 4 m_wbs_dat_o_6[8]
port 518 nsew signal input
rlabel metal3 s -800 7760 800 7880 4 m_wbs_dat_o_6[9]
port 519 nsew signal input
rlabel metal3 s -800 26800 800 26920 4 m_wbs_dat_o_7[0]
port 520 nsew signal input
rlabel metal3 s -800 35096 800 35216 4 m_wbs_dat_o_7[10]
port 521 nsew signal input
rlabel metal3 s -800 35912 800 36032 4 m_wbs_dat_o_7[11]
port 522 nsew signal input
rlabel metal3 s -800 36728 800 36848 4 m_wbs_dat_o_7[12]
port 523 nsew signal input
rlabel metal3 s -800 37544 800 37664 4 m_wbs_dat_o_7[13]
port 524 nsew signal input
rlabel metal3 s -800 38360 800 38480 4 m_wbs_dat_o_7[14]
port 525 nsew signal input
rlabel metal3 s -800 39176 800 39296 4 m_wbs_dat_o_7[15]
port 526 nsew signal input
rlabel metal3 s -800 39992 800 40112 4 m_wbs_dat_o_7[16]
port 527 nsew signal input
rlabel metal3 s -800 40944 800 41064 4 m_wbs_dat_o_7[17]
port 528 nsew signal input
rlabel metal3 s -800 41760 800 41880 4 m_wbs_dat_o_7[18]
port 529 nsew signal input
rlabel metal3 s -800 42576 800 42696 4 m_wbs_dat_o_7[19]
port 530 nsew signal input
rlabel metal3 s -800 27616 800 27736 4 m_wbs_dat_o_7[1]
port 531 nsew signal input
rlabel metal3 s -800 43392 800 43512 4 m_wbs_dat_o_7[20]
port 532 nsew signal input
rlabel metal3 s -800 44208 800 44328 4 m_wbs_dat_o_7[21]
port 533 nsew signal input
rlabel metal3 s -800 45024 800 45144 4 m_wbs_dat_o_7[22]
port 534 nsew signal input
rlabel metal3 s -800 45840 800 45960 4 m_wbs_dat_o_7[23]
port 535 nsew signal input
rlabel metal3 s -800 46656 800 46776 4 m_wbs_dat_o_7[24]
port 536 nsew signal input
rlabel metal3 s -800 47472 800 47592 4 m_wbs_dat_o_7[25]
port 537 nsew signal input
rlabel metal3 s -800 48288 800 48408 4 m_wbs_dat_o_7[26]
port 538 nsew signal input
rlabel metal3 s -800 49104 800 49224 4 m_wbs_dat_o_7[27]
port 539 nsew signal input
rlabel metal3 s -800 49920 800 50040 4 m_wbs_dat_o_7[28]
port 540 nsew signal input
rlabel metal3 s -800 50872 800 50992 4 m_wbs_dat_o_7[29]
port 541 nsew signal input
rlabel metal3 s -800 28432 800 28552 4 m_wbs_dat_o_7[2]
port 542 nsew signal input
rlabel metal3 s -800 51688 800 51808 4 m_wbs_dat_o_7[30]
port 543 nsew signal input
rlabel metal3 s -800 52504 800 52624 4 m_wbs_dat_o_7[31]
port 544 nsew signal input
rlabel metal3 s -800 29248 800 29368 4 m_wbs_dat_o_7[3]
port 545 nsew signal input
rlabel metal3 s -800 30064 800 30184 4 m_wbs_dat_o_7[4]
port 546 nsew signal input
rlabel metal3 s -800 31016 800 31136 4 m_wbs_dat_o_7[5]
port 547 nsew signal input
rlabel metal3 s -800 31832 800 31952 4 m_wbs_dat_o_7[6]
port 548 nsew signal input
rlabel metal3 s -800 32648 800 32768 4 m_wbs_dat_o_7[7]
port 549 nsew signal input
rlabel metal3 s -800 33464 800 33584 4 m_wbs_dat_o_7[8]
port 550 nsew signal input
rlabel metal3 s -800 34280 800 34400 4 m_wbs_dat_o_7[9]
port 551 nsew signal input
rlabel metal3 s -800 53320 800 53440 4 m_wbs_dat_o_8[0]
port 552 nsew signal input
rlabel metal3 s -800 61616 800 61736 4 m_wbs_dat_o_8[10]
port 553 nsew signal input
rlabel metal3 s -800 62432 800 62552 4 m_wbs_dat_o_8[11]
port 554 nsew signal input
rlabel metal3 s -800 63248 800 63368 4 m_wbs_dat_o_8[12]
port 555 nsew signal input
rlabel metal3 s -800 64064 800 64184 4 m_wbs_dat_o_8[13]
port 556 nsew signal input
rlabel metal3 s -800 64880 800 65000 4 m_wbs_dat_o_8[14]
port 557 nsew signal input
rlabel metal3 s -800 65696 800 65816 4 m_wbs_dat_o_8[15]
port 558 nsew signal input
rlabel metal3 s -800 66512 800 66632 4 m_wbs_dat_o_8[16]
port 559 nsew signal input
rlabel metal3 s -800 67328 800 67448 4 m_wbs_dat_o_8[17]
port 560 nsew signal input
rlabel metal3 s -800 68144 800 68264 4 m_wbs_dat_o_8[18]
port 561 nsew signal input
rlabel metal3 s -800 68960 800 69080 4 m_wbs_dat_o_8[19]
port 562 nsew signal input
rlabel metal3 s -800 54136 800 54256 4 m_wbs_dat_o_8[1]
port 563 nsew signal input
rlabel metal3 s -800 69776 800 69896 4 m_wbs_dat_o_8[20]
port 564 nsew signal input
rlabel metal3 s -800 70728 800 70848 4 m_wbs_dat_o_8[21]
port 565 nsew signal input
rlabel metal3 s -800 71544 800 71664 4 m_wbs_dat_o_8[22]
port 566 nsew signal input
rlabel metal3 s -800 72360 800 72480 4 m_wbs_dat_o_8[23]
port 567 nsew signal input
rlabel metal3 s -800 73176 800 73296 4 m_wbs_dat_o_8[24]
port 568 nsew signal input
rlabel metal3 s -800 73992 800 74112 4 m_wbs_dat_o_8[25]
port 569 nsew signal input
rlabel metal3 s -800 74808 800 74928 4 m_wbs_dat_o_8[26]
port 570 nsew signal input
rlabel metal3 s -800 75624 800 75744 4 m_wbs_dat_o_8[27]
port 571 nsew signal input
rlabel metal3 s -800 76440 800 76560 4 m_wbs_dat_o_8[28]
port 572 nsew signal input
rlabel metal3 s -800 77256 800 77376 4 m_wbs_dat_o_8[29]
port 573 nsew signal input
rlabel metal3 s -800 54952 800 55072 4 m_wbs_dat_o_8[2]
port 574 nsew signal input
rlabel metal3 s -800 78072 800 78192 4 m_wbs_dat_o_8[30]
port 575 nsew signal input
rlabel metal3 s -800 78888 800 79008 4 m_wbs_dat_o_8[31]
port 576 nsew signal input
rlabel metal3 s -800 55768 800 55888 4 m_wbs_dat_o_8[3]
port 577 nsew signal input
rlabel metal3 s -800 56584 800 56704 4 m_wbs_dat_o_8[4]
port 578 nsew signal input
rlabel metal3 s -800 57400 800 57520 4 m_wbs_dat_o_8[5]
port 579 nsew signal input
rlabel metal3 s -800 58216 800 58336 4 m_wbs_dat_o_8[6]
port 580 nsew signal input
rlabel metal3 s -800 59032 800 59152 4 m_wbs_dat_o_8[7]
port 581 nsew signal input
rlabel metal3 s -800 59848 800 59968 4 m_wbs_dat_o_8[8]
port 582 nsew signal input
rlabel metal3 s -800 60800 800 60920 4 m_wbs_dat_o_8[9]
port 583 nsew signal input
rlabel metal3 s -800 79704 800 79824 4 m_wbs_dat_o_9[0]
port 584 nsew signal input
rlabel metal3 s -800 88000 800 88120 4 m_wbs_dat_o_9[10]
port 585 nsew signal input
rlabel metal3 s -800 88816 800 88936 4 m_wbs_dat_o_9[11]
port 586 nsew signal input
rlabel metal3 s -800 89632 800 89752 4 m_wbs_dat_o_9[12]
port 587 nsew signal input
rlabel metal3 s -800 90584 800 90704 4 m_wbs_dat_o_9[13]
port 588 nsew signal input
rlabel metal3 s -800 91400 800 91520 4 m_wbs_dat_o_9[14]
port 589 nsew signal input
rlabel metal3 s -800 92216 800 92336 4 m_wbs_dat_o_9[15]
port 590 nsew signal input
rlabel metal3 s -800 93032 800 93152 4 m_wbs_dat_o_9[16]
port 591 nsew signal input
rlabel metal3 s -800 93848 800 93968 4 m_wbs_dat_o_9[17]
port 592 nsew signal input
rlabel metal3 s -800 94664 800 94784 4 m_wbs_dat_o_9[18]
port 593 nsew signal input
rlabel metal3 s -800 95480 800 95600 4 m_wbs_dat_o_9[19]
port 594 nsew signal input
rlabel metal3 s -800 80656 800 80776 4 m_wbs_dat_o_9[1]
port 595 nsew signal input
rlabel metal3 s -800 96296 800 96416 4 m_wbs_dat_o_9[20]
port 596 nsew signal input
rlabel metal3 s -800 97112 800 97232 4 m_wbs_dat_o_9[21]
port 597 nsew signal input
rlabel metal3 s -800 97928 800 98048 4 m_wbs_dat_o_9[22]
port 598 nsew signal input
rlabel metal3 s -800 98744 800 98864 4 m_wbs_dat_o_9[23]
port 599 nsew signal input
rlabel metal3 s -800 99560 800 99680 4 m_wbs_dat_o_9[24]
port 600 nsew signal input
rlabel metal3 s -800 100512 800 100632 4 m_wbs_dat_o_9[25]
port 601 nsew signal input
rlabel metal3 s -800 101328 800 101448 4 m_wbs_dat_o_9[26]
port 602 nsew signal input
rlabel metal3 s -800 102144 800 102264 4 m_wbs_dat_o_9[27]
port 603 nsew signal input
rlabel metal3 s -800 102960 800 103080 4 m_wbs_dat_o_9[28]
port 604 nsew signal input
rlabel metal3 s -800 103776 800 103896 4 m_wbs_dat_o_9[29]
port 605 nsew signal input
rlabel metal3 s -800 81472 800 81592 4 m_wbs_dat_o_9[2]
port 606 nsew signal input
rlabel metal3 s -800 104592 800 104712 4 m_wbs_dat_o_9[30]
port 607 nsew signal input
rlabel metal3 s -800 105408 800 105528 4 m_wbs_dat_o_9[31]
port 608 nsew signal input
rlabel metal3 s -800 82288 800 82408 4 m_wbs_dat_o_9[3]
port 609 nsew signal input
rlabel metal3 s -800 83104 800 83224 4 m_wbs_dat_o_9[4]
port 610 nsew signal input
rlabel metal3 s -800 83920 800 84040 4 m_wbs_dat_o_9[5]
port 611 nsew signal input
rlabel metal3 s -800 84736 800 84856 4 m_wbs_dat_o_9[6]
port 612 nsew signal input
rlabel metal3 s -800 85552 800 85672 4 m_wbs_dat_o_9[7]
port 613 nsew signal input
rlabel metal3 s -800 86368 800 86488 4 m_wbs_dat_o_9[8]
port 614 nsew signal input
rlabel metal3 s -800 87184 800 87304 4 m_wbs_dat_o_9[9]
port 615 nsew signal input
rlabel metal2 s 36726 119200 36782 120800 6 m_wbs_we_i
port 616 nsew signal output
rlabel metal2 s 25870 119200 25926 120800 6 mt_QEI_ChA_0
port 617 nsew signal output
rlabel metal2 s 26146 119200 26202 120800 6 mt_QEI_ChA_1
port 618 nsew signal output
rlabel metal2 s 26330 119200 26386 120800 6 mt_QEI_ChA_2
port 619 nsew signal output
rlabel metal2 s 26514 119200 26570 120800 6 mt_QEI_ChA_3
port 620 nsew signal output
rlabel metal2 s 26790 119200 26846 120800 6 mt_QEI_ChB_0
port 621 nsew signal output
rlabel metal2 s 26974 119200 27030 120800 6 mt_QEI_ChB_1
port 622 nsew signal output
rlabel metal2 s 27158 119200 27214 120800 6 mt_QEI_ChB_2
port 623 nsew signal output
rlabel metal2 s 27342 119200 27398 120800 6 mt_QEI_ChB_3
port 624 nsew signal output
rlabel metal2 s 27618 119200 27674 120800 6 mt_clo_test
port 625 nsew signal output
rlabel metal2 s 27802 119200 27858 120800 6 mt_pwm_h_0
port 626 nsew signal input
rlabel metal2 s 27986 119200 28042 120800 6 mt_pwm_h_1
port 627 nsew signal input
rlabel metal2 s 28262 119200 28318 120800 6 mt_pwm_h_2
port 628 nsew signal input
rlabel metal2 s 28446 119200 28502 120800 6 mt_pwm_h_3
port 629 nsew signal input
rlabel metal2 s 28630 119200 28686 120800 6 mt_pwm_l_0
port 630 nsew signal input
rlabel metal2 s 28906 119200 28962 120800 6 mt_pwm_l_1
port 631 nsew signal input
rlabel metal2 s 29090 119200 29146 120800 6 mt_pwm_l_2
port 632 nsew signal input
rlabel metal2 s 29274 119200 29330 120800 6 mt_pwm_l_3
port 633 nsew signal input
rlabel metal2 s 29458 119200 29514 120800 6 mt_pwm_test
port 634 nsew signal output
rlabel metal2 s 29918 119200 29974 120800 6 mt_sync_in[0]
port 635 nsew signal input
rlabel metal2 s 30102 119200 30158 120800 6 mt_sync_in[1]
port 636 nsew signal input
rlabel metal2 s 30378 119200 30434 120800 6 mt_sync_in[2]
port 637 nsew signal input
rlabel metal2 s 30562 119200 30618 120800 6 mt_sync_in[3]
port 638 nsew signal input
rlabel metal2 s 30746 119200 30802 120800 6 mt_sync_in[4]
port 639 nsew signal input
rlabel metal2 s 31022 119200 31078 120800 6 mt_sync_in[5]
port 640 nsew signal input
rlabel metal2 s 31206 119200 31262 120800 6 mt_sync_in[6]
port 641 nsew signal input
rlabel metal2 s 31390 119200 31446 120800 6 mt_sync_in[7]
port 642 nsew signal input
rlabel metal2 s 29734 119200 29790 120800 6 mt_sync_out
port 643 nsew signal output
rlabel metal2 s 110 -800 166 800 8 wb_clk_i
port 644 nsew signal input
rlabel metal2 s 386 -800 442 800 8 wb_rst_i
port 645 nsew signal input
rlabel metal2 s 1490 -800 1546 800 8 wbs_ack_o
port 646 nsew signal output
rlabel metal2 s 2686 -800 2742 800 8 wbs_adr_i[0]
port 647 nsew signal input
rlabel metal2 s 12622 -800 12678 800 8 wbs_adr_i[10]
port 648 nsew signal input
rlabel metal2 s 13542 -800 13598 800 8 wbs_adr_i[11]
port 649 nsew signal input
rlabel metal2 s 14370 -800 14426 800 8 wbs_adr_i[12]
port 650 nsew signal input
rlabel metal2 s 15290 -800 15346 800 8 wbs_adr_i[13]
port 651 nsew signal input
rlabel metal2 s 16118 -800 16174 800 8 wbs_adr_i[14]
port 652 nsew signal input
rlabel metal2 s 17038 -800 17094 800 8 wbs_adr_i[15]
port 653 nsew signal input
rlabel metal2 s 17866 -800 17922 800 8 wbs_adr_i[16]
port 654 nsew signal input
rlabel metal2 s 18786 -800 18842 800 8 wbs_adr_i[17]
port 655 nsew signal input
rlabel metal2 s 19614 -800 19670 800 8 wbs_adr_i[18]
port 656 nsew signal input
rlabel metal2 s 20534 -800 20590 800 8 wbs_adr_i[19]
port 657 nsew signal input
rlabel metal2 s 3882 -800 3938 800 8 wbs_adr_i[1]
port 658 nsew signal input
rlabel metal2 s 21362 -800 21418 800 8 wbs_adr_i[20]
port 659 nsew signal input
rlabel metal2 s 22282 -800 22338 800 8 wbs_adr_i[21]
port 660 nsew signal input
rlabel metal2 s 23110 -800 23166 800 8 wbs_adr_i[22]
port 661 nsew signal input
rlabel metal2 s 24030 -800 24086 800 8 wbs_adr_i[23]
port 662 nsew signal input
rlabel metal2 s 24858 -800 24914 800 8 wbs_adr_i[24]
port 663 nsew signal input
rlabel metal2 s 25778 -800 25834 800 8 wbs_adr_i[25]
port 664 nsew signal input
rlabel metal2 s 26606 -800 26662 800 8 wbs_adr_i[26]
port 665 nsew signal input
rlabel metal2 s 27526 -800 27582 800 8 wbs_adr_i[27]
port 666 nsew signal input
rlabel metal2 s 28354 -800 28410 800 8 wbs_adr_i[28]
port 667 nsew signal input
rlabel metal2 s 29274 -800 29330 800 8 wbs_adr_i[29]
port 668 nsew signal input
rlabel metal2 s 4986 -800 5042 800 8 wbs_adr_i[2]
port 669 nsew signal input
rlabel metal2 s 30194 -800 30250 800 8 wbs_adr_i[30]
port 670 nsew signal input
rlabel metal2 s 31022 -800 31078 800 8 wbs_adr_i[31]
port 671 nsew signal input
rlabel metal2 s 6182 -800 6238 800 8 wbs_adr_i[3]
port 672 nsew signal input
rlabel metal2 s 7378 -800 7434 800 8 wbs_adr_i[4]
port 673 nsew signal input
rlabel metal2 s 8206 -800 8262 800 8 wbs_adr_i[5]
port 674 nsew signal input
rlabel metal2 s 9126 -800 9182 800 8 wbs_adr_i[6]
port 675 nsew signal input
rlabel metal2 s 9954 -800 10010 800 8 wbs_adr_i[7]
port 676 nsew signal input
rlabel metal2 s 10874 -800 10930 800 8 wbs_adr_i[8]
port 677 nsew signal input
rlabel metal2 s 11794 -800 11850 800 8 wbs_adr_i[9]
port 678 nsew signal input
rlabel metal2 s 1858 -800 1914 800 8 wbs_cyc_i
port 679 nsew signal input
rlabel metal2 s 2962 -800 3018 800 8 wbs_dat_i[0]
port 680 nsew signal input
rlabel metal2 s 12898 -800 12954 800 8 wbs_dat_i[10]
port 681 nsew signal input
rlabel metal2 s 13818 -800 13874 800 8 wbs_dat_i[11]
port 682 nsew signal input
rlabel metal2 s 14646 -800 14702 800 8 wbs_dat_i[12]
port 683 nsew signal input
rlabel metal2 s 15566 -800 15622 800 8 wbs_dat_i[13]
port 684 nsew signal input
rlabel metal2 s 16394 -800 16450 800 8 wbs_dat_i[14]
port 685 nsew signal input
rlabel metal2 s 17314 -800 17370 800 8 wbs_dat_i[15]
port 686 nsew signal input
rlabel metal2 s 18142 -800 18198 800 8 wbs_dat_i[16]
port 687 nsew signal input
rlabel metal2 s 19062 -800 19118 800 8 wbs_dat_i[17]
port 688 nsew signal input
rlabel metal2 s 19890 -800 19946 800 8 wbs_dat_i[18]
port 689 nsew signal input
rlabel metal2 s 20810 -800 20866 800 8 wbs_dat_i[19]
port 690 nsew signal input
rlabel metal2 s 4158 -800 4214 800 8 wbs_dat_i[1]
port 691 nsew signal input
rlabel metal2 s 21638 -800 21694 800 8 wbs_dat_i[20]
port 692 nsew signal input
rlabel metal2 s 22558 -800 22614 800 8 wbs_dat_i[21]
port 693 nsew signal input
rlabel metal2 s 23478 -800 23534 800 8 wbs_dat_i[22]
port 694 nsew signal input
rlabel metal2 s 24306 -800 24362 800 8 wbs_dat_i[23]
port 695 nsew signal input
rlabel metal2 s 25226 -800 25282 800 8 wbs_dat_i[24]
port 696 nsew signal input
rlabel metal2 s 26054 -800 26110 800 8 wbs_dat_i[25]
port 697 nsew signal input
rlabel metal2 s 26974 -800 27030 800 8 wbs_dat_i[26]
port 698 nsew signal input
rlabel metal2 s 27802 -800 27858 800 8 wbs_dat_i[27]
port 699 nsew signal input
rlabel metal2 s 28722 -800 28778 800 8 wbs_dat_i[28]
port 700 nsew signal input
rlabel metal2 s 29550 -800 29606 800 8 wbs_dat_i[29]
port 701 nsew signal input
rlabel metal2 s 5354 -800 5410 800 8 wbs_dat_i[2]
port 702 nsew signal input
rlabel metal2 s 30470 -800 30526 800 8 wbs_dat_i[30]
port 703 nsew signal input
rlabel metal2 s 31298 -800 31354 800 8 wbs_dat_i[31]
port 704 nsew signal input
rlabel metal2 s 6458 -800 6514 800 8 wbs_dat_i[3]
port 705 nsew signal input
rlabel metal2 s 7654 -800 7710 800 8 wbs_dat_i[4]
port 706 nsew signal input
rlabel metal2 s 8574 -800 8630 800 8 wbs_dat_i[5]
port 707 nsew signal input
rlabel metal2 s 9402 -800 9458 800 8 wbs_dat_i[6]
port 708 nsew signal input
rlabel metal2 s 10322 -800 10378 800 8 wbs_dat_i[7]
port 709 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 wbs_dat_i[8]
port 710 nsew signal input
rlabel metal2 s 12070 -800 12126 800 8 wbs_dat_i[9]
port 711 nsew signal input
rlabel metal2 s 3238 -800 3294 800 8 wbs_dat_o[0]
port 712 nsew signal output
rlabel metal2 s 13174 -800 13230 800 8 wbs_dat_o[10]
port 713 nsew signal output
rlabel metal2 s 14094 -800 14150 800 8 wbs_dat_o[11]
port 714 nsew signal output
rlabel metal2 s 14922 -800 14978 800 8 wbs_dat_o[12]
port 715 nsew signal output
rlabel metal2 s 15842 -800 15898 800 8 wbs_dat_o[13]
port 716 nsew signal output
rlabel metal2 s 16670 -800 16726 800 8 wbs_dat_o[14]
port 717 nsew signal output
rlabel metal2 s 17590 -800 17646 800 8 wbs_dat_o[15]
port 718 nsew signal output
rlabel metal2 s 18510 -800 18566 800 8 wbs_dat_o[16]
port 719 nsew signal output
rlabel metal2 s 19338 -800 19394 800 8 wbs_dat_o[17]
port 720 nsew signal output
rlabel metal2 s 20258 -800 20314 800 8 wbs_dat_o[18]
port 721 nsew signal output
rlabel metal2 s 21086 -800 21142 800 8 wbs_dat_o[19]
port 722 nsew signal output
rlabel metal2 s 4434 -800 4490 800 8 wbs_dat_o[1]
port 723 nsew signal output
rlabel metal2 s 22006 -800 22062 800 8 wbs_dat_o[20]
port 724 nsew signal output
rlabel metal2 s 22834 -800 22890 800 8 wbs_dat_o[21]
port 725 nsew signal output
rlabel metal2 s 23754 -800 23810 800 8 wbs_dat_o[22]
port 726 nsew signal output
rlabel metal2 s 24582 -800 24638 800 8 wbs_dat_o[23]
port 727 nsew signal output
rlabel metal2 s 25502 -800 25558 800 8 wbs_dat_o[24]
port 728 nsew signal output
rlabel metal2 s 26330 -800 26386 800 8 wbs_dat_o[25]
port 729 nsew signal output
rlabel metal2 s 27250 -800 27306 800 8 wbs_dat_o[26]
port 730 nsew signal output
rlabel metal2 s 28078 -800 28134 800 8 wbs_dat_o[27]
port 731 nsew signal output
rlabel metal2 s 28998 -800 29054 800 8 wbs_dat_o[28]
port 732 nsew signal output
rlabel metal2 s 29826 -800 29882 800 8 wbs_dat_o[29]
port 733 nsew signal output
rlabel metal2 s 5630 -800 5686 800 8 wbs_dat_o[2]
port 734 nsew signal output
rlabel metal2 s 30746 -800 30802 800 8 wbs_dat_o[30]
port 735 nsew signal output
rlabel metal2 s 31574 -800 31630 800 8 wbs_dat_o[31]
port 736 nsew signal output
rlabel metal2 s 6826 -800 6882 800 8 wbs_dat_o[3]
port 737 nsew signal output
rlabel metal2 s 7930 -800 7986 800 8 wbs_dat_o[4]
port 738 nsew signal output
rlabel metal2 s 8850 -800 8906 800 8 wbs_dat_o[5]
port 739 nsew signal output
rlabel metal2 s 9678 -800 9734 800 8 wbs_dat_o[6]
port 740 nsew signal output
rlabel metal2 s 10598 -800 10654 800 8 wbs_dat_o[7]
port 741 nsew signal output
rlabel metal2 s 11426 -800 11482 800 8 wbs_dat_o[8]
port 742 nsew signal output
rlabel metal2 s 12346 -800 12402 800 8 wbs_dat_o[9]
port 743 nsew signal output
rlabel metal2 s 3606 -800 3662 800 8 wbs_sel_i[0]
port 744 nsew signal input
rlabel metal2 s 4710 -800 4766 800 8 wbs_sel_i[1]
port 745 nsew signal input
rlabel metal2 s 5906 -800 5962 800 8 wbs_sel_i[2]
port 746 nsew signal input
rlabel metal2 s 7102 -800 7158 800 8 wbs_sel_i[3]
port 747 nsew signal input
rlabel metal2 s 2134 -800 2190 800 8 wbs_stb_i
port 748 nsew signal input
rlabel metal2 s 2410 -800 2466 800 8 wbs_we_i
port 749 nsew signal input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 750 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 751 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 752 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 40000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/wb_local/runs/wb_local/results/magic/wb_local.gds
string GDS_END 4674038
string GDS_START 332948
<< end >>

