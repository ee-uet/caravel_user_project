magic
tech sky130A
magscale 1 2
timestamp 1624043987
<< obsli1 >>
rect 1104 2159 58880 117521
<< obsm1 >>
rect 1104 2128 58880 117552
<< metal2 >>
rect 3698 119200 3754 120800
rect 11150 119200 11206 120800
rect 18694 119200 18750 120800
rect 26146 119200 26202 120800
rect 33690 119200 33746 120800
rect 41142 119200 41198 120800
rect 48686 119200 48742 120800
rect 56138 119200 56194 120800
rect 4986 -800 5042 800
rect 14922 -800 14978 800
rect 24950 -800 25006 800
rect 34978 -800 35034 800
rect 44914 -800 44970 800
rect 54942 -800 54998 800
<< obsm2 >>
rect 1768 119144 3642 119200
rect 3810 119144 11094 119200
rect 11262 119144 18638 119200
rect 18806 119144 26090 119200
rect 26258 119144 33634 119200
rect 33802 119144 41086 119200
rect 41254 119144 48630 119200
rect 48798 119144 56082 119200
rect 56250 119144 58218 119200
rect 1768 856 58218 119144
rect 1768 800 4930 856
rect 5098 800 14866 856
rect 15034 800 24894 856
rect 25062 800 34922 856
rect 35090 800 44858 856
rect 45026 800 54886 856
rect 55054 800 58218 856
<< metal3 >>
rect 59200 118464 60800 118584
rect -800 117920 800 118040
rect 59200 115744 60800 115864
rect -800 114112 800 114232
rect 59200 113024 60800 113144
rect -800 110440 800 110560
rect 59200 110304 60800 110424
rect 59200 107584 60800 107704
rect -800 106632 800 106752
rect 59200 104864 60800 104984
rect -800 102960 800 103080
rect 59200 102144 60800 102264
rect 59200 99424 60800 99544
rect -800 99152 800 99272
rect 59200 96704 60800 96824
rect -800 95480 800 95600
rect 59200 93984 60800 94104
rect -800 91672 800 91792
rect 59200 91264 60800 91384
rect 59200 88544 60800 88664
rect -800 87864 800 87984
rect 59200 85824 60800 85944
rect -800 84192 800 84312
rect 59200 83104 60800 83224
rect -800 80384 800 80504
rect 59200 80384 60800 80504
rect 59200 77664 60800 77784
rect -800 76712 800 76832
rect 59200 74944 60800 75064
rect -800 72904 800 73024
rect 59200 72224 60800 72344
rect 59200 69504 60800 69624
rect -800 69232 800 69352
rect 59200 66784 60800 66904
rect -800 65424 800 65544
rect 59200 64064 60800 64184
rect -800 61752 800 61872
rect 59200 61344 60800 61464
rect 59200 58488 60800 58608
rect -800 57944 800 58064
rect 59200 55768 60800 55888
rect -800 54136 800 54256
rect 59200 53048 60800 53168
rect -800 50464 800 50584
rect 59200 50328 60800 50448
rect 59200 47608 60800 47728
rect -800 46656 800 46776
rect 59200 44888 60800 45008
rect -800 42984 800 43104
rect 59200 42168 60800 42288
rect 59200 39448 60800 39568
rect -800 39176 800 39296
rect 59200 36728 60800 36848
rect -800 35504 800 35624
rect 59200 34008 60800 34128
rect -800 31696 800 31816
rect 59200 31288 60800 31408
rect 59200 28568 60800 28688
rect -800 27888 800 28008
rect 59200 25848 60800 25968
rect -800 24216 800 24336
rect 59200 23128 60800 23248
rect -800 20408 800 20528
rect 59200 20408 60800 20528
rect 59200 17688 60800 17808
rect -800 16736 800 16856
rect 59200 14968 60800 15088
rect -800 12928 800 13048
rect 59200 12248 60800 12368
rect 59200 9528 60800 9648
rect -800 9256 800 9376
rect 59200 6808 60800 6928
rect -800 5448 800 5568
rect 59200 4088 60800 4208
rect -800 1776 800 1896
rect 59200 1368 60800 1488
<< obsm3 >>
rect 800 118384 59120 118557
rect 800 118120 59200 118384
rect 880 117840 59200 118120
rect 800 115944 59200 117840
rect 800 115664 59120 115944
rect 800 114312 59200 115664
rect 880 114032 59200 114312
rect 800 113224 59200 114032
rect 800 112944 59120 113224
rect 800 110640 59200 112944
rect 880 110504 59200 110640
rect 880 110360 59120 110504
rect 800 110224 59120 110360
rect 800 107784 59200 110224
rect 800 107504 59120 107784
rect 800 106832 59200 107504
rect 880 106552 59200 106832
rect 800 105064 59200 106552
rect 800 104784 59120 105064
rect 800 103160 59200 104784
rect 880 102880 59200 103160
rect 800 102344 59200 102880
rect 800 102064 59120 102344
rect 800 99624 59200 102064
rect 800 99352 59120 99624
rect 880 99344 59120 99352
rect 880 99072 59200 99344
rect 800 96904 59200 99072
rect 800 96624 59120 96904
rect 800 95680 59200 96624
rect 880 95400 59200 95680
rect 800 94184 59200 95400
rect 800 93904 59120 94184
rect 800 91872 59200 93904
rect 880 91592 59200 91872
rect 800 91464 59200 91592
rect 800 91184 59120 91464
rect 800 88744 59200 91184
rect 800 88464 59120 88744
rect 800 88064 59200 88464
rect 880 87784 59200 88064
rect 800 86024 59200 87784
rect 800 85744 59120 86024
rect 800 84392 59200 85744
rect 880 84112 59200 84392
rect 800 83304 59200 84112
rect 800 83024 59120 83304
rect 800 80584 59200 83024
rect 880 80304 59120 80584
rect 800 77864 59200 80304
rect 800 77584 59120 77864
rect 800 76912 59200 77584
rect 880 76632 59200 76912
rect 800 75144 59200 76632
rect 800 74864 59120 75144
rect 800 73104 59200 74864
rect 880 72824 59200 73104
rect 800 72424 59200 72824
rect 800 72144 59120 72424
rect 800 69704 59200 72144
rect 800 69432 59120 69704
rect 880 69424 59120 69432
rect 880 69152 59200 69424
rect 800 66984 59200 69152
rect 800 66704 59120 66984
rect 800 65624 59200 66704
rect 880 65344 59200 65624
rect 800 64264 59200 65344
rect 800 63984 59120 64264
rect 800 61952 59200 63984
rect 880 61672 59200 61952
rect 800 61544 59200 61672
rect 800 61264 59120 61544
rect 800 58688 59200 61264
rect 800 58408 59120 58688
rect 800 58144 59200 58408
rect 880 57864 59200 58144
rect 800 55968 59200 57864
rect 800 55688 59120 55968
rect 800 54336 59200 55688
rect 880 54056 59200 54336
rect 800 53248 59200 54056
rect 800 52968 59120 53248
rect 800 50664 59200 52968
rect 880 50528 59200 50664
rect 880 50384 59120 50528
rect 800 50248 59120 50384
rect 800 47808 59200 50248
rect 800 47528 59120 47808
rect 800 46856 59200 47528
rect 880 46576 59200 46856
rect 800 45088 59200 46576
rect 800 44808 59120 45088
rect 800 43184 59200 44808
rect 880 42904 59200 43184
rect 800 42368 59200 42904
rect 800 42088 59120 42368
rect 800 39648 59200 42088
rect 800 39376 59120 39648
rect 880 39368 59120 39376
rect 880 39096 59200 39368
rect 800 36928 59200 39096
rect 800 36648 59120 36928
rect 800 35704 59200 36648
rect 880 35424 59200 35704
rect 800 34208 59200 35424
rect 800 33928 59120 34208
rect 800 31896 59200 33928
rect 880 31616 59200 31896
rect 800 31488 59200 31616
rect 800 31208 59120 31488
rect 800 28768 59200 31208
rect 800 28488 59120 28768
rect 800 28088 59200 28488
rect 880 27808 59200 28088
rect 800 26048 59200 27808
rect 800 25768 59120 26048
rect 800 24416 59200 25768
rect 880 24136 59200 24416
rect 800 23328 59200 24136
rect 800 23048 59120 23328
rect 800 20608 59200 23048
rect 880 20328 59120 20608
rect 800 17888 59200 20328
rect 800 17608 59120 17888
rect 800 16936 59200 17608
rect 880 16656 59200 16936
rect 800 15168 59200 16656
rect 800 14888 59120 15168
rect 800 13128 59200 14888
rect 880 12848 59200 13128
rect 800 12448 59200 12848
rect 800 12168 59120 12448
rect 800 9728 59200 12168
rect 800 9456 59120 9728
rect 880 9448 59120 9456
rect 880 9176 59200 9448
rect 800 7008 59200 9176
rect 800 6728 59120 7008
rect 800 5648 59200 6728
rect 880 5368 59200 5648
rect 800 4288 59200 5368
rect 800 4008 59120 4288
rect 800 1976 59200 4008
rect 880 1696 59200 1976
rect 800 1568 59200 1696
rect 800 1395 59120 1568
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
<< labels >>
rlabel metal2 s 4986 -800 5042 800 8 clock
port 1 nsew signal input
rlabel metal2 s 26146 119200 26202 120800 6 io_QEI_ChA
port 2 nsew signal input
rlabel metal2 s 33690 119200 33746 120800 6 io_QEI_ChB
port 3 nsew signal input
rlabel metal2 s 56138 119200 56194 120800 6 io_clo_test
port 4 nsew signal input
rlabel metal2 s 54942 -800 54998 800 8 io_irq
port 5 nsew signal output
rlabel metal2 s 3698 119200 3754 120800 6 io_pwm_h
port 6 nsew signal output
rlabel metal2 s 11150 119200 11206 120800 6 io_pwm_l
port 7 nsew signal output
rlabel metal2 s 18694 119200 18750 120800 6 io_pwm_test
port 8 nsew signal input
rlabel metal2 s 41142 119200 41198 120800 6 io_sync_in
port 9 nsew signal input
rlabel metal2 s 48686 119200 48742 120800 6 io_sync_out
port 10 nsew signal output
rlabel metal2 s 44914 -800 44970 800 8 io_wb_ack_o
port 11 nsew signal output
rlabel metal3 s 59200 1368 60800 1488 6 io_wb_adr_i[0]
port 12 nsew signal input
rlabel metal3 s 59200 28568 60800 28688 6 io_wb_adr_i[10]
port 13 nsew signal input
rlabel metal3 s 59200 31288 60800 31408 6 io_wb_adr_i[11]
port 14 nsew signal input
rlabel metal3 s 59200 4088 60800 4208 6 io_wb_adr_i[1]
port 15 nsew signal input
rlabel metal3 s 59200 6808 60800 6928 6 io_wb_adr_i[2]
port 16 nsew signal input
rlabel metal3 s 59200 9528 60800 9648 6 io_wb_adr_i[3]
port 17 nsew signal input
rlabel metal3 s 59200 12248 60800 12368 6 io_wb_adr_i[4]
port 18 nsew signal input
rlabel metal3 s 59200 14968 60800 15088 6 io_wb_adr_i[5]
port 19 nsew signal input
rlabel metal3 s 59200 17688 60800 17808 6 io_wb_adr_i[6]
port 20 nsew signal input
rlabel metal3 s 59200 20408 60800 20528 6 io_wb_adr_i[7]
port 21 nsew signal input
rlabel metal3 s 59200 23128 60800 23248 6 io_wb_adr_i[8]
port 22 nsew signal input
rlabel metal3 s 59200 25848 60800 25968 6 io_wb_adr_i[9]
port 23 nsew signal input
rlabel metal2 s 34978 -800 35034 800 8 io_wb_cs_i
port 24 nsew signal input
rlabel metal3 s 59200 34008 60800 34128 6 io_wb_dat_i[0]
port 25 nsew signal input
rlabel metal3 s 59200 61344 60800 61464 6 io_wb_dat_i[10]
port 26 nsew signal input
rlabel metal3 s 59200 64064 60800 64184 6 io_wb_dat_i[11]
port 27 nsew signal input
rlabel metal3 s 59200 66784 60800 66904 6 io_wb_dat_i[12]
port 28 nsew signal input
rlabel metal3 s 59200 69504 60800 69624 6 io_wb_dat_i[13]
port 29 nsew signal input
rlabel metal3 s 59200 72224 60800 72344 6 io_wb_dat_i[14]
port 30 nsew signal input
rlabel metal3 s 59200 74944 60800 75064 6 io_wb_dat_i[15]
port 31 nsew signal input
rlabel metal3 s 59200 77664 60800 77784 6 io_wb_dat_i[16]
port 32 nsew signal input
rlabel metal3 s 59200 80384 60800 80504 6 io_wb_dat_i[17]
port 33 nsew signal input
rlabel metal3 s 59200 83104 60800 83224 6 io_wb_dat_i[18]
port 34 nsew signal input
rlabel metal3 s 59200 85824 60800 85944 6 io_wb_dat_i[19]
port 35 nsew signal input
rlabel metal3 s 59200 36728 60800 36848 6 io_wb_dat_i[1]
port 36 nsew signal input
rlabel metal3 s 59200 88544 60800 88664 6 io_wb_dat_i[20]
port 37 nsew signal input
rlabel metal3 s 59200 91264 60800 91384 6 io_wb_dat_i[21]
port 38 nsew signal input
rlabel metal3 s 59200 93984 60800 94104 6 io_wb_dat_i[22]
port 39 nsew signal input
rlabel metal3 s 59200 96704 60800 96824 6 io_wb_dat_i[23]
port 40 nsew signal input
rlabel metal3 s 59200 99424 60800 99544 6 io_wb_dat_i[24]
port 41 nsew signal input
rlabel metal3 s 59200 102144 60800 102264 6 io_wb_dat_i[25]
port 42 nsew signal input
rlabel metal3 s 59200 104864 60800 104984 6 io_wb_dat_i[26]
port 43 nsew signal input
rlabel metal3 s 59200 107584 60800 107704 6 io_wb_dat_i[27]
port 44 nsew signal input
rlabel metal3 s 59200 110304 60800 110424 6 io_wb_dat_i[28]
port 45 nsew signal input
rlabel metal3 s 59200 113024 60800 113144 6 io_wb_dat_i[29]
port 46 nsew signal input
rlabel metal3 s 59200 39448 60800 39568 6 io_wb_dat_i[2]
port 47 nsew signal input
rlabel metal3 s 59200 115744 60800 115864 6 io_wb_dat_i[30]
port 48 nsew signal input
rlabel metal3 s 59200 118464 60800 118584 6 io_wb_dat_i[31]
port 49 nsew signal input
rlabel metal3 s 59200 42168 60800 42288 6 io_wb_dat_i[3]
port 50 nsew signal input
rlabel metal3 s 59200 44888 60800 45008 6 io_wb_dat_i[4]
port 51 nsew signal input
rlabel metal3 s 59200 47608 60800 47728 6 io_wb_dat_i[5]
port 52 nsew signal input
rlabel metal3 s 59200 50328 60800 50448 6 io_wb_dat_i[6]
port 53 nsew signal input
rlabel metal3 s 59200 53048 60800 53168 6 io_wb_dat_i[7]
port 54 nsew signal input
rlabel metal3 s 59200 55768 60800 55888 6 io_wb_dat_i[8]
port 55 nsew signal input
rlabel metal3 s 59200 58488 60800 58608 6 io_wb_dat_i[9]
port 56 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 io_wb_dat_o[0]
port 57 nsew signal output
rlabel metal3 s -800 39176 800 39296 4 io_wb_dat_o[10]
port 58 nsew signal output
rlabel metal3 s -800 42984 800 43104 4 io_wb_dat_o[11]
port 59 nsew signal output
rlabel metal3 s -800 46656 800 46776 4 io_wb_dat_o[12]
port 60 nsew signal output
rlabel metal3 s -800 50464 800 50584 4 io_wb_dat_o[13]
port 61 nsew signal output
rlabel metal3 s -800 54136 800 54256 4 io_wb_dat_o[14]
port 62 nsew signal output
rlabel metal3 s -800 57944 800 58064 4 io_wb_dat_o[15]
port 63 nsew signal output
rlabel metal3 s -800 61752 800 61872 4 io_wb_dat_o[16]
port 64 nsew signal output
rlabel metal3 s -800 65424 800 65544 4 io_wb_dat_o[17]
port 65 nsew signal output
rlabel metal3 s -800 69232 800 69352 4 io_wb_dat_o[18]
port 66 nsew signal output
rlabel metal3 s -800 72904 800 73024 4 io_wb_dat_o[19]
port 67 nsew signal output
rlabel metal3 s -800 5448 800 5568 4 io_wb_dat_o[1]
port 68 nsew signal output
rlabel metal3 s -800 76712 800 76832 4 io_wb_dat_o[20]
port 69 nsew signal output
rlabel metal3 s -800 80384 800 80504 4 io_wb_dat_o[21]
port 70 nsew signal output
rlabel metal3 s -800 84192 800 84312 4 io_wb_dat_o[22]
port 71 nsew signal output
rlabel metal3 s -800 87864 800 87984 4 io_wb_dat_o[23]
port 72 nsew signal output
rlabel metal3 s -800 91672 800 91792 4 io_wb_dat_o[24]
port 73 nsew signal output
rlabel metal3 s -800 95480 800 95600 4 io_wb_dat_o[25]
port 74 nsew signal output
rlabel metal3 s -800 99152 800 99272 4 io_wb_dat_o[26]
port 75 nsew signal output
rlabel metal3 s -800 102960 800 103080 4 io_wb_dat_o[27]
port 76 nsew signal output
rlabel metal3 s -800 106632 800 106752 4 io_wb_dat_o[28]
port 77 nsew signal output
rlabel metal3 s -800 110440 800 110560 4 io_wb_dat_o[29]
port 78 nsew signal output
rlabel metal3 s -800 9256 800 9376 4 io_wb_dat_o[2]
port 79 nsew signal output
rlabel metal3 s -800 114112 800 114232 4 io_wb_dat_o[30]
port 80 nsew signal output
rlabel metal3 s -800 117920 800 118040 4 io_wb_dat_o[31]
port 81 nsew signal output
rlabel metal3 s -800 12928 800 13048 4 io_wb_dat_o[3]
port 82 nsew signal output
rlabel metal3 s -800 16736 800 16856 4 io_wb_dat_o[4]
port 83 nsew signal output
rlabel metal3 s -800 20408 800 20528 4 io_wb_dat_o[5]
port 84 nsew signal output
rlabel metal3 s -800 24216 800 24336 4 io_wb_dat_o[6]
port 85 nsew signal output
rlabel metal3 s -800 27888 800 28008 4 io_wb_dat_o[7]
port 86 nsew signal output
rlabel metal3 s -800 31696 800 31816 4 io_wb_dat_o[8]
port 87 nsew signal output
rlabel metal3 s -800 35504 800 35624 4 io_wb_dat_o[9]
port 88 nsew signal output
rlabel metal2 s 24950 -800 25006 800 8 io_wb_we_i
port 89 nsew signal input
rlabel metal2 s 14922 -800 14978 800 8 reset
port 90 nsew signal input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 91 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 94 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/motor_top/runs/motor_top/results/magic/motor_top.gds
string GDS_END 16570526
string GDS_START 892868
<< end >>

