* NGSPICE file created from motor_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt motor_top clock io_QEI_ChA io_QEI_ChB io_clo_test io_irq io_pwm_h io_pwm_l
+ io_pwm_test io_sync_in io_sync_out io_wb_ack_o io_wb_adr_i[0] io_wb_adr_i[10] io_wb_adr_i[11]
+ io_wb_adr_i[1] io_wb_adr_i[2] io_wb_adr_i[3] io_wb_adr_i[4] io_wb_adr_i[5] io_wb_adr_i[6]
+ io_wb_adr_i[7] io_wb_adr_i[8] io_wb_adr_i[9] io_wb_cs_i io_wb_dat_i[0] io_wb_dat_i[10]
+ io_wb_dat_i[11] io_wb_dat_i[12] io_wb_dat_i[13] io_wb_dat_i[14] io_wb_dat_i[15]
+ io_wb_dat_i[16] io_wb_dat_i[17] io_wb_dat_i[18] io_wb_dat_i[19] io_wb_dat_i[1] io_wb_dat_i[20]
+ io_wb_dat_i[21] io_wb_dat_i[22] io_wb_dat_i[23] io_wb_dat_i[24] io_wb_dat_i[25]
+ io_wb_dat_i[26] io_wb_dat_i[27] io_wb_dat_i[28] io_wb_dat_i[29] io_wb_dat_i[2] io_wb_dat_i[30]
+ io_wb_dat_i[31] io_wb_dat_i[3] io_wb_dat_i[4] io_wb_dat_i[5] io_wb_dat_i[6] io_wb_dat_i[7]
+ io_wb_dat_i[8] io_wb_dat_i[9] io_wb_dat_o[0] io_wb_dat_o[10] io_wb_dat_o[11] io_wb_dat_o[12]
+ io_wb_dat_o[13] io_wb_dat_o[14] io_wb_dat_o[15] io_wb_dat_o[16] io_wb_dat_o[17]
+ io_wb_dat_o[18] io_wb_dat_o[19] io_wb_dat_o[1] io_wb_dat_o[20] io_wb_dat_o[21] io_wb_dat_o[22]
+ io_wb_dat_o[23] io_wb_dat_o[24] io_wb_dat_o[25] io_wb_dat_o[26] io_wb_dat_o[27]
+ io_wb_dat_o[28] io_wb_dat_o[29] io_wb_dat_o[2] io_wb_dat_o[30] io_wb_dat_o[31] io_wb_dat_o[3]
+ io_wb_dat_o[4] io_wb_dat_o[5] io_wb_dat_o[6] io_wb_dat_o[7] io_wb_dat_o[8] io_wb_dat_o[9]
+ io_wb_we_i reset vccd1 vssd1
XFILLER_100_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05903_ _05911_/A vssd1 vssd1 vccd1 vccd1 _05903_/X sky130_fd_sc_hd__clkbuf_2
X_09671_ _10152_/Q _10168_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06883_ _06911_/A _07031_/B _07100_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _06885_/A
+ sky130_fd_sc_hd__o22a_1
X_08622_ _08623_/A _09940_/X vssd1 vssd1 vccd1 vccd1 _10042_/D sky130_fd_sc_hd__or2_1
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05834_ _10022_/S vssd1 vssd1 vccd1 vccd1 _05834_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08553_ _08464_/X _08552_/X _08464_/X _08552_/X vssd1 vssd1 vccd1 vccd1 _08554_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_05765_ _07421_/A _05759_/X _09631_/X _05761_/X _05764_/X vssd1 vssd1 vccd1 vccd1
+ _10269_/D sky130_fd_sc_hd__o221a_1
X_08484_ _10066_/Q _08484_/B vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__or2_1
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07504_ _07806_/A _07504_/B vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__or2_2
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05696_ _10299_/Q vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__inv_2
X_07435_ _05804_/A _07428_/B _07429_/B vssd1 vssd1 vccd1 vccd1 _07435_/X sky130_fd_sc_hd__a21bo_1
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07366_ _07071_/X _07074_/X _07075_/X _07096_/X _07054_/X vssd1 vssd1 vccd1 vccd1
+ _07366_/X sky130_fd_sc_hd__o221a_1
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ _09105_/A vssd1 vssd1 vccd1 vccd1 _09105_/Y sky130_fd_sc_hd__inv_2
X_06317_ _10238_/Q _08355_/A _06304_/A _06302_/X vssd1 vssd1 vccd1 vccd1 _06317_/X
+ sky130_fd_sc_hd__o22a_1
X_07297_ _07064_/C _07278_/X _07064_/C _07278_/X vssd1 vssd1 vccd1 vccd1 _07297_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06248_ _10182_/Q _08198_/A vssd1 vssd1 vccd1 vccd1 _06249_/B sky130_fd_sc_hd__or2_1
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09036_ _09036_/A _09036_/B vssd1 vssd1 vccd1 vccd1 _09083_/B sky130_fd_sc_hd__nor2_2
XFILLER_184_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06179_ _06181_/A _09664_/X vssd1 vssd1 vccd1 vccd1 _10114_/D sky130_fd_sc_hd__and2_1
XFILLER_2_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _08956_/X _08954_/Y _09986_/S vssd1 vssd1 vccd1 vccd1 _09938_/X sky130_fd_sc_hd__mux2_2
X_09869_ _09868_/X input39/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09869_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10009_ _07984_/Y _08028_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05550_ _05550_/A vssd1 vssd1 vccd1 vccd1 _05550_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05481_ _05481_/A _05481_/B vssd1 vssd1 vccd1 vccd1 _05481_/Y sky130_fd_sc_hd__nor2_1
X_07220_ _07223_/C _07220_/B vssd1 vssd1 vccd1 vccd1 _07220_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater93 _09944_/S vssd1 vssd1 vccd1 vccd1 _09709_/S sky130_fd_sc_hd__buf_8
XFILLER_118_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07151_ _07147_/A _07164_/B _10219_/Q _07152_/B vssd1 vssd1 vccd1 vccd1 _07151_/X
+ sky130_fd_sc_hd__o211a_1
X_06102_ _06102_/A vssd1 vssd1 vccd1 vccd1 _06102_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07082_ _10225_/Q _07082_/B _07093_/A vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__and3_1
X_06033_ _09841_/X _06028_/X _06030_/X _06031_/X _06032_/X vssd1 vssd1 vccd1 vccd1
+ _10197_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07984_ _07984_/A vssd1 vssd1 vccd1 vccd1 _07984_/Y sky130_fd_sc_hd__inv_2
X_09723_ _06792_/Y _10388_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10054_/D sky130_fd_sc_hd__mux2_1
X_06935_ _07023_/C _07021_/B vssd1 vssd1 vccd1 vccd1 _06935_/X sky130_fd_sc_hd__or2_2
X_09654_ _10120_/Q input50/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06866_ _06866_/A vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08605_ _08289_/A _08499_/X _08604_/X vssd1 vssd1 vccd1 vccd1 _08605_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05817_ _07415_/A _10253_/Q _05811_/Y _05816_/X vssd1 vssd1 vccd1 vccd1 _05817_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06797_ _06818_/A vssd1 vssd1 vccd1 vccd1 _06802_/A sky130_fd_sc_hd__clkbuf_2
X_09585_ _08419_/Y _08418_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _10056_/Q _08474_/B _08475_/B vssd1 vssd1 vccd1 vccd1 _08574_/B sky130_fd_sc_hd__a21bo_1
X_05748_ _05786_/A _05741_/X _09641_/X _05743_/X _05747_/X vssd1 vssd1 vccd1 vccd1
+ _10279_/D sky130_fd_sc_hd__o221a_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _08467_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__nand2_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05679_ _05679_/A vssd1 vssd1 vccd1 vccd1 _05679_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08398_ _09499_/X _08414_/B vssd1 vssd1 vccd1 vccd1 _08398_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07418_ _10270_/Q _07418_/B vssd1 vssd1 vccd1 vccd1 _07427_/B sky130_fd_sc_hd__or2_1
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ _05964_/X _06912_/B _07108_/A _06868_/Y _07348_/X vssd1 vssd1 vccd1 vccd1
+ _07349_/X sky130_fd_sc_hd__a41o_1
X_10360_ _10426_/CLK _10360_/D vssd1 vssd1 vccd1 vccd1 _10360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09019_ _09018_/A _09018_/B _09063_/A vssd1 vssd1 vccd1 vccd1 _09019_/X sky130_fd_sc_hd__a21bo_1
X_10291_ _10420_/CLK _10291_/D vssd1 vssd1 vccd1 vccd1 _10291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06720_ _06635_/Y _06719_/Y _08734_/A vssd1 vssd1 vccd1 vccd1 _06802_/B sky130_fd_sc_hd__o21a_1
XFILLER_110_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ _08457_/A vssd1 vssd1 vccd1 vccd1 _08624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05602_ _05649_/A _05649_/B vssd1 vssd1 vccd1 vccd1 _05648_/A sky130_fd_sc_hd__nand2_1
X_06582_ _06563_/X _06566_/X _06580_/X _06571_/X _06581_/X vssd1 vssd1 vccd1 vccd1
+ _06583_/B sky130_fd_sc_hd__o311a_1
X_09370_ _09368_/X _09369_/X _09368_/X _09369_/X vssd1 vssd1 vccd1 vccd1 _09370_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
X_08321_ _08321_/A _09997_/S _10000_/S vssd1 vssd1 vccd1 vccd1 _08322_/C sky130_fd_sc_hd__or3_1
X_05533_ _05533_/A vssd1 vssd1 vccd1 vccd1 _05534_/B sky130_fd_sc_hd__clkbuf_1
X_08252_ _10194_/Q vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__inv_2
XFILLER_177_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05464_ _10315_/Q _05372_/X _05457_/Y _05409_/X vssd1 vssd1 vccd1 vccd1 _10315_/D
+ sky130_fd_sc_hd__o22ai_1
X_07203_ _07129_/X _07202_/Y _07129_/X _07202_/Y vssd1 vssd1 vccd1 vccd1 _07204_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _08183_/A vssd1 vssd1 vccd1 vccd1 _08184_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_118_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05395_ _05395_/A _05406_/A vssd1 vssd1 vccd1 vccd1 _05404_/A sky130_fd_sc_hd__or2_1
XFILLER_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07134_ _07134_/A vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__inv_2
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07065_ _07068_/C _07065_/B vssd1 vssd1 vccd1 vccd1 _07065_/Y sky130_fd_sc_hd__nand2_1
X_06016_ _10202_/Q vssd1 vssd1 vccd1 vccd1 _06268_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_4 _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07967_ _07963_/X _07964_/X _07963_/X _07964_/X vssd1 vssd1 vccd1 vccd1 _07971_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09706_ _06584_/Y input39/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09706_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06918_ _06903_/A _06913_/Y _06910_/X _06914_/X vssd1 vssd1 vccd1 vccd1 _06925_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07898_ _07878_/X _07897_/Y _07878_/X _07897_/Y vssd1 vssd1 vccd1 vccd1 _07898_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09637_ _06346_/Y _06347_/Y _10175_/Q vssd1 vssd1 vccd1 vccd1 _09637_/X sky130_fd_sc_hd__mux2_1
X_06849_ _06835_/A _06835_/B _06836_/B vssd1 vssd1 vccd1 vccd1 _06849_/X sky130_fd_sc_hd__a21bo_1
XFILLER_43_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ _08391_/Y _09567_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _10061_/Q _08479_/B _08480_/B vssd1 vssd1 vccd1 vccd1 _08519_/X sky130_fd_sc_hd__a21bo_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _09498_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09499_/X sky130_fd_sc_hd__mux2_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ _10414_/CLK _10412_/D vssd1 vssd1 vccd1 vccd1 _10412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _10343_/CLK _10343_/D vssd1 vssd1 vccd1 vccd1 _10343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10274_ _10274_/CLK _10274_/D vssd1 vssd1 vccd1 vccd1 _10274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05180_ _05678_/A vssd1 vssd1 vccd1 vccd1 _05646_/A sky130_fd_sc_hd__buf_2
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _10295_/Q _07458_/Y _08843_/X _08869_/X vssd1 vssd1 vccd1 vccd1 _08870_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07821_ _07824_/C _07821_/B vssd1 vssd1 vccd1 vccd1 _07821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07752_ _07737_/X _07750_/Y _07751_/X vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__a21oi_2
X_06703_ _08717_/A vssd1 vssd1 vccd1 vccd1 _06703_/Y sky130_fd_sc_hd__inv_2
X_07683_ _07671_/A _07671_/B _07671_/X vssd1 vssd1 vccd1 vccd1 _07684_/B sky130_fd_sc_hd__a21bo_1
X_06634_ _10365_/Q vssd1 vssd1 vccd1 vccd1 _06634_/Y sky130_fd_sc_hd__inv_2
X_09422_ _09171_/X _09421_/X _09171_/X _09421_/X vssd1 vssd1 vccd1 vccd1 _09424_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09353_ _09470_/A _09452_/B _09408_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09356_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08304_ _08304_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__or2_1
X_06565_ _10104_/Q vssd1 vssd1 vccd1 vccd1 _08439_/A sky130_fd_sc_hd__inv_2
XFILLER_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09284_ _08377_/A _09282_/A _09283_/A vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__o21ai_1
X_06496_ _06496_/A vssd1 vssd1 vccd1 vccd1 _06496_/X sky130_fd_sc_hd__buf_1
XFILLER_100_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05516_ _06887_/A _07234_/B _07660_/A _07814_/A vssd1 vssd1 vccd1 vccd1 _05516_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_193_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _08166_/X _08230_/Y _06257_/B vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__o21ai_1
X_05447_ _05447_/A vssd1 vssd1 vccd1 vccd1 _10320_/D sky130_fd_sc_hd__inv_2
XFILLER_193_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08166_ _08578_/A vssd1 vssd1 vccd1 vccd1 _08166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05378_ _10324_/Q vssd1 vssd1 vccd1 vccd1 _05391_/A sky130_fd_sc_hd__inv_2
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07117_ _07117_/A vssd1 vssd1 vccd1 vccd1 _07118_/C sky130_fd_sc_hd__inv_2
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08097_ _06657_/Y _08657_/A _08763_/A _08093_/X _08096_/X vssd1 vssd1 vccd1 vccd1
+ _08098_/D sky130_fd_sc_hd__o221a_1
XFILLER_133_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07048_ _07050_/B vssd1 vssd1 vccd1 vccd1 _07048_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08999_ _09948_/X vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10326_ _10328_/CLK _10326_/D vssd1 vssd1 vccd1 vccd1 _10326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10257_ _10274_/CLK _10257_/D vssd1 vssd1 vccd1 vccd1 _10257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10188_ _10426_/CLK _10188_/D vssd1 vssd1 vccd1 vccd1 _10188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06350_ _10243_/Q vssd1 vssd1 vccd1 vccd1 _06351_/A sky130_fd_sc_hd__inv_2
XFILLER_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05301_ _05301_/A _05347_/A vssd1 vssd1 vccd1 vccd1 _05343_/A sky130_fd_sc_hd__or2_1
X_06281_ _10236_/Q vssd1 vssd1 vccd1 vccd1 _06281_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05232_ _10370_/Q _05230_/X input34/X _05231_/X _05227_/X vssd1 vssd1 vccd1 vccd1
+ _10370_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_19_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10426_/CLK sky130_fd_sc_hd__clkbuf_16
X_08020_ _08020_/A _08020_/B vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__or2_1
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05163_ _05179_/A _05163_/B vssd1 vssd1 vccd1 vccd1 _10400_/D sky130_fd_sc_hd__nor2_1
XFILLER_155_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05094_ _05094_/A vssd1 vssd1 vccd1 vccd1 _05094_/X sky130_fd_sc_hd__clkbuf_2
X_09971_ _09970_/X _06961_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08922_ _08920_/A _08920_/B _08942_/A vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08853_ _10287_/Q _07434_/X _10287_/Q _07434_/X vssd1 vssd1 vccd1 vccd1 _08853_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08784_ _08625_/A _08625_/B _08625_/Y vssd1 vssd1 vccd1 vccd1 _08784_/X sky130_fd_sc_hd__a21o_1
X_05996_ _06069_/A vssd1 vssd1 vccd1 vccd1 _06067_/A sky130_fd_sc_hd__inv_2
XFILLER_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07804_ _05966_/X _07800_/X _07802_/X _07803_/Y vssd1 vssd1 vccd1 vccd1 _07804_/X
+ sky130_fd_sc_hd__a31o_1
X_07735_ _07630_/X _07646_/X _07630_/X _07646_/X vssd1 vssd1 vccd1 vccd1 _07737_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ _09474_/B vssd1 vssd1 vccd1 vccd1 _09405_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07667_/B _07677_/A vssd1 vssd1 vccd1 vccd1 _07672_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06617_ _06606_/X _06607_/Y _06614_/X _06615_/X _06616_/X vssd1 vssd1 vccd1 vccd1
+ _06617_/X sky130_fd_sc_hd__o2111a_1
X_07597_ _07597_/A _09920_/X _07597_/C vssd1 vssd1 vccd1 vccd1 _07597_/X sky130_fd_sc_hd__or3_1
XFILLER_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06548_ _06560_/B _06547_/X _06560_/B _06547_/X vssd1 vssd1 vccd1 vccd1 _06548_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09336_ _09336_/A _09336_/B vssd1 vssd1 vccd1 vccd1 _09457_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09267_ _09268_/A _09268_/B vssd1 vssd1 vccd1 vccd1 _09267_/X sky130_fd_sc_hd__and2_1
XFILLER_138_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08093_/X _08213_/Y _06253_/B vssd1 vssd1 vccd1 vccd1 _08218_/Y sky130_fd_sc_hd__o21ai_1
X_06479_ _06482_/B _06478_/Y _06482_/B _06478_/Y vssd1 vssd1 vccd1 vccd1 _06479_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_193_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ _09259_/B vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__buf_2
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08149_ _10196_/Q vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__inv_2
XFILLER_146_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _10450_/CLK _10111_/D vssd1 vssd1 vccd1 vccd1 _10111_/Q sky130_fd_sc_hd__dfxtp_1
X_10042_ _10450_/CLK _10042_/D vssd1 vssd1 vccd1 vccd1 _10042_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _10420_/CLK _10309_/D vssd1 vssd1 vccd1 vccd1 _10309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05850_ _10261_/Q _05780_/X _05842_/X _06837_/A _05845_/X vssd1 vssd1 vccd1 vccd1
+ _10261_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07520_ _07499_/X _07500_/X _07499_/X _07500_/X vssd1 vssd1 vccd1 vccd1 _07521_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_05781_ _10281_/Q vssd1 vssd1 vccd1 vccd1 _07854_/A sky130_fd_sc_hd__inv_2
X_07451_ _07837_/A vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__buf_1
XFILLER_194_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06402_ _06399_/X _06401_/X _06399_/X _06401_/X vssd1 vssd1 vccd1 vccd1 _06402_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_07382_ _07176_/A _07176_/B _07177_/B vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__a21bo_1
X_09121_ _09229_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__inv_2
X_06333_ _10240_/Q _08370_/A _06322_/A _06324_/Y vssd1 vssd1 vccd1 vccd1 _06333_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06264_ _08504_/A _08267_/A vssd1 vssd1 vccd1 vccd1 _06265_/B sky130_fd_sc_hd__or2_1
XFILLER_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _09050_/X _09094_/A _09050_/X _09094_/A vssd1 vssd1 vccd1 vccd1 _09053_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06195_ _09705_/X _06187_/X _10106_/Q _06190_/X vssd1 vssd1 vccd1 vccd1 _10106_/D
+ sky130_fd_sc_hd__a22o_1
X_05215_ _05263_/A vssd1 vssd1 vccd1 vccd1 _05215_/X sky130_fd_sc_hd__clkbuf_2
X_08003_ _08003_/A vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__inv_2
XFILLER_190_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05146_ _10435_/Q vssd1 vssd1 vccd1 vccd1 _05146_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09954_ _06616_/B _08273_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__mux2_1
X_05077_ _10425_/Q _05072_/X input24/X _05073_/X _05070_/X vssd1 vssd1 vccd1 vccd1
+ _10425_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08905_ _08904_/A _08904_/B _08926_/A vssd1 vssd1 vccd1 vccd1 _08905_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09885_ _06823_/X _05883_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__mux2_2
X_08836_ _06272_/A _08708_/X _06271_/A _08710_/X _08835_/X vssd1 vssd1 vccd1 vccd1
+ _08836_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08767_ _08762_/A _08762_/B _08763_/B vssd1 vssd1 vccd1 vccd1 _08767_/X sky130_fd_sc_hd__a21bo_1
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05979_ _07885_/A _05970_/X input45/X _05971_/X _05978_/X vssd1 vssd1 vccd1 vccd1
+ _10214_/D sky130_fd_sc_hd__o221a_1
X_08698_ _08693_/X _08697_/X _08695_/B vssd1 vssd1 vccd1 vccd1 _08698_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_198_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07718_ _07569_/X _07648_/Y _07652_/A vssd1 vssd1 vccd1 vccd1 _07718_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_198_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07649_ _07569_/X _07648_/Y _07569_/X _07648_/Y vssd1 vssd1 vccd1 vccd1 _07650_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ _09319_/A _09319_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__and2_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput75 _09594_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput64 _09584_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput53 _10209_/Q vssd1 vssd1 vccd1 vccd1 io_irq sky130_fd_sc_hd__clkbuf_2
Xoutput86 _10030_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[6] sky130_fd_sc_hd__clkbuf_2
X_10025_ _10044_/Q _09539_/X _08338_/Y _09541_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10025_/X sky130_fd_sc_hd__mux4_2
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05000_ input9/X input6/X input10/X vssd1 vssd1 vccd1 vccd1 _06183_/A sky130_fd_sc_hd__or3_4
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06951_ _06943_/X _06947_/X _06943_/X _06947_/X vssd1 vssd1 vccd1 vccd1 _06951_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ _10151_/Q _10167_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__mux2_1
X_05902_ _05910_/A vssd1 vssd1 vccd1 vccd1 _05902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _10043_/D _10077_/Q vssd1 vssd1 vccd1 vccd1 _08621_/X sky130_fd_sc_hd__and2_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06882_ _09891_/X vssd1 vssd1 vccd1 vccd1 _07031_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05833_ _05830_/Y _05832_/X _05830_/Y _05832_/X vssd1 vssd1 vccd1 vccd1 _10022_/S
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08552_ _08625_/A _10047_/Q _08459_/Y vssd1 vssd1 vccd1 vccd1 _08552_/X sky130_fd_sc_hd__a21o_1
X_05764_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05764_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08483_ _10065_/Q _08511_/A vssd1 vssd1 vccd1 vccd1 _08484_/B sky130_fd_sc_hd__or2_1
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07503_ _07777_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _07506_/A sky130_fd_sc_hd__or2_1
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05695_ _05695_/A _08899_/C vssd1 vssd1 vccd1 vccd1 _05695_/X sky130_fd_sc_hd__and2_1
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07434_/X sky130_fd_sc_hd__buf_2
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07365_ _07317_/X _07318_/X _07316_/X _07319_/X vssd1 vssd1 vccd1 vccd1 _07365_/Y
+ sky130_fd_sc_hd__o22ai_2
X_09104_ _09104_/A vssd1 vssd1 vccd1 vccd1 _09201_/C sky130_fd_sc_hd__inv_2
X_06316_ _06313_/Y _06315_/A _06313_/A _06315_/Y vssd1 vssd1 vccd1 vccd1 _06316_/X
+ sky130_fd_sc_hd__o22a_1
X_07296_ _07296_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _07296_/Y sky130_fd_sc_hd__nand2_2
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06247_ _10181_/Q _06247_/B vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__or2_1
X_09035_ _09034_/A _09034_/B _09083_/A vssd1 vssd1 vccd1 vccd1 _09036_/B sky130_fd_sc_hd__a21o_1
XFILLER_190_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06178_ _06181_/A _09665_/X vssd1 vssd1 vccd1 vccd1 _10115_/D sky130_fd_sc_hd__and2_1
X_05129_ _05202_/A vssd1 vssd1 vccd1 vccd1 _05129_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09937_ _10044_/Q input30/X _09940_/S vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09868_ _09867_/X _08300_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09868_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08819_ _08819_/A _08819_/B _08819_/C _08780_/X vssd1 vssd1 vccd1 vccd1 _08820_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_133_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09799_ _10358_/Q _09798_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09799_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _08035_/X _07389_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10008_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05480_ _10013_/X vssd1 vssd1 vccd1 vccd1 _05481_/B sky130_fd_sc_hd__inv_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater94 _09554_/S vssd1 vssd1 vccd1 vccd1 _09582_/S sky130_fd_sc_hd__buf_4
X_07150_ _07150_/A _09885_/X vssd1 vssd1 vccd1 vccd1 _07155_/C sky130_fd_sc_hd__nor2_2
XFILLER_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06101_ _06101_/A vssd1 vssd1 vccd1 vccd1 _06101_/X sky130_fd_sc_hd__clkbuf_2
X_07081_ _07234_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__or2_1
XFILLER_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06032_ _06032_/A vssd1 vssd1 vccd1 vccd1 _06032_/X sky130_fd_sc_hd__buf_1
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _06791_/Y _10387_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10053_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07983_ _07983_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__nand2_1
X_06934_ _10220_/Q _06929_/Y _05964_/X _06930_/Y _06933_/X vssd1 vssd1 vccd1 vccd1
+ _06937_/A sky130_fd_sc_hd__a41o_1
X_09653_ _10119_/Q input49/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09653_/X sky130_fd_sc_hd__mux2_1
X_06865_ _07063_/A vssd1 vssd1 vccd1 vccd1 _06866_/A sky130_fd_sc_hd__clkbuf_2
X_08604_ _08289_/A _08499_/X _08285_/A _08500_/X _08603_/X vssd1 vssd1 vccd1 vccd1
+ _08604_/X sky130_fd_sc_hd__o221a_1
X_09584_ _08416_/X _09583_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09584_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05816_ _07421_/A _10252_/Q _05812_/Y _05815_/Y vssd1 vssd1 vccd1 vccd1 _05816_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06796_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__clkbuf_2
X_08535_ _08804_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08594_/C sky130_fd_sc_hd__nor2_1
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05747_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _08457_/A _08456_/X _08457_/Y _08465_/X vssd1 vssd1 vccd1 vccd1 _08467_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05678_ _05678_/A vssd1 vssd1 vccd1 vccd1 _08618_/A sky130_fd_sc_hd__clkbuf_2
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__buf_1
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07417_ _10269_/Q _07417_/B vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__or2_1
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07348_ _07023_/C _06960_/B _06961_/A _06949_/D vssd1 vssd1 vccd1 vccd1 _07348_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07279_ _07276_/X _07277_/X _07064_/C _07278_/X vssd1 vssd1 vccd1 vccd1 _07279_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__or2_1
X_10290_ _10420_/CLK _10290_/D vssd1 vssd1 vccd1 vccd1 _10290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06650_ _10450_/Q vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__inv_2
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05601_ _09947_/X _05556_/X _05654_/A vssd1 vssd1 vccd1 vccd1 _05649_/B sky130_fd_sc_hd__o21ai_1
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06581_ _08442_/A _06437_/A _08444_/A _06436_/A vssd1 vssd1 vccd1 vccd1 _06581_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08320_ _08413_/B vssd1 vssd1 vccd1 vccd1 _09748_/S sky130_fd_sc_hd__clkbuf_2
X_05532_ _10009_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _05533_/A sky130_fd_sc_hd__and2_1
X_08251_ _08125_/X _08249_/B _08240_/X _08250_/Y vssd1 vssd1 vccd1 vccd1 _08251_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_177_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05463_ _05456_/Y _05409_/X _05372_/X _05462_/X vssd1 vssd1 vccd1 vccd1 _10316_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07202_ _07202_/A _07202_/B vssd1 vssd1 vccd1 vccd1 _07202_/Y sky130_fd_sc_hd__nor2_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08182_ _08182_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08183_/A sky130_fd_sc_hd__or2_1
XFILLER_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05394_ _05394_/A _05412_/A vssd1 vssd1 vccd1 vccd1 _05406_/A sky130_fd_sc_hd__or2_1
XFILLER_145_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ _07133_/A _07139_/A vssd1 vssd1 vccd1 vccd1 _07133_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07064_ _07219_/A _07126_/B _07064_/C vssd1 vssd1 vccd1 vccd1 _07065_/B sky130_fd_sc_hd__and3_1
X_06015_ _06028_/A vssd1 vssd1 vccd1 vccd1 _06015_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_5 _07777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _07960_/X _07965_/X _07960_/X _07965_/X vssd1 vssd1 vccd1 vccd1 _07966_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09705_ _06577_/X input38/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__mux2_1
X_06917_ _06917_/A vssd1 vssd1 vccd1 vccd1 _06919_/A sky130_fd_sc_hd__inv_2
XFILLER_114_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09636_ _06334_/X _06336_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07897_ _07897_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _07897_/Y sky130_fd_sc_hd__nor2_1
X_06848_ _06836_/A _06836_/B _06837_/B vssd1 vssd1 vccd1 vccd1 _06848_/X sky130_fd_sc_hd__a21bo_1
XFILLER_203_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06779_ _10403_/Q _06811_/B _06778_/Y vssd1 vssd1 vccd1 vccd1 _06779_/X sky130_fd_sc_hd__a21bo_1
XFILLER_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09567_ _08392_/Y _10121_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__mux2_1
X_08518_ _10062_/Q _08480_/B _08481_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__a21bo_1
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09498_ _09497_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09498_/X sky130_fd_sc_hd__mux2_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _09980_/X _08449_/B vssd1 vssd1 vccd1 vccd1 _08449_/Y sky130_fd_sc_hd__nor2_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10414_/CLK _10411_/D vssd1 vssd1 vccd1 vccd1 _10411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ _10343_/CLK _10342_/D vssd1 vssd1 vccd1 vccd1 _10342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10273_ _10298_/CLK _10273_/D vssd1 vssd1 vccd1 vccd1 _10273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07820_ _07820_/A _07885_/B _07820_/C vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__and3_1
X_07751_ _07493_/C _07732_/X _07493_/C _07732_/X vssd1 vssd1 vccd1 vccd1 _07751_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06702_ _10373_/Q _08715_/A _06700_/Y vssd1 vssd1 vccd1 vccd1 _06813_/B sky130_fd_sc_hd__a21oi_2
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07682_ _07770_/A _07662_/B _07662_/X vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__a21bo_1
X_06633_ _06633_/A vssd1 vssd1 vccd1 vccd1 _06633_/Y sky130_fd_sc_hd__inv_2
X_09421_ _09416_/X _09420_/X _09416_/X _09420_/X vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06564_ _06563_/A _06563_/B _06563_/X vssd1 vssd1 vccd1 vccd1 _06564_/Y sky130_fd_sc_hd__a21boi_1
X_09352_ _09341_/X _09351_/X _09341_/X _09351_/X vssd1 vssd1 vccd1 vccd1 _09352_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08303_ _08303_/A vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__buf_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05515_ _07819_/A vssd1 vssd1 vccd1 vccd1 _07814_/A sky130_fd_sc_hd__clkbuf_2
X_09283_ _09283_/A vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__inv_2
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06495_ _06495_/A _06495_/B _06495_/C vssd1 vssd1 vccd1 vccd1 _06498_/A sky130_fd_sc_hd__or3_4
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08234_ _08107_/X _08232_/B _08184_/A _08233_/Y vssd1 vssd1 vccd1 vccd1 _08234_/Y
+ sky130_fd_sc_hd__a211oi_4
X_05446_ _05441_/B _05439_/X _05445_/Y _05387_/A _05424_/A vssd1 vssd1 vccd1 vccd1
+ _05447_/A sky130_fd_sc_hd__o32a_1
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08165_ _10190_/Q vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__inv_2
X_05377_ _10325_/Q vssd1 vssd1 vccd1 vccd1 _05392_/A sky130_fd_sc_hd__inv_2
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07116_ _07125_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07117_/A sky130_fd_sc_hd__or2_2
XFILLER_173_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _06626_/Y _10205_/Q _08625_/B _08554_/A vssd1 vssd1 vccd1 vccd1 _08096_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_118_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07047_ _07311_/A _07228_/A _07213_/A _07047_/D vssd1 vssd1 vccd1 vccd1 _07050_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_102_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08998_ _08998_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _09074_/C sky130_fd_sc_hd__or2_2
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ _07850_/A _07850_/B _07881_/B vssd1 vssd1 vccd1 vccd1 _07949_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _09618_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09619_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10325_ _10328_/CLK _10325_/D vssd1 vssd1 vccd1 vccd1 _10325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10274_/CLK _10256_/D vssd1 vssd1 vccd1 vccd1 _10256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10421_/CLK _10187_/D vssd1 vssd1 vccd1 vccd1 _10187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05300_ _05300_/A _05351_/A vssd1 vssd1 vccd1 vccd1 _05347_/A sky130_fd_sc_hd__or2_1
X_06280_ _10129_/Q vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__inv_2
X_05231_ _05240_/A vssd1 vssd1 vccd1 vccd1 _05231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05162_ _05153_/X _06616_/C _05160_/Y _05161_/X vssd1 vssd1 vccd1 vccd1 _05163_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09970_ _09969_/X _09468_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__mux2_1
X_05093_ input46/X vssd1 vssd1 vccd1 vccd1 _05093_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08921_ _08921_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__inv_2
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ _10288_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _08852_/Y sky130_fd_sc_hd__nor2_1
X_07803_ _05966_/X _07800_/X _07802_/X vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__a21oi_1
X_08783_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__and2_1
X_05995_ _10043_/D _09781_/S vssd1 vssd1 vccd1 vccd1 _06069_/A sky130_fd_sc_hd__or2_2
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07734_ _07729_/X _07733_/X _07729_/X _07733_/X vssd1 vssd1 vccd1 vccd1 _07734_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07665_ _07663_/X _07664_/X _07663_/X _07664_/X vssd1 vssd1 vccd1 vccd1 _07671_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06616_ _06616_/A _06616_/B _06616_/C _06616_/D vssd1 vssd1 vccd1 vccd1 _06616_/X
+ sky130_fd_sc_hd__and4_1
X_09404_ _09396_/X _09403_/X _09396_/X _09403_/X vssd1 vssd1 vccd1 vccd1 _09404_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07596_ _07596_/A _07596_/B vssd1 vssd1 vccd1 vccd1 _07596_/X sky130_fd_sc_hd__or2_1
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06547_ _10099_/Q _06466_/X _06538_/A _06543_/A vssd1 vssd1 vccd1 vccd1 _06547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _08870_/X _09334_/X _08870_/X _09334_/X vssd1 vssd1 vccd1 vccd1 _09336_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _09188_/X _09196_/X _09197_/X _09207_/X vssd1 vssd1 vccd1 vccd1 _09268_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06478_ _08385_/A _06438_/X _06482_/A vssd1 vssd1 vccd1 vccd1 _06478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08217_ _08081_/X _08215_/B _08184_/A _08216_/Y vssd1 vssd1 vccd1 vccd1 _08217_/Y
+ sky130_fd_sc_hd__a211oi_4
X_05429_ _05422_/B _05416_/X _05428_/Y _05391_/A _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05430_/A sky130_fd_sc_hd__o32a_1
X_09197_ _09188_/X _09196_/X _09188_/X _09196_/X vssd1 vssd1 vccd1 vccd1 _09197_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08148_ _08241_/A vssd1 vssd1 vccd1 vccd1 _08533_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08079_ _08600_/A vssd1 vssd1 vccd1 vccd1 _08079_/X sky130_fd_sc_hd__buf_2
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _10207_/CLK _10110_/D vssd1 vssd1 vccd1 vccd1 _10110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10041_ _10450_/CLK _10041_/D vssd1 vssd1 vccd1 vccd1 _10041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _10420_/CLK _10308_/D vssd1 vssd1 vccd1 vccd1 _10308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10239_ _10447_/CLK _10239_/D vssd1 vssd1 vccd1 vccd1 _10239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05780_ _05871_/A vssd1 vssd1 vccd1 vccd1 _05780_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_207_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07450_ _07603_/A vssd1 vssd1 vccd1 vccd1 _07837_/A sky130_fd_sc_hd__buf_1
X_06401_ _06384_/X _06391_/A _06400_/X vssd1 vssd1 vccd1 vccd1 _06401_/X sky130_fd_sc_hd__o21ba_1
XFILLER_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07381_ _07177_/A _07177_/B _07178_/B vssd1 vssd1 vccd1 vccd1 _07398_/A sky130_fd_sc_hd__a21bo_1
X_09120_ _09918_/X vssd1 vssd1 vccd1 vccd1 _09229_/B sky130_fd_sc_hd__clkbuf_2
X_06332_ _06332_/A vssd1 vssd1 vccd1 vccd1 _06332_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _09097_/A _09010_/B _08979_/A _09009_/X _09010_/X vssd1 vssd1 vccd1 vccd1
+ _09094_/A sky130_fd_sc_hd__o32a_1
X_06263_ _06263_/A _06263_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__or2_1
X_08002_ _08002_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__inv_2
X_06194_ _09706_/X _06187_/X _10107_/Q _06190_/X vssd1 vssd1 vccd1 vccd1 _10107_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05214_ _05239_/A vssd1 vssd1 vccd1 vccd1 _05263_/A sky130_fd_sc_hd__clkbuf_4
X_05145_ _10403_/Q vssd1 vssd1 vccd1 vccd1 _06615_/D sky130_fd_sc_hd__inv_2
XFILLER_143_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _09952_/X _06632_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09953_/X sky130_fd_sc_hd__mux2_1
X_05076_ _10426_/Q _05072_/X input25/X _05073_/X _05070_/X vssd1 vssd1 vccd1 vccd1
+ _10426_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__nand2_1
X_09884_ _06822_/X _06412_/Y _10022_/S vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__mux2_2
X_08835_ _10205_/Q _08710_/X _06270_/A _08712_/X _08834_/X vssd1 vssd1 vccd1 vccd1
+ _08835_/X sky130_fd_sc_hd__o221a_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08766_ _08766_/A vssd1 vssd1 vccd1 vccd1 _08766_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05978_ _06111_/A vssd1 vssd1 vccd1 vccd1 _05978_/X sky130_fd_sc_hd__buf_2
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07717_ _07713_/X _07714_/X _07713_/X _07714_/X vssd1 vssd1 vccd1 vccd1 _07717_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08697_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__or2_1
XFILLER_82_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07648_ _07648_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _07648_/Y sky130_fd_sc_hd__nor2_2
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07579_ _07579_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _07579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _09313_/X _09317_/X _09313_/X _09317_/X vssd1 vssd1 vccd1 vccd1 _09321_/A
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09249_ _09451_/A _09462_/B _09073_/A _09248_/X vssd1 vssd1 vccd1 vccd1 _09249_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_5_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput54 _08620_/X vssd1 vssd1 vccd1 vccd1 io_pwm_h sky130_fd_sc_hd__clkbuf_2
Xoutput76 _09595_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput65 _09585_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput87 _10031_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_130_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10024_ _10443_/Q _09535_/X _08323_/X _09537_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10024_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_18_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10312_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ _06950_/A _06949_/X vssd1 vssd1 vccd1 vccd1 _06950_/X sky130_fd_sc_hd__or2b_1
X_05901_ _10247_/Q _05896_/X input23/X _05897_/X _05900_/X vssd1 vssd1 vccd1 vccd1
+ _10247_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06881_ _06880_/A _06880_/B _06880_/Y vssd1 vssd1 vccd1 vccd1 _06881_/X sky130_fd_sc_hd__a21o_1
X_08620_ _10043_/D _10078_/Q vssd1 vssd1 vccd1 vccd1 _08620_/X sky130_fd_sc_hd__and2_1
XFILLER_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05832_ _05831_/Y _10265_/Q _05831_/Y _10265_/Q vssd1 vssd1 vccd1 vccd1 _05832_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08551_ _08551_/A vssd1 vssd1 vccd1 vccd1 _08551_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05763_ _08855_/B _05759_/X _09632_/X _05761_/X _05756_/X vssd1 vssd1 vccd1 vccd1
+ _10270_/D sky130_fd_sc_hd__o221a_1
X_08482_ _10064_/Q _08482_/B vssd1 vssd1 vccd1 vccd1 _08511_/A sky130_fd_sc_hd__or2_1
X_05694_ _05694_/A vssd1 vssd1 vccd1 vccd1 _05694_/Y sky130_fd_sc_hd__inv_2
X_07502_ _07766_/A vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__buf_6
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07433_ _05800_/A _07429_/B _07430_/B vssd1 vssd1 vccd1 vccd1 _07433_/X sky130_fd_sc_hd__a21bo_1
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _09088_/X _09102_/X _09088_/X _09102_/X vssd1 vssd1 vccd1 vccd1 _09105_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07364_ _07320_/X _07325_/X _07326_/X _07363_/X vssd1 vssd1 vccd1 vccd1 _07364_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06315_ _06315_/A vssd1 vssd1 vccd1 vccd1 _06315_/Y sky130_fd_sc_hd__inv_2
X_07295_ _07285_/X _07286_/Y _07287_/X _07294_/X vssd1 vssd1 vccd1 vccd1 _07296_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_163_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06246_ _08137_/A _06246_/B vssd1 vssd1 vccd1 vccd1 _06247_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09034_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06177_ _06181_/A _09666_/X vssd1 vssd1 vccd1 vccd1 _10116_/D sky130_fd_sc_hd__and2_1
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05128_ _05133_/A _05128_/B vssd1 vssd1 vccd1 vccd1 _10407_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05059_ _10437_/Q _05055_/X input37/X _05057_/X _05053_/X vssd1 vssd1 vccd1 vccd1
+ _10437_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _07434_/X _07436_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _09936_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09867_ _10375_/Q _09866_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09867_/X sky130_fd_sc_hd__mux2_1
X_08818_ _08818_/A vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__inv_2
XFILLER_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _08223_/X _10358_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08749_ _08745_/A _08745_/B _06638_/Y _08748_/Y vssd1 vssd1 vccd1 vccd1 _08751_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ _05534_/A _05534_/B _10007_/S vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater95 _09849_/S vssd1 vssd1 vccd1 vccd1 _09881_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06100_ _10339_/Q _06093_/X _10167_/Q _06094_/X _06099_/X vssd1 vssd1 vccd1 vccd1
+ _10167_/D sky130_fd_sc_hd__a221o_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ _07067_/X _07068_/X _07067_/X _07068_/X vssd1 vssd1 vccd1 vccd1 _07080_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_06031_ _06031_/A vssd1 vssd1 vccd1 vccd1 _06031_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_133_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07982_ _07982_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _07983_/B sky130_fd_sc_hd__nand2_1
X_09721_ _06790_/X _10386_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10052_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06933_ _06962_/A _07021_/B _07023_/C _09896_/X vssd1 vssd1 vccd1 vccd1 _06933_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09652_ _10118_/Q input48/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09652_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06864_ _07218_/A vssd1 vssd1 vccd1 vccd1 _07063_/A sky130_fd_sc_hd__buf_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ _08285_/A _08500_/X _08281_/A _08599_/B _08602_/Y vssd1 vssd1 vccd1 vccd1
+ _08603_/X sky130_fd_sc_hd__a221o_1
X_06795_ _06795_/A _06795_/B vssd1 vssd1 vccd1 vccd1 _06795_/Y sky130_fd_sc_hd__nor2_1
X_09583_ _08414_/Y _09582_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09583_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05815_ _05815_/A vssd1 vssd1 vccd1 vccd1 _05815_/Y sky130_fd_sc_hd__inv_2
X_08534_ _10058_/Q _08476_/B _08477_/B vssd1 vssd1 vccd1 vccd1 _08535_/B sky130_fd_sc_hd__a21bo_1
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05746_ _06119_/A vssd1 vssd1 vccd1 vccd1 _05866_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ _10449_/Q _08657_/B _08459_/Y _08464_/X vssd1 vssd1 vccd1 vccd1 _08465_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05677_ _05677_/A _05677_/B vssd1 vssd1 vccd1 vccd1 _10303_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08396_ _08396_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08396_/X sky130_fd_sc_hd__or2_1
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ _10268_/Q _07594_/C vssd1 vssd1 vccd1 vccd1 _07417_/B sky130_fd_sc_hd__or2_2
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07347_ _07343_/X _07344_/X _07343_/X _07344_/X vssd1 vssd1 vccd1 vccd1 _07347_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09017_ _09017_/A vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__inv_2
X_07278_ _07276_/X _07277_/X _07276_/X _07277_/X vssd1 vssd1 vccd1 vccd1 _07278_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06229_ _09681_/X _06224_/X _10082_/Q _06225_/X vssd1 vssd1 vccd1 vccd1 _10082_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09919_ _07423_/Y _07426_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _09919_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05600_ _05655_/A _05655_/B vssd1 vssd1 vccd1 vccd1 _05654_/A sky130_fd_sc_hd__or2_1
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06580_ _06580_/A _06570_/X vssd1 vssd1 vccd1 vccd1 _06580_/X sky130_fd_sc_hd__or2b_1
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05531_ _10009_/X _09905_/X vssd1 vssd1 vccd1 vccd1 _05534_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08250_ _08255_/B vssd1 vssd1 vccd1 vccd1 _08250_/Y sky130_fd_sc_hd__inv_2
X_05462_ _10316_/Q _10315_/Q _05456_/Y _05457_/Y vssd1 vssd1 vccd1 vccd1 _05462_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__nor2_2
X_07201_ _07142_/X _07184_/X _07185_/X _07200_/X vssd1 vssd1 vccd1 vccd1 _07204_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07132_ _07117_/A _07127_/Y _07124_/X _07128_/X vssd1 vssd1 vccd1 vccd1 _07139_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05393_ _05393_/A _05417_/A vssd1 vssd1 vccd1 vccd1 _05412_/A sky130_fd_sc_hd__or2_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07063_ _07063_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07064_/C sky130_fd_sc_hd__or2_2
X_06014_ _09865_/X _05998_/X _06269_/A _06002_/X _06005_/X vssd1 vssd1 vccd1 vccd1
+ _10203_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_6 _08618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07965_ _07919_/X _07962_/X _07963_/X _07964_/X vssd1 vssd1 vccd1 vccd1 _07965_/X
+ sky130_fd_sc_hd__o22a_1
X_09704_ _06573_/X input37/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06916_ _06899_/X _06900_/X _06899_/X _06900_/X vssd1 vssd1 vccd1 vccd1 _06917_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09635_ _06325_/X _06328_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09635_/X sky130_fd_sc_hd__mux2_1
X_07896_ _07874_/X _07895_/Y _07874_/X _07895_/Y vssd1 vssd1 vccd1 vccd1 _07896_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06847_ _07100_/A vssd1 vssd1 vccd1 vccd1 _07118_/A sky130_fd_sc_hd__clkbuf_2
X_06778_ _10403_/Q _06811_/B _06777_/Y vssd1 vssd1 vccd1 vccd1 _06778_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09566_ _08388_/Y _10120_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09566_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08517_ _10195_/Q _08513_/B _10194_/Q _08516_/Y vssd1 vssd1 vccd1 vccd1 _08517_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _09496_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09497_/X sky130_fd_sc_hd__mux2_1
X_05729_ _10287_/Q _05728_/X _10271_/Q _05719_/X _05724_/X vssd1 vssd1 vccd1 vccd1
+ _10287_/D sky130_fd_sc_hd__o221a_1
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08448_ _08448_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08448_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10410_ _10442_/CLK _10410_/D vssd1 vssd1 vccd1 vccd1 _10410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08379_ _09621_/X _08391_/B vssd1 vssd1 vccd1 vccd1 _08379_/Y sky130_fd_sc_hd__nor2_1
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10341_ _10343_/CLK _10341_/D vssd1 vssd1 vccd1 vccd1 _10341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ _10298_/CLK _10272_/D vssd1 vssd1 vccd1 vccd1 _10272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07750_/Y sky130_fd_sc_hd__nand2_2
X_06701_ _06699_/Y _06700_/Y _08711_/A vssd1 vssd1 vccd1 vccd1 _06814_/B sky130_fd_sc_hd__o21a_1
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07681_ _07675_/X _07680_/X _07675_/X _07680_/X vssd1 vssd1 vccd1 vccd1 _07681_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06632_ _10368_/Q vssd1 vssd1 vccd1 vccd1 _06632_/Y sky130_fd_sc_hd__inv_2
X_09420_ _05922_/X _09417_/Y _09423_/B _09464_/A vssd1 vssd1 vccd1 vccd1 _09420_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06563_ _06563_/A _06563_/B vssd1 vssd1 vccd1 vccd1 _06563_/X sky130_fd_sc_hd__or2_2
X_09351_ _09392_/A _09304_/B _09350_/Y _09304_/Y _09350_/A vssd1 vssd1 vccd1 vccd1
+ _09351_/X sky130_fd_sc_hd__o32a_2
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08302_ _06271_/A _06271_/B _08301_/Y vssd1 vssd1 vccd1 vccd1 _08302_/X sky130_fd_sc_hd__a21o_1
X_09282_ _09282_/A vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__inv_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05514_ _07591_/A vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__buf_1
X_08233_ _08236_/B vssd1 vssd1 vccd1 vccd1 _08233_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06494_ _06494_/A vssd1 vssd1 vccd1 vccd1 _06516_/A sky130_fd_sc_hd__inv_2
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05445_ _10320_/Q _05445_/B vssd1 vssd1 vccd1 vccd1 _05445_/Y sky130_fd_sc_hd__nor2_1
X_08164_ _06653_/Y _10179_/Q _06636_/Y _10192_/Q _08163_/X vssd1 vssd1 vccd1 vccd1
+ _08175_/C sky130_fd_sc_hd__o221a_1
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05376_ _10326_/Q vssd1 vssd1 vccd1 vccd1 _05393_/A sky130_fd_sc_hd__inv_2
X_08095_ _08788_/A vssd1 vssd1 vccd1 vccd1 _08554_/A sky130_fd_sc_hd__clkbuf_2
X_07115_ _07101_/X _07102_/X _07113_/X _07114_/X vssd1 vssd1 vccd1 vccd1 _07115_/X
+ sky130_fd_sc_hd__o22a_1
X_07046_ _05943_/X _07082_/B _07050_/A _07008_/A vssd1 vssd1 vccd1 vccd1 _07046_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08997_ _08994_/X _08996_/X _08994_/X _08996_/X vssd1 vssd1 vccd1 vccd1 _08997_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _07944_/X _07945_/X _07944_/X _07945_/X vssd1 vssd1 vccd1 vccd1 _07948_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07879_ _07879_/A _07878_/X vssd1 vssd1 vccd1 vccd1 _07879_/X sky130_fd_sc_hd__or2b_1
XFILLER_204_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09618_ _08378_/X _06330_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09618_/X sky130_fd_sc_hd__mux2_1
X_09549_ _10383_/Q _10180_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__mux2_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ _10329_/CLK _10324_/D vssd1 vssd1 vccd1 vccd1 _10324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10255_ _10274_/CLK _10255_/D vssd1 vssd1 vccd1 vccd1 _10255_/Q sky130_fd_sc_hd__dfxtp_1
X_10186_ _10421_/CLK _10186_/D vssd1 vssd1 vccd1 vccd1 _10186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05230_ _05239_/A vssd1 vssd1 vccd1 vccd1 _05230_/X sky130_fd_sc_hd__clkbuf_2
X_05161_ _05161_/A vssd1 vssd1 vccd1 vccd1 _05161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05092_ _05091_/X _05082_/X _10417_/Q _05083_/X _05086_/X vssd1 vssd1 vccd1 vccd1
+ _10417_/D sky130_fd_sc_hd__a221o_1
XFILLER_6_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__or2_1
XFILLER_130_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08851_ _10289_/Q _05801_/X _10289_/Q _05801_/X vssd1 vssd1 vccd1 vccd1 _08851_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07802_ _07802_/A _07864_/A vssd1 vssd1 vccd1 vccd1 _07802_/X sky130_fd_sc_hd__or2_1
X_08782_ _08782_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _08818_/A sky130_fd_sc_hd__or2_1
X_05994_ _05116_/X _05990_/Y _05990_/A _05992_/X _05993_/X vssd1 vssd1 vccd1 vccd1
+ _10208_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07733_ _07730_/X _07731_/X _07493_/C _07732_/X vssd1 vssd1 vccd1 vccd1 _07733_/X
+ sky130_fd_sc_hd__o22a_1
X_07664_ _07672_/A _07677_/A vssd1 vssd1 vccd1 vccd1 _07664_/X sky130_fd_sc_hd__or2_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06615_ _06615_/A _06615_/B _06615_/C _06615_/D vssd1 vssd1 vccd1 vccd1 _06615_/X
+ sky130_fd_sc_hd__and4_1
X_09403_ _09402_/A _09402_/B _09402_/Y vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__a21o_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _07597_/C _07593_/X _08000_/A vssd1 vssd1 vccd1 vccd1 _07596_/B sky130_fd_sc_hd__a21oi_1
XFILLER_178_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06546_ _10100_/Q _06464_/A _08430_/A _06540_/A vssd1 vssd1 vccd1 vccd1 _06560_/B
+ sky130_fd_sc_hd__a22o_1
X_09334_ _08842_/A _05704_/X _08842_/Y vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09265_ _09250_/X _09264_/X _09250_/X _09264_/X vssd1 vssd1 vccd1 vccd1 _09268_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06477_ _10088_/Q _06461_/A _08388_/A _06487_/A vssd1 vssd1 vccd1 vccd1 _06482_/B
+ sky130_fd_sc_hd__a22o_1
X_08216_ _08220_/B vssd1 vssd1 vccd1 vccd1 _08216_/Y sky130_fd_sc_hd__inv_2
X_09196_ _09191_/X _09195_/Y _09191_/X _09195_/Y vssd1 vssd1 vccd1 vccd1 _09196_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05428_ _10324_/Q _05428_/B vssd1 vssd1 vccd1 vccd1 _05428_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08147_ _10191_/Q vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__inv_2
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05359_ _05298_/A _05362_/A _05298_/C vssd1 vssd1 vccd1 vccd1 _05359_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08078_ _10199_/Q vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__inv_2
XFILLER_134_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07029_ _05943_/X _06868_/Y _07028_/X vssd1 vssd1 vccd1 vccd1 _07029_/Y sky130_fd_sc_hd__a21oi_1
X_10040_ _10244_/CLK _10040_/D vssd1 vssd1 vccd1 vccd1 _10040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10307_ _10420_/CLK _10307_/D vssd1 vssd1 vccd1 vccd1 _10307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10238_ _10447_/CLK _10238_/D vssd1 vssd1 vccd1 vccd1 _10238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ _10343_/CLK _10169_/D vssd1 vssd1 vccd1 vccd1 _10169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06400_ _10247_/Q _08405_/A _06391_/B _06394_/X vssd1 vssd1 vccd1 vccd1 _06400_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07380_ _07293_/A _07293_/B _07293_/X vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__a21bo_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06331_ _06330_/A _10134_/Q _06330_/Y vssd1 vssd1 vccd1 vccd1 _06332_/A sky130_fd_sc_hd__a21oi_2
X_06262_ _06262_/A _08257_/A vssd1 vssd1 vccd1 vccd1 _06263_/B sky130_fd_sc_hd__or2_1
X_09050_ _05931_/X _09168_/B _09048_/X _09049_/Y vssd1 vssd1 vccd1 vccd1 _09050_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05213_ _05240_/A vssd1 vssd1 vccd1 vccd1 _05239_/A sky130_fd_sc_hd__inv_2
X_08001_ _08001_/A vssd1 vssd1 vccd1 vccd1 _08001_/X sky130_fd_sc_hd__clkbuf_1
X_06193_ _09707_/X _06187_/X _10108_/Q _06190_/X vssd1 vssd1 vccd1 vccd1 _10108_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05144_ _05157_/A _05144_/B vssd1 vssd1 vccd1 vccd1 _10404_/D sky130_fd_sc_hd__nor2_1
X_09952_ _06616_/C _08269_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__mux2_1
X_05075_ _10427_/Q _05072_/X input26/X _05073_/X _05070_/X vssd1 vssd1 vccd1 vccd1
+ _10427_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08903_ _08903_/A vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__inv_2
X_09883_ _10446_/Q input3/X _10042_/Q vssd1 vssd1 vccd1 vccd1 _09899_/S sky130_fd_sc_hd__mux2_8
X_08834_ _06270_/A _08712_/X _06269_/A _08714_/X _08833_/X vssd1 vssd1 vccd1 vccd1
+ _08834_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08765_ _08765_/A _08766_/A vssd1 vssd1 vccd1 vccd1 _08765_/X sky130_fd_sc_hd__or2_1
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05977_ _10214_/Q vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__clkbuf_2
X_07716_ _07710_/X _07715_/X _07710_/X _07715_/X vssd1 vssd1 vccd1 vccd1 _07716_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08696_ _08681_/X _08685_/X _08705_/C vssd1 vssd1 vccd1 vccd1 _08696_/X sky130_fd_sc_hd__o21ba_1
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07647_ _07582_/X _07629_/X _07630_/X _07646_/X vssd1 vssd1 vccd1 vccd1 _07650_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07578_ _07578_/A _07578_/B vssd1 vssd1 vccd1 vccd1 _07648_/B sky130_fd_sc_hd__nor2_2
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09317_ _09315_/Y _09316_/X _09315_/Y _09316_/X vssd1 vssd1 vccd1 vccd1 _09317_/X
+ sky130_fd_sc_hd__o2bb2a_2
X_06529_ _06539_/C _06529_/B vssd1 vssd1 vccd1 vccd1 _06529_/X sky130_fd_sc_hd__and2_1
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09248_ _09186_/X _09187_/X _09181_/X _09185_/X vssd1 vssd1 vccd1 vccd1 _09248_/X
+ sky130_fd_sc_hd__o211a_1
X_09179_ _09026_/X _09133_/X _09134_/X _09135_/X vssd1 vssd1 vccd1 vccd1 _09181_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput55 _08621_/X vssd1 vssd1 vccd1 vccd1 io_pwm_l sky130_fd_sc_hd__clkbuf_2
XFILLER_122_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput66 _09586_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[17] sky130_fd_sc_hd__clkbuf_2
Xoutput77 _09596_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput88 _10032_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _08007_/A _08040_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10023_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05900_ _05934_/A vssd1 vssd1 vccd1 vccd1 _05900_/X sky130_fd_sc_hd__clkbuf_2
X_06880_ _06880_/A _06880_/B vssd1 vssd1 vccd1 vccd1 _06880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05831_ _10282_/Q vssd1 vssd1 vccd1 vccd1 _05831_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08550_ _08204_/A _08569_/B _08200_/A _08549_/X vssd1 vssd1 vccd1 vccd1 _08551_/A
+ sky130_fd_sc_hd__o22a_1
X_05762_ _10271_/Q _05759_/X _09633_/X _05761_/X _05756_/X vssd1 vssd1 vccd1 vccd1
+ _10271_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08481_ _10063_/Q _08481_/B vssd1 vssd1 vccd1 vccd1 _08482_/B sky130_fd_sc_hd__or2_2
X_05693_ _08618_/A _05693_/B vssd1 vssd1 vccd1 vccd1 _10300_/D sky130_fd_sc_hd__nor2_1
X_07501_ _07477_/X _07484_/Y _07499_/X _07500_/X vssd1 vssd1 vccd1 vccd1 _07501_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _08850_/B _07430_/B _07431_/Y vssd1 vssd1 vccd1 vccd1 _07432_/X sky130_fd_sc_hd__a21o_1
XFILLER_148_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _09192_/A _09101_/B _09101_/Y vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__a21o_1
X_07363_ _07333_/X _07361_/X _07371_/B vssd1 vssd1 vccd1 vccd1 _07363_/X sky130_fd_sc_hd__o21a_1
X_06314_ _06299_/Y _10131_/Q _06305_/A vssd1 vssd1 vccd1 vccd1 _06315_/A sky130_fd_sc_hd__o21ai_1
X_07294_ _07288_/X _07290_/X _07291_/X _07293_/X vssd1 vssd1 vccd1 vccd1 _07294_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06245_ _10179_/Q _06245_/B vssd1 vssd1 vccd1 vccd1 _06246_/B sky130_fd_sc_hd__nor2_2
X_09033_ _09031_/X _09077_/A _09031_/X _09077_/A vssd1 vssd1 vccd1 vccd1 _09034_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06176_ _06176_/A vssd1 vssd1 vccd1 vccd1 _06181_/A sky130_fd_sc_hd__buf_1
XFILLER_190_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05127_ _05116_/X _06614_/D _05126_/Y _05113_/X vssd1 vssd1 vccd1 vccd1 _05128_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05058_ _10438_/Q _05055_/X input38/X _05057_/X _05053_/X vssd1 vssd1 vccd1 vccd1
+ _10438_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09935_ _05801_/X _07433_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__mux2_2
X_09866_ _08298_/Y _10375_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09866_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08817_ _08817_/A _08817_/B _08797_/X vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__or3b_1
X_09797_ _09796_/X input20/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09797_/X sky130_fd_sc_hd__mux2_1
X_08748_ _08748_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _08748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08679_ _06030_/X _08671_/Y _06026_/X _08668_/Y vssd1 vssd1 vccd1 vccd1 _08679_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10006_ _08029_/X _07386_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10006_/X sky130_fd_sc_hd__mux2_2
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater96 _09821_/S vssd1 vssd1 vccd1 vccd1 _09849_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_200_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06030_ _06263_/A vssd1 vssd1 vccd1 vccd1 _06030_/X sky130_fd_sc_hd__buf_2
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07981_ _07982_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__or2_1
X_09720_ _06789_/X _10385_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10051_/D sky130_fd_sc_hd__mux2_1
X_06932_ _06942_/A vssd1 vssd1 vccd1 vccd1 _07023_/C sky130_fd_sc_hd__clkbuf_2
X_09651_ _10117_/Q input47/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09651_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06863_ _10222_/Q vssd1 vssd1 vccd1 vccd1 _07218_/A sky130_fd_sc_hd__inv_2
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08602_ _08602_/A _08602_/B vssd1 vssd1 vccd1 vccd1 _08602_/Y sky130_fd_sc_hd__nor2_1
X_06794_ _06795_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _08415_/Y _10126_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05814_ _07423_/A _10251_/Q _05505_/Y _05888_/A vssd1 vssd1 vccd1 vccd1 _05815_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08533_ _08533_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__or2_1
XFILLER_82_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05745_ _05704_/X _05741_/X _09642_/X _05743_/X _05737_/X vssd1 vssd1 vccd1 vccd1
+ _10280_/D sky130_fd_sc_hd__o221a_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _05024_/A _08460_/Y _08461_/Y _08463_/Y vssd1 vssd1 vccd1 vccd1 _08464_/X
+ sky130_fd_sc_hd__o22a_1
X_05676_ _05653_/X _05672_/Y _05673_/Y _08063_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05677_/B sky130_fd_sc_hd__o32a_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _09529_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08395_/Y sky130_fd_sc_hd__nor2_2
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07415_ _07415_/A vssd1 vssd1 vccd1 vccd1 _07415_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07346_ _07341_/X _07345_/X _07341_/X _07345_/X vssd1 vssd1 vccd1 vccd1 _07346_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_17_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10433_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09016_ _09014_/X _09015_/X _09014_/X _09015_/X vssd1 vssd1 vccd1 vccd1 _09017_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07277_ _07269_/A _07269_/B _07269_/X vssd1 vssd1 vccd1 vccd1 _07277_/X sky130_fd_sc_hd__a21bo_1
XFILLER_191_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06228_ _09682_/X _06224_/X _10083_/Q _06225_/X vssd1 vssd1 vccd1 vccd1 _10083_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06159_ _09649_/X _06156_/X _10131_/Q _06157_/X _06154_/X vssd1 vssd1 vccd1 vccd1
+ _10131_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _09118_/X _09116_/Y _09994_/S vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__mux2_1
X_09849_ _09848_/X input34/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05530_ _10018_/X _10006_/X _05469_/X _05529_/X vssd1 vssd1 vccd1 vccd1 _05530_/Y
+ sky130_fd_sc_hd__o22ai_4
X_05461_ _05461_/A vssd1 vssd1 vccd1 vccd1 _10317_/D sky130_fd_sc_hd__inv_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08180_ _08180_/A vssd1 vssd1 vccd1 vccd1 _08182_/A sky130_fd_sc_hd__inv_2
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07200_ _07186_/X _07187_/X _07188_/X _07199_/X vssd1 vssd1 vccd1 vccd1 _07200_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05392_ _05392_/A _05421_/A vssd1 vssd1 vccd1 vccd1 _05417_/A sky130_fd_sc_hd__or2_1
X_07131_ _07131_/A vssd1 vssd1 vccd1 vccd1 _07133_/A sky130_fd_sc_hd__inv_2
XFILLER_158_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07062_ _07063_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07068_/C sky130_fd_sc_hd__nor2_1
X_06013_ _10203_/Q vssd1 vssd1 vccd1 vccd1 _06269_/A sky130_fd_sc_hd__buf_1
XFILLER_173_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_7 _05934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07964_ _07919_/X _07962_/X _07919_/X _07962_/X vssd1 vssd1 vccd1 vccd1 _07964_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09703_ _06568_/X input36/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07895_ _07875_/X _07888_/X _07889_/X _07894_/X vssd1 vssd1 vccd1 vccd1 _07895_/Y
+ sky130_fd_sc_hd__o22ai_1
X_06915_ _06910_/X _06914_/X _06910_/X _06914_/X vssd1 vssd1 vccd1 vccd1 _06946_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _06316_/X _06318_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09634_/X sky130_fd_sc_hd__mux2_1
X_06846_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07100_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06777_ _06616_/A _06710_/A _06776_/Y vssd1 vssd1 vccd1 vccd1 _06777_/Y sky130_fd_sc_hd__o21ai_1
X_09565_ _09564_/X _10356_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08516_ _08516_/A vssd1 vssd1 vccd1 vccd1 _08516_/Y sky130_fd_sc_hd__inv_2
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05728_ _05741_/A vssd1 vssd1 vccd1 vccd1 _05728_/X sky130_fd_sc_hd__clkbuf_2
X_09496_ _08396_/X _06370_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _09959_/X _08449_/B vssd1 vssd1 vccd1 vccd1 _08447_/Y sky130_fd_sc_hd__nor2_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05659_ _05561_/X _05598_/X _05561_/X _05598_/X vssd1 vssd1 vccd1 vccd1 _05659_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _08378_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08378_/X sky130_fd_sc_hd__or2_1
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07329_ _06878_/X _06956_/X _06878_/X _06956_/X vssd1 vssd1 vccd1 vccd1 _07329_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10340_ _10343_/CLK _10340_/D vssd1 vssd1 vccd1 vccd1 _10340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _10300_/CLK _10271_/D vssd1 vssd1 vccd1 vccd1 _10271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06700_ _08713_/A vssd1 vssd1 vccd1 vccd1 _06700_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07680_ _07773_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07680_/X sky130_fd_sc_hd__or2_1
XFILLER_25_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06631_ _10369_/Q vssd1 vssd1 vccd1 vccd1 _06631_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06562_ _06542_/A _06560_/X _06542_/B _06561_/X vssd1 vssd1 vccd1 vccd1 _06563_/B
+ sky130_fd_sc_hd__o211a_1
X_09350_ _09350_/A vssd1 vssd1 vccd1 vccd1 _09350_/Y sky130_fd_sc_hd__inv_2
X_08301_ _08301_/A vssd1 vssd1 vccd1 vccd1 _08301_/Y sky130_fd_sc_hd__inv_2
X_09281_ _09280_/A _09280_/B _09336_/A vssd1 vssd1 vccd1 vccd1 _09281_/X sky130_fd_sc_hd__a21o_1
X_05513_ _07588_/A vssd1 vssd1 vccd1 vccd1 _07591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08236_/B sky130_fd_sc_hd__or2_1
X_06493_ _10091_/Q _06461_/A _08403_/A _06496_/A vssd1 vssd1 vccd1 vccd1 _06494_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05444_ _05444_/A vssd1 vssd1 vccd1 vccd1 _05445_/B sky130_fd_sc_hd__inv_2
X_08163_ _10358_/Q _08160_/X _10372_/Q _08162_/X vssd1 vssd1 vccd1 vccd1 _08163_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05375_ _10327_/Q vssd1 vssd1 vccd1 vccd1 _05394_/A sky130_fd_sc_hd__inv_2
X_08094_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__inv_2
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07114_ _07101_/X _07102_/X _07101_/X _07102_/X vssd1 vssd1 vccd1 vccd1 _07114_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07045_ _07013_/X _07016_/X _07013_/X _07016_/X vssd1 vssd1 vccd1 vccd1 _07052_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _08921_/A _08943_/A _08972_/Y _08970_/A _08995_/Y vssd1 vssd1 vccd1 vccd1
+ _08996_/X sky130_fd_sc_hd__o32a_1
XFILLER_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07947_ _07941_/X _07946_/X _07941_/X _07946_/X vssd1 vssd1 vccd1 vccd1 _07947_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07878_ _07878_/A _09924_/X _07878_/C _07878_/D vssd1 vssd1 vccd1 vccd1 _07878_/X
+ sky130_fd_sc_hd__or4_4
X_09617_ _09616_/X _10362_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09617_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06829_ _06829_/A _06829_/B vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__or2_1
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09548_ _08351_/Y _10114_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09548_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09479_ _09436_/X _09437_/X _09438_/X _09439_/X vssd1 vssd1 vccd1 vccd1 _09479_/Y
+ sky130_fd_sc_hd__o22ai_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _10329_/CLK _10323_/D vssd1 vssd1 vccd1 vccd1 _10323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10254_ _10274_/CLK _10254_/D vssd1 vssd1 vccd1 vccd1 _10254_/Q sky130_fd_sc_hd__dfxtp_1
X_10185_ _10421_/CLK _10185_/D vssd1 vssd1 vccd1 vccd1 _10185_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05160_ _10432_/Q vssd1 vssd1 vccd1 vccd1 _05160_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05091_ input47/X vssd1 vssd1 vccd1 vccd1 _05091_/X sky130_fd_sc_hd__buf_4
XFILLER_170_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08850_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07801_ _09914_/X vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__clkbuf_2
X_08781_ _08632_/A _08632_/B _08752_/B vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__o21ai_1
XFILLER_97_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05993_ _06111_/A vssd1 vssd1 vccd1 vccd1 _05993_/X sky130_fd_sc_hd__buf_2
XFILLER_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07732_ _07730_/X _07731_/X _07730_/X _07731_/X vssd1 vssd1 vccd1 vccd1 _07732_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07663_ _07663_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07663_/X sky130_fd_sc_hd__or2_1
XFILLER_198_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06614_ _06614_/A _06614_/B _06614_/C _06614_/D vssd1 vssd1 vccd1 vccd1 _06614_/X
+ sky130_fd_sc_hd__and4_1
X_09402_ _09402_/A _09402_/B vssd1 vssd1 vccd1 vccd1 _09402_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09333_ _09332_/A _09332_/B _09384_/A vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__a21bo_1
X_07594_ _10210_/Q _07612_/A _07594_/C _10211_/Q vssd1 vssd1 vccd1 vccd1 _08000_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06545_ _10100_/Q vssd1 vssd1 vccd1 vccd1 _08430_/A sky130_fd_sc_hd__inv_2
XFILLER_193_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09264_ _09319_/A _09319_/B _09319_/A _09319_/B vssd1 vssd1 vccd1 vccd1 _09264_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06476_ _10088_/Q vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__inv_2
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08215_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__or2_1
X_09195_ _09195_/A vssd1 vssd1 vccd1 vccd1 _09195_/Y sky130_fd_sc_hd__inv_2
X_05427_ _05427_/A vssd1 vssd1 vccd1 vccd1 _05428_/B sky130_fd_sc_hd__inv_2
XFILLER_193_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _10348_/Q vssd1 vssd1 vccd1 vccd1 _08146_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05358_ _05358_/A vssd1 vssd1 vccd1 vccd1 _10335_/D sky130_fd_sc_hd__inv_2
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08077_ _08181_/B vssd1 vssd1 vccd1 vccd1 _08077_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05289_ _10338_/Q vssd1 vssd1 vccd1 vccd1 _05302_/A sky130_fd_sc_hd__inv_2
XFILLER_161_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07028_ _07028_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__or2_1
XFILLER_121_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ _08979_/A vssd1 vssd1 vccd1 vccd1 _09010_/C sky130_fd_sc_hd__inv_2
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _10420_/CLK _10306_/D vssd1 vssd1 vccd1 vccd1 _10306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10237_ _10447_/CLK _10237_/D vssd1 vssd1 vccd1 vccd1 _10237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10343_/CLK _10168_/D vssd1 vssd1 vccd1 vccd1 _10168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10099_ _10442_/CLK _10099_/D vssd1 vssd1 vccd1 vccd1 _10099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
X_06330_ _06330_/A _10134_/Q vssd1 vssd1 vccd1 vccd1 _06330_/Y sky130_fd_sc_hd__nor2_1
X_06261_ _08733_/A _06261_/B vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__or2_1
XFILLER_148_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05212_ _05968_/A _08328_/A vssd1 vssd1 vccd1 vccd1 _05240_/A sky130_fd_sc_hd__or2_4
X_08000_ _08000_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__or2_1
X_06192_ _09708_/X _06187_/X _10109_/Q _06190_/X vssd1 vssd1 vccd1 vccd1 _10109_/D
+ sky130_fd_sc_hd__a22o_1
X_05143_ _05129_/X _06615_/C _05142_/Y _05138_/X vssd1 vssd1 vccd1 vccd1 _05144_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09951_ _09950_/X _10366_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__mux2_2
X_05074_ _10428_/Q _05072_/X input27/X _05073_/X _05070_/X vssd1 vssd1 vccd1 vccd1
+ _10428_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08902_ _08936_/C _08901_/B _08923_/A vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__a21bo_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09882_ _10414_/Q _08062_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__mux2_1
X_08833_ _06268_/A _08716_/X _06269_/A _08714_/X _08832_/X vssd1 vssd1 vccd1 vccd1
+ _08833_/X sky130_fd_sc_hd__o221a_1
X_08764_ _08084_/Y _08763_/Y _08753_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__o21ai_2
X_05976_ _07885_/C _05970_/X input46/X _05971_/X _05960_/X vssd1 vssd1 vccd1 vccd1
+ _10215_/D sky130_fd_sc_hd__o221a_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07715_ _07711_/X _07712_/X _07713_/X _07714_/X vssd1 vssd1 vccd1 vccd1 _07715_/X
+ sky130_fd_sc_hd__o22a_1
X_08695_ _08695_/A _08695_/B _08695_/C _08695_/D vssd1 vssd1 vccd1 vccd1 _08705_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07646_ _07631_/X _07632_/X _07633_/X _07645_/X vssd1 vssd1 vccd1 vccd1 _07646_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07578_/B sky130_fd_sc_hd__or2_1
X_09316_ _09354_/C _09462_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__or3_1
X_06528_ _08418_/A _06434_/A _08420_/A _06434_/A vssd1 vssd1 vccd1 vccd1 _06529_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_178_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _09247_/A vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06459_ _08382_/A _06442_/X _10086_/Q _06460_/A vssd1 vssd1 vccd1 vccd1 _06471_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _09171_/X _09177_/X _09171_/A _09177_/X vssd1 vssd1 vccd1 vccd1 _09178_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08129_ _08181_/A vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput56 _09874_/S vssd1 vssd1 vccd1 vccd1 io_sync_out sky130_fd_sc_hd__clkbuf_2
XFILLER_162_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput67 _09587_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput78 _09597_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput89 _10033_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10022_ _08039_/X _07392_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05830_ _05782_/X _05783_/Y _05784_/X _05829_/X vssd1 vssd1 vccd1 vccd1 _05830_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05761_ _05761_/A vssd1 vssd1 vccd1 vccd1 _05761_/X sky130_fd_sc_hd__buf_2
X_07500_ _07477_/X _07484_/Y _07477_/X _07484_/Y vssd1 vssd1 vccd1 vccd1 _07500_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08480_ _10062_/Q _08480_/B vssd1 vssd1 vccd1 vccd1 _08481_/B sky130_fd_sc_hd__or2_1
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05692_ _05771_/A _05689_/Y _05690_/X _08060_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05693_/B sky130_fd_sc_hd__o32a_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07431_ _07438_/B vssd1 vssd1 vccd1 vccd1 _07431_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__or2_1
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09101_ _09192_/A _09101_/B vssd1 vssd1 vccd1 vccd1 _09101_/Y sky130_fd_sc_hd__nor2_1
X_06313_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06313_/Y sky130_fd_sc_hd__inv_2
X_07293_ _07293_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07293_/X sky130_fd_sc_hd__or2_1
XFILLER_191_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06244_ _10178_/Q _08180_/A vssd1 vssd1 vccd1 vccd1 _06245_/B sky130_fd_sc_hd__or2_2
X_09032_ _09029_/A _09128_/A _08959_/A _09000_/X _09001_/X vssd1 vssd1 vccd1 vccd1
+ _09077_/A sky130_fd_sc_hd__o32a_1
X_06175_ _06175_/A _09667_/X vssd1 vssd1 vccd1 vccd1 _10117_/D sky130_fd_sc_hd__and2_1
X_05126_ _10439_/Q vssd1 vssd1 vccd1 vccd1 _05126_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05057_ _05095_/A vssd1 vssd1 vccd1 vccd1 _05057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _08852_/B _07435_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09934_/X sky130_fd_sc_hd__mux2_2
X_09865_ _09864_/X input38/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09865_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08816_ _08772_/A _08772_/B _08772_/Y vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__o21ai_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09796_ _09795_/X _08221_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09796_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08747_ _10191_/Q _08747_/B vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__or2_1
X_05959_ _07165_/A _05947_/A input44/X _05948_/A _05950_/X vssd1 vssd1 vccd1 vccd1
+ _10221_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08678_ _06038_/X _08676_/Y _06035_/X _08524_/Y _08677_/X vssd1 vssd1 vccd1 vccd1
+ _08678_/X sky130_fd_sc_hd__o221a_1
XFILLER_26_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07629_ _07600_/X _07605_/X _07606_/X _07628_/X _07584_/X vssd1 vssd1 vccd1 vccd1
+ _07629_/X sky130_fd_sc_hd__o221a_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10005_ _08051_/X _07398_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__mux2_2
XFILLER_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater97 _09801_/S vssd1 vssd1 vccd1 vccd1 _09821_/S sky130_fd_sc_hd__buf_2
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07980_ _07976_/Y _07979_/Y _07976_/Y _07979_/Y vssd1 vssd1 vccd1 vccd1 _07982_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06931_ _06931_/A vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__clkbuf_2
X_09650_ _10116_/Q input46/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09650_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08601_ _08586_/A _08586_/B _08598_/Y _08599_/Y _08600_/Y vssd1 vssd1 vccd1 vccd1
+ _08602_/B sky130_fd_sc_hd__a311o_1
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
X_06862_ _07234_/A vssd1 vssd1 vccd1 vccd1 _07054_/C sky130_fd_sc_hd__clkbuf_2
X_06793_ _09717_/S _06793_/B vssd1 vssd1 vccd1 vccd1 _06793_/X sky130_fd_sc_hd__and2_1
X_09581_ _08412_/Y _09580_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09581_/X sky130_fd_sc_hd__mux2_1
X_05813_ _07423_/A _10251_/Q _10268_/Q _10251_/Q vssd1 vssd1 vccd1 vccd1 _05888_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_08532_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _08587_/A sky130_fd_sc_hd__or2_1
X_05744_ _10281_/Q _05741_/X _09643_/X _05743_/X _05737_/X vssd1 vssd1 vccd1 vccd1
+ _10281_/D sky130_fd_sc_hd__o221a_1
X_08463_ _08463_/A vssd1 vssd1 vccd1 vccd1 _08463_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05675_ _05750_/A vssd1 vssd1 vccd1 vccd1 _05675_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ _07369_/X _07413_/Y _07369_/X _07413_/Y vssd1 vssd1 vccd1 vccd1 _07414_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08394_ _08453_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__buf_2
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07345_ _07016_/X _07342_/X _07343_/X _07344_/X vssd1 vssd1 vccd1 vccd1 _07345_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_1
X_07276_ _07204_/A _07204_/B _07206_/A vssd1 vssd1 vccd1 vccd1 _07276_/X sky130_fd_sc_hd__a21bo_1
XFILLER_163_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06227_ _09683_/X _06224_/X _10084_/Q _06225_/X vssd1 vssd1 vccd1 vccd1 _10084_/D
+ sky130_fd_sc_hd__a22o_1
X_09015_ _08977_/X _08981_/X _08947_/X _08982_/X vssd1 vssd1 vccd1 vccd1 _09015_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06158_ _09650_/X _06156_/X _10132_/Q _06157_/X _06154_/X vssd1 vssd1 vccd1 vccd1
+ _10132_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05109_ _10442_/Q vssd1 vssd1 vccd1 vccd1 _05109_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06089_ _06102_/A vssd1 vssd1 vccd1 vccd1 _06089_/X sky130_fd_sc_hd__clkbuf_2
X_09917_ _07437_/Y _07443_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09917_/X sky130_fd_sc_hd__mux2_1
X_09848_ _09847_/X _08279_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09779_ _10353_/Q _09778_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05460_ _05452_/B _05439_/X _05459_/X _05458_/Y _05424_/A vssd1 vssd1 vccd1 vccd1
+ _05461_/A sky130_fd_sc_hd__o32a_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05391_ _05391_/A _05427_/A vssd1 vssd1 vccd1 vccd1 _05421_/A sky130_fd_sc_hd__or2_1
XFILLER_201_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _07113_/X _07114_/X _07113_/X _07114_/X vssd1 vssd1 vccd1 vccd1 _07131_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_173_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07061_ _09889_/X vssd1 vssd1 vccd1 vccd1 _07102_/B sky130_fd_sc_hd__clkbuf_2
X_06012_ _09869_/X _05998_/X _06270_/A _06002_/X _06005_/X vssd1 vssd1 vccd1 vccd1
+ _10204_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_8 _10226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _07734_/X _07753_/Y _07734_/X _07753_/Y vssd1 vssd1 vccd1 vccd1 _07963_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09702_ _06564_/Y input35/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07894_ _07894_/A _07894_/B vssd1 vssd1 vccd1 vccd1 _07894_/X sky130_fd_sc_hd__or2_1
X_06914_ _06904_/C _06913_/A _06903_/A _06913_/Y vssd1 vssd1 vccd1 vccd1 _06914_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09633_ _06306_/Y _06307_/Y _10175_/Q vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__mux2_1
X_06845_ _07146_/C vssd1 vssd1 vccd1 vccd1 _07161_/A sky130_fd_sc_hd__clkbuf_2
X_09564_ _10388_/Q _10185_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__mux2_1
X_08515_ _10063_/Q _08481_/B _08482_/B vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__a21bo_1
X_06776_ _10401_/Q _06808_/B _10402_/Q _06810_/B _06775_/X vssd1 vssd1 vccd1 vccd1
+ _06776_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ _09494_/X _10358_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09495_/X sky130_fd_sc_hd__mux2_1
X_05727_ _10288_/Q _05715_/X _05804_/A _05719_/X _05724_/X vssd1 vssd1 vccd1 vccd1
+ _10288_/D sky130_fd_sc_hd__o221a_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08446_ _08446_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08446_/Y sky130_fd_sc_hd__nor2_1
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05658_ _05677_/A _05658_/B vssd1 vssd1 vccd1 vccd1 _10307_/D sky130_fd_sc_hd__nor2_1
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08377_ _08377_/A vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__buf_6
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05589_ _05685_/A _05685_/B vssd1 vssd1 vccd1 vccd1 _05684_/A sky130_fd_sc_hd__nand2_1
X_07328_ _07050_/A _07050_/B _07050_/Y vssd1 vssd1 vccd1 vccd1 _07328_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07259_ _07141_/X _07206_/X _07141_/X _07206_/X vssd1 vssd1 vccd1 vccd1 _07259_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _10298_/CLK _10270_/D vssd1 vssd1 vccd1 vccd1 _10270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10399_ _10399_/CLK _10399_/D vssd1 vssd1 vccd1 vccd1 _10399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06630_ _10371_/Q vssd1 vssd1 vccd1 vccd1 _06630_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10066_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06561_ _08432_/A _06435_/A _08434_/A _06540_/X _06551_/X vssd1 vssd1 vccd1 vccd1
+ _06561_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08300_ _06270_/A _08295_/Y _08264_/X _08304_/B vssd1 vssd1 vccd1 vccd1 _08300_/X
+ sky130_fd_sc_hd__o211a_1
X_06492_ _10091_/Q vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__inv_2
X_09280_ _09280_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__nor2_2
X_05512_ _10210_/Q vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__inv_2
X_08231_ _10189_/Q _06255_/B _08230_/Y vssd1 vssd1 vccd1 vccd1 _08231_/X sky130_fd_sc_hd__a21o_1
X_05443_ _05443_/A vssd1 vssd1 vccd1 vccd1 _10321_/D sky130_fd_sc_hd__inv_2
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08162_ _08285_/A vssd1 vssd1 vccd1 vccd1 _08162_/X sky130_fd_sc_hd__buf_2
XFILLER_158_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05374_ _10328_/Q vssd1 vssd1 vccd1 vccd1 _05395_/A sky130_fd_sc_hd__inv_2
X_08093_ _08220_/A vssd1 vssd1 vccd1 vccd1 _08093_/X sky130_fd_sc_hd__clkbuf_2
X_07113_ _07103_/X _07104_/X _07111_/X _07112_/X vssd1 vssd1 vccd1 vccd1 _07113_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07044_ _07032_/X _07043_/X _07032_/X _07043_/X vssd1 vssd1 vccd1 vccd1 _07044_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08995_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ _07942_/Y _07943_/X _07944_/X _07945_/X vssd1 vssd1 vccd1 vccd1 _07946_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07877_ _07877_/A vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__clkbuf_2
X_09616_ _10394_/Q _10191_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09616_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06828_ _06828_/A _06828_/B vssd1 vssd1 vccd1 vccd1 _06829_/B sky130_fd_sc_hd__or2_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06759_ _10388_/Q _06792_/B _10387_/Q _06791_/B _06758_/X vssd1 vssd1 vccd1 vccd1
+ _06759_/Y sky130_fd_sc_hd__o221ai_2
X_09547_ _09546_/X _10350_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09461_/X _09477_/Y _09461_/X _09477_/Y vssd1 vssd1 vccd1 vccd1 _09478_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08429_ _08452_/B vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _10329_/CLK _10322_/D vssd1 vssd1 vccd1 vccd1 _10322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10253_ _10274_/CLK _10253_/D vssd1 vssd1 vccd1 vccd1 _10253_/Q sky130_fd_sc_hd__dfxtp_1
X_10184_ _10421_/CLK _10184_/D vssd1 vssd1 vccd1 vccd1 _10184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05090_ _05089_/X _05082_/X _10418_/Q _05083_/X _05086_/X vssd1 vssd1 vccd1 vccd1
+ _10418_/D sky130_fd_sc_hd__a221o_1
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08780_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__or2_1
XFILLER_97_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07800_ _07885_/D vssd1 vssd1 vccd1 vccd1 _07800_/X sky130_fd_sc_hd__clkbuf_2
X_05992_ _10043_/Q _09973_/X vssd1 vssd1 vccd1 vccd1 _05992_/X sky130_fd_sc_hd__and2_2
XFILLER_84_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07731_ _07722_/A _07722_/B _07722_/X vssd1 vssd1 vccd1 vccd1 _07731_/X sky130_fd_sc_hd__a21bo_1
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _07770_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07662_/X sky130_fd_sc_hd__or2_2
X_09401_ _09468_/A _09922_/X _09291_/X vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__or3b_1
X_06613_ _06613_/A _06613_/B _06613_/C _06613_/D vssd1 vssd1 vccd1 vccd1 _06613_/Y
+ sky130_fd_sc_hd__nor4_2
X_07593_ _05510_/A _07591_/A _10211_/Q _07612_/A vssd1 vssd1 vccd1 vccd1 _07593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06544_ _06560_/A _06543_/Y _06538_/A _06543_/A vssd1 vssd1 vccd1 vccd1 _06544_/X
+ sky130_fd_sc_hd__o22a_1
X_09332_ _09332_/A _09332_/B vssd1 vssd1 vccd1 vccd1 _09384_/A sky130_fd_sc_hd__or2_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _09262_/A _09262_/B _09320_/A vssd1 vssd1 vccd1 vccd1 _09319_/B sky130_fd_sc_hd__a21oi_1
X_06475_ _06474_/A _06474_/B _06482_/A vssd1 vssd1 vccd1 vccd1 _06475_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _09100_/A _09192_/Y _09150_/Y _09147_/Y _09193_/X vssd1 vssd1 vccd1 vccd1
+ _09195_/A sky130_fd_sc_hd__a32o_1
X_08214_ _10185_/Q _06251_/B _08213_/Y vssd1 vssd1 vccd1 vccd1 _08214_/X sky130_fd_sc_hd__a21o_1
X_05426_ _05426_/A vssd1 vssd1 vccd1 vccd1 _10325_/D sky130_fd_sc_hd__inv_2
X_08145_ _08204_/A vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__clkbuf_2
X_05357_ _05352_/B _05333_/A _05356_/Y _05336_/A _05299_/A vssd1 vssd1 vccd1 vccd1
+ _05358_/A sky130_fd_sc_hd__o32a_1
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _10176_/Q vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__inv_2
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05288_ _10339_/Q vssd1 vssd1 vccd1 vccd1 _05303_/A sky130_fd_sc_hd__inv_2
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ _06965_/X _07026_/Y _06965_/X _07026_/Y vssd1 vssd1 vccd1 vccd1 _07027_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08978_ _08978_/A vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07929_ _07929_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07982_/A sky130_fd_sc_hd__nand2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10305_ _10420_/CLK _10305_/D vssd1 vssd1 vccd1 vccd1 _10305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10236_ _10447_/CLK _10236_/D vssd1 vssd1 vccd1 vccd1 _10236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10167_ _10343_/CLK _10167_/D vssd1 vssd1 vccd1 vccd1 _10167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10098_ _10442_/CLK _10098_/D vssd1 vssd1 vccd1 vccd1 _10098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06260_ _06260_/A _08247_/A vssd1 vssd1 vccd1 vccd1 _06261_/B sky130_fd_sc_hd__or2_1
XFILLER_148_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05211_ _08329_/D _08324_/A _08324_/C vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__or3_4
X_06191_ _09709_/X _06187_/X _10110_/Q _06190_/X vssd1 vssd1 vccd1 vccd1 _10110_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05142_ _10436_/Q vssd1 vssd1 vccd1 vccd1 _05142_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09950_ _10398_/Q _10195_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__mux2_1
X_05073_ _05073_/A vssd1 vssd1 vccd1 vccd1 _05073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08901_ _08936_/C _08901_/B vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__or2_2
X_09881_ _09880_/X input43/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08832_ _06268_/A _08716_/X _06020_/X _08718_/X _08831_/Y vssd1 vssd1 vccd1 vccd1
+ _08832_/X sky130_fd_sc_hd__a221o_1
X_08763_ _08763_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _08763_/Y sky130_fd_sc_hd__nor2_2
X_05975_ _10215_/Q vssd1 vssd1 vccd1 vccd1 _07885_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07714_ _07711_/X _07712_/X _07711_/X _07712_/X vssd1 vssd1 vccd1 vccd1 _07714_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08694_ _08697_/B _08694_/B _08697_/A _08693_/X vssd1 vssd1 vccd1 vccd1 _08695_/D
+ sky130_fd_sc_hd__or4bb_4
XFILLER_93_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07645_ _07637_/X _07641_/X _07642_/X _07644_/X vssd1 vssd1 vccd1 vccd1 _07645_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07576_ _07552_/C _07548_/B _07548_/Y vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__o21ai_1
X_09315_ _09315_/A vssd1 vssd1 vccd1 vccd1 _09315_/Y sky130_fd_sc_hd__inv_2
X_06527_ _06527_/A _06527_/B vssd1 vssd1 vccd1 vccd1 _06539_/C sky130_fd_sc_hd__or2_1
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ _09189_/X _09190_/X _09191_/X _09195_/Y _09245_/X vssd1 vssd1 vccd1 vccd1
+ _09246_/X sky130_fd_sc_hd__o221a_1
X_06458_ _10086_/Q vssd1 vssd1 vccd1 vccd1 _08382_/A sky130_fd_sc_hd__inv_2
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05409_ _05423_/A vssd1 vssd1 vccd1 vccd1 _05409_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _09294_/C _09176_/B _09240_/A vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__a21bo_1
X_06389_ _10247_/Q vssd1 vssd1 vccd1 vccd1 _06390_/A sky130_fd_sc_hd__inv_2
X_08128_ _10177_/Q vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__inv_2
XFILLER_107_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ _08059_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08059_/Y sky130_fd_sc_hd__nor2_1
Xoutput57 _08839_/X vssd1 vssd1 vccd1 vccd1 io_wb_ack_o sky130_fd_sc_hd__clkbuf_2
Xoutput79 _09598_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput68 _09588_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10021_ _08041_/X _07393_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10021_/X sky130_fd_sc_hd__mux2_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10219_ _10300_/CLK _10219_/D vssd1 vssd1 vccd1 vccd1 _10219_/Q sky130_fd_sc_hd__dfxtp_2
X_05760_ _05804_/A _05759_/X _09634_/X _05753_/X _05756_/X vssd1 vssd1 vccd1 vccd1
+ _10272_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05691_ _10300_/Q vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__inv_2
XFILLER_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07430_ _10274_/Q _07430_/B vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__or2_1
XFILLER_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07361_ _07334_/X _07339_/X _07340_/X _07360_/X vssd1 vssd1 vccd1 vccd1 _07361_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09100_ _09100_/A _09193_/A vssd1 vssd1 vccd1 vccd1 _09101_/B sky130_fd_sc_hd__nor2_2
X_06312_ _06312_/A _06312_/B vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__or2_2
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ _05941_/X _09251_/A _09029_/X _09030_/Y vssd1 vssd1 vccd1 vccd1 _09031_/X
+ sky130_fd_sc_hd__a31o_1
X_07292_ _07197_/A _07197_/B _07197_/X vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__a21bo_1
X_06243_ _10177_/Q _10176_/Q vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__or2_1
XFILLER_163_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06174_ _06175_/A _09669_/X vssd1 vssd1 vccd1 vccd1 _10118_/D sky130_fd_sc_hd__and2_1
X_05125_ _10407_/Q vssd1 vssd1 vccd1 vccd1 _06614_/D sky130_fd_sc_hd__inv_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05056_ _05073_/A vssd1 vssd1 vccd1 vccd1 _05095_/A sky130_fd_sc_hd__clkbuf_4
X_09933_ _05797_/Y _07432_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__mux2_1
X_09864_ _09863_/X _08296_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08815_ _08815_/A _08815_/B _08815_/C _08774_/X vssd1 vssd1 vccd1 vccd1 _08820_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09795_ _10357_/Q _09794_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08746_ _08742_/A _08745_/B _06722_/Y _08745_/Y vssd1 vssd1 vccd1 vccd1 _08747_/B
+ sky130_fd_sc_hd__o22a_1
X_05958_ _10221_/Q vssd1 vssd1 vccd1 vccd1 _07165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08677_ _08260_/A _10064_/Q _08253_/X _10063_/Q vssd1 vssd1 vccd1 vccd1 _08677_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05889_ _07686_/A _05505_/B _05888_/Y _05505_/Y _05888_/A vssd1 vssd1 vccd1 vccd1
+ _06819_/B sky130_fd_sc_hd__o32a_1
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07628_ _07622_/A _07640_/A _07621_/Y _07619_/A _07627_/Y vssd1 vssd1 vccd1 vccd1
+ _07628_/X sky130_fd_sc_hd__o32a_1
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07559_ _07555_/X _07558_/X _07555_/X _07558_/X vssd1 vssd1 vccd1 vccd1 _07559_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ _09451_/A _09229_/B _09294_/C vssd1 vssd1 vccd1 vccd1 _09229_/X sky130_fd_sc_hd__or3_4
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10443_/Q input4/X _10042_/Q vssd1 vssd1 vccd1 vccd1 _10043_/D sky130_fd_sc_hd__mux2_4
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater98 _09781_/S vssd1 vssd1 vccd1 vccd1 _09801_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06930_ _09896_/X vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__inv_2
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08600_/Y sky130_fd_sc_hd__nor2_1
X_06861_ _07212_/A vssd1 vssd1 vccd1 vccd1 _07234_/A sky130_fd_sc_hd__clkbuf_2
X_06792_ _06795_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06792_/Y sky130_fd_sc_hd__nor2_1
X_09580_ _08410_/Y _09579_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__mux2_1
X_05812_ _10269_/Q _10252_/Q vssd1 vssd1 vccd1 vccd1 _05812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_208_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08531_ _10059_/Q _08477_/B _08478_/B vssd1 vssd1 vccd1 vccd1 _08578_/B sky130_fd_sc_hd__a21bo_1
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05743_ _05761_/A vssd1 vssd1 vccd1 vccd1 _05743_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08462_ _05024_/A _08460_/Y _06658_/Y _10046_/Q vssd1 vssd1 vccd1 vccd1 _08463_/A
+ sky130_fd_sc_hd__o22a_1
X_05674_ _10303_/Q vssd1 vssd1 vccd1 vccd1 _08063_/A sky130_fd_sc_hd__inv_2
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07413_ _07413_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07413_/Y sky130_fd_sc_hd__nor2_2
XFILLER_195_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08393_ _08445_/B vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__inv_2
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ _07300_/X _07301_/X _07300_/X _07301_/X vssd1 vssd1 vccd1 vccd1 _07344_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07275_ _07272_/X _07273_/X _07272_/X _07273_/X vssd1 vssd1 vccd1 vccd1 _07275_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_163_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06226_ _09684_/X _06224_/X _10085_/Q _06225_/X vssd1 vssd1 vccd1 vccd1 _10085_/D
+ sky130_fd_sc_hd__a22o_1
X_09014_ _09007_/X _09013_/X _09007_/X _09013_/X vssd1 vssd1 vccd1 vccd1 _09014_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06157_ _06157_/A vssd1 vssd1 vccd1 vccd1 _06157_/X sky130_fd_sc_hd__buf_1
XFILLER_208_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05108_ _05202_/A vssd1 vssd1 vccd1 vccd1 _05193_/A sky130_fd_sc_hd__clkbuf_4
X_06088_ _06101_/A vssd1 vssd1 vccd1 vccd1 _06088_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05039_ _10443_/Q _05012_/A _05038_/X _05013_/A _05036_/X vssd1 vssd1 vccd1 vccd1
+ _10443_/D sky130_fd_sc_hd__o221a_1
X_09916_ _07445_/X _07447_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _09916_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09847_ _10370_/Q _09846_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09847_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09778_ _08203_/Y _10353_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09778_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ _08729_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08729_/X sky130_fd_sc_hd__or2_1
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05390_ _05390_/A _05431_/A vssd1 vssd1 vccd1 vccd1 _05427_/A sky130_fd_sc_hd__or2_1
XFILLER_192_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07060_ _07058_/X _07059_/X _07058_/X _07059_/X vssd1 vssd1 vccd1 vccd1 _07067_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06011_ _10204_/Q vssd1 vssd1 vccd1 vccd1 _06270_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _06557_/X input34/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09701_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_9 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07962_ _07854_/D _07885_/B _07820_/A _07800_/X _07961_/X vssd1 vssd1 vccd1 vccd1
+ _07962_/X sky130_fd_sc_hd__a41o_1
XFILLER_114_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07893_ _07792_/X _07891_/X _07867_/X _07892_/X vssd1 vssd1 vccd1 vccd1 _07894_/B
+ sky130_fd_sc_hd__o22a_1
X_06913_ _06913_/A vssd1 vssd1 vccd1 vccd1 _06913_/Y sky130_fd_sc_hd__inv_2
X_09632_ _06296_/X _06298_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09632_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06844_ _10221_/Q vssd1 vssd1 vccd1 vccd1 _07146_/C sky130_fd_sc_hd__inv_2
X_09563_ _08385_/Y _10119_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__mux2_1
X_08514_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08514_/Y sky130_fd_sc_hd__inv_2
X_06775_ _10401_/Q _06808_/B _10400_/Q _06807_/B _06774_/X vssd1 vssd1 vccd1 vccd1
+ _06775_/X sky130_fd_sc_hd__a221o_1
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09494_ _10390_/Q _10187_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05726_ _10272_/Q vssd1 vssd1 vccd1 vccd1 _05804_/A sky130_fd_sc_hd__buf_2
XFILLER_211_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08445_ _09965_/X _08445_/B vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__and2_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05657_ _05653_/X _05654_/Y _05655_/X _08069_/A _05644_/X vssd1 vssd1 vccd1 vccd1
+ _05658_/B sky130_fd_sc_hd__o32a_1
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08376_ _09245_/A vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05588_ _09978_/X _05576_/X _09978_/X _05576_/X vssd1 vssd1 vccd1 vccd1 _05685_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07327_ _07323_/X _07324_/X _07323_/X _07324_/X vssd1 vssd1 vccd1 vccd1 _07362_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07258_ _07229_/X _07248_/X _07229_/X _07248_/X vssd1 vssd1 vccd1 vccd1 _07258_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06209_ _09695_/X _06203_/X _10096_/Q _06204_/X vssd1 vssd1 vccd1 vccd1 _10096_/D
+ sky130_fd_sc_hd__a22o_1
X_07189_ _07189_/A vssd1 vssd1 vccd1 vccd1 _07189_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10398_ _10433_/CLK _10398_/D vssd1 vssd1 vccd1 vccd1 _10398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06560_ _06560_/A _06560_/B _06560_/C _06560_/D vssd1 vssd1 vccd1 vccd1 _06560_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_178_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06491_ _06495_/B _06490_/Y _06495_/B _06490_/Y vssd1 vssd1 vccd1 vccd1 _06491_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05511_ _07667_/A vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__clkbuf_2
X_08230_ _08230_/A vssd1 vssd1 vccd1 vccd1 _08230_/Y sky130_fd_sc_hd__inv_2
X_05442_ _05436_/B _05439_/X _05441_/Y _05388_/A _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05443_/A sky130_fd_sc_hd__o32a_1
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ _10201_/Q vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__inv_2
XFILLER_158_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05373_ _10329_/Q vssd1 vssd1 vccd1 vccd1 _05396_/A sky130_fd_sc_hd__inv_2
XFILLER_173_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _10186_/Q vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__inv_2
X_07112_ _07112_/A _09887_/X _07112_/C vssd1 vssd1 vccd1 vccd1 _07112_/X sky130_fd_sc_hd__or3_1
X_07043_ _07038_/X _07042_/Y _07038_/X _07042_/Y vssd1 vssd1 vccd1 vccd1 _07043_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ _08991_/X _08993_/X _08991_/X _08993_/X vssd1 vssd1 vccd1 vccd1 _08994_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07945_ _07942_/Y _07943_/X _07942_/Y _07943_/X vssd1 vssd1 vccd1 vccd1 _07945_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _09614_/X _06642_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09615_/X sky130_fd_sc_hd__mux2_2
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _07877_/A _09924_/X _07855_/A _07878_/D vssd1 vssd1 vccd1 vccd1 _07879_/A
+ sky130_fd_sc_hd__o22a_1
X_06827_ _06827_/A _06827_/B vssd1 vssd1 vccd1 vccd1 _06828_/B sky130_fd_sc_hd__or2_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06758_ _10387_/Q _06791_/B _06747_/Y _06753_/Y _06757_/Y vssd1 vssd1 vccd1 vccd1
+ _06758_/X sky130_fd_sc_hd__a221o_1
X_09546_ _10382_/Q _10179_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09477_ _09467_/X _09476_/Y _09467_/X _09476_/Y vssd1 vssd1 vccd1 vccd1 _09477_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05709_ _10278_/Q vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__clkbuf_2
X_06689_ _10377_/Q _08707_/A vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__or2_2
X_08428_ _09957_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08428_/Y sky130_fd_sc_hd__nor2_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08359_ _09097_/A vssd1 vssd1 vccd1 vccd1 _09252_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10329_/CLK _10321_/D vssd1 vssd1 vccd1 vccd1 _10321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10252_ _10274_/CLK _10252_/D vssd1 vssd1 vccd1 vccd1 _10252_/Q sky130_fd_sc_hd__dfxtp_1
X_10183_ _10421_/CLK _10183_/D vssd1 vssd1 vccd1 vccd1 _10183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05991_ _05990_/A _05989_/X _10209_/Q _05990_/Y _05978_/X vssd1 vssd1 vccd1 vccd1
+ _10209_/D sky130_fd_sc_hd__o221a_1
XFILLER_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ _07650_/A _07650_/B _07652_/A vssd1 vssd1 vccd1 vccd1 _07730_/X sky130_fd_sc_hd__a21bo_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07661_ _07686_/B _07765_/A vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__or2_1
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09400_ _10228_/Q _09397_/Y _05941_/X _09398_/Y _09399_/X vssd1 vssd1 vccd1 vccd1
+ _09402_/A sky130_fd_sc_hd__a41o_1
X_06612_ _10390_/Q _10389_/Q _10388_/Q _10387_/Q vssd1 vssd1 vccd1 vccd1 _06613_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07592_ _09919_/X vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__inv_2
XFILLER_206_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06543_ _06543_/A vssd1 vssd1 vccd1 vccd1 _06543_/Y sky130_fd_sc_hd__inv_2
X_09331_ _09331_/A vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__inv_2
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06474_ _06474_/A _06474_/B vssd1 vssd1 vccd1 vccd1 _06482_/A sky130_fd_sc_hd__or2_1
X_08213_ _08213_/A vssd1 vssd1 vccd1 vccd1 _08213_/Y sky130_fd_sc_hd__inv_2
X_09193_ _09193_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__or2_1
XFILLER_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05425_ _05418_/B _05416_/X _05422_/Y _05392_/A _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05426_/A sky130_fd_sc_hd__o32a_1
XFILLER_174_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08144_ _10182_/Q vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__inv_2
X_05356_ _10335_/Q _05356_/B vssd1 vssd1 vccd1 vccd1 _05356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08075_/Y sky130_fd_sc_hd__nor2_1
X_05287_ _10340_/Q vssd1 vssd1 vccd1 vccd1 _05304_/A sky130_fd_sc_hd__inv_2
XFILLER_161_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07026_ _07020_/X _07025_/Y _07020_/X _07025_/Y vssd1 vssd1 vccd1 vccd1 _07026_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08977_ _08945_/X _08976_/X _08945_/X _08976_/X vssd1 vssd1 vccd1 vccd1 _08977_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__nand2_1
X_07859_ _07808_/X _07858_/X _07808_/X _07858_/X vssd1 vssd1 vccd1 vccd1 _07859_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09528_/X _06644_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09529_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10399_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _10422_/CLK _10304_/D vssd1 vssd1 vccd1 vccd1 _10304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10235_ _10414_/CLK _10235_/D vssd1 vssd1 vccd1 vccd1 _10235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10166_ _10334_/CLK _10166_/D vssd1 vssd1 vccd1 vccd1 _10166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10097_ _10176_/CLK _10097_/D vssd1 vssd1 vccd1 vccd1 _10097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06190_ _06204_/A vssd1 vssd1 vccd1 vccd1 _06190_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05210_ _05116_/X _10379_/Q _05203_/A _09746_/X _05206_/X vssd1 vssd1 vccd1 vccd1
+ _10379_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05141_ _10404_/Q vssd1 vssd1 vccd1 vccd1 _06615_/C sky130_fd_sc_hd__inv_2
XFILLER_128_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05072_ _05072_/A vssd1 vssd1 vccd1 vccd1 _05072_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09880_ _09879_/X _08314_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _08939_/C _08899_/X _08939_/C _08899_/X vssd1 vssd1 vccd1 vccd1 _08901_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_08831_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08831_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08762_ _08762_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__or2_1
X_05974_ _07483_/A _05970_/X input47/X _05971_/X _05960_/X vssd1 vssd1 vccd1 vccd1
+ _10216_/D sky130_fd_sc_hd__o221a_1
X_08693_ _08294_/A _10072_/Q _08134_/X _10071_/Q vssd1 vssd1 vccd1 vccd1 _08693_/X
+ sky130_fd_sc_hd__o22a_1
X_07713_ _07527_/A _07527_/B _07528_/B vssd1 vssd1 vccd1 vccd1 _07713_/X sky130_fd_sc_hd__a21bo_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07644_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07644_/X sky130_fd_sc_hd__or2_1
XFILLER_202_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07575_ _07563_/A _07563_/B _07648_/A vssd1 vssd1 vccd1 vccd1 _07578_/A sky130_fd_sc_hd__a21o_1
X_06526_ _10097_/Q _06464_/A _08423_/A _06434_/A vssd1 vssd1 vccd1 vccd1 _06539_/A
+ sky130_fd_sc_hd__a22o_1
X_09314_ _09314_/A _09254_/X vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__or2b_1
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _09245_/X sky130_fd_sc_hd__or3_1
X_06457_ _06454_/X _06456_/Y _06454_/X _06456_/Y vssd1 vssd1 vccd1 vccd1 _06457_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_193_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05408_ _06185_/A _05465_/A vssd1 vssd1 vccd1 vccd1 _05423_/A sky130_fd_sc_hd__or2_1
X_09176_ _09294_/C _09176_/B vssd1 vssd1 vccd1 vccd1 _09240_/A sky130_fd_sc_hd__or2_1
X_06388_ _10247_/Q _08405_/A vssd1 vssd1 vccd1 vccd1 _06391_/A sky130_fd_sc_hd__nor2_1
XFILLER_193_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08127_ _06755_/B _08545_/A _08760_/A _08121_/X _08126_/X vssd1 vssd1 vccd1 vccd1
+ _08143_/A sky130_fd_sc_hd__o221a_1
XFILLER_134_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05339_ _05339_/A vssd1 vssd1 vccd1 vccd1 _05340_/B sky130_fd_sc_hd__inv_2
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08058_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08063_/B sky130_fd_sc_hd__buf_1
XFILLER_122_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 _10024_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[0] sky130_fd_sc_hd__clkbuf_2
X_07009_ _07235_/A vssd1 vssd1 vccd1 vccd1 _07054_/A sky130_fd_sc_hd__buf_4
X_10020_ _08033_/X _07388_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__mux2_1
Xoutput69 _10025_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10218_ _10225_/CLK _10218_/D vssd1 vssd1 vccd1 vccd1 _10218_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _10330_/CLK _10149_/D vssd1 vssd1 vccd1 vccd1 _10149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05690_ _05694_/A _05690_/B vssd1 vssd1 vccd1 vccd1 _05690_/X sky130_fd_sc_hd__and2_1
XFILLER_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07360_ _07341_/X _07345_/X _07346_/X _07359_/X vssd1 vssd1 vccd1 vccd1 _07360_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06311_ _06311_/A _10132_/Q vssd1 vssd1 vccd1 vccd1 _06312_/B sky130_fd_sc_hd__nor2_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09030_ _05941_/X _09251_/A _09029_/X vssd1 vssd1 vccd1 vccd1 _09030_/Y sky130_fd_sc_hd__a21oi_1
X_07291_ _07288_/X _07290_/X _07288_/X _07290_/X vssd1 vssd1 vccd1 vccd1 _07291_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06242_ _10180_/Q vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__inv_2
XFILLER_175_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06173_ _06175_/A _09670_/X vssd1 vssd1 vccd1 vccd1 _10119_/D sky130_fd_sc_hd__and2_1
X_05124_ _05133_/A _05124_/B vssd1 vssd1 vccd1 vccd1 _10408_/D sky130_fd_sc_hd__nor2_1
XFILLER_171_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05055_ _05072_/A vssd1 vssd1 vccd1 vccd1 _05055_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09932_ _09931_/X _07830_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__mux2_1
X_09863_ _10374_/Q _09862_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09863_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08814_ _08179_/A _08790_/A _08788_/X _08792_/X vssd1 vssd1 vccd1 vccd1 _08815_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09794_ _08218_/Y _10357_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09794_/X sky130_fd_sc_hd__mux2_1
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _08745_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05957_ _05956_/X _05947_/X input45/X _05948_/X _05950_/X vssd1 vssd1 vccd1 vccd1
+ _10222_/D sky130_fd_sc_hd__o221a_1
X_08676_ _10064_/Q vssd1 vssd1 vccd1 vccd1 _08676_/Y sky130_fd_sc_hd__inv_2
X_05888_ _05888_/A vssd1 vssd1 vccd1 vccd1 _05888_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07627_ _07627_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07627_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07558_ _07830_/A _07558_/B _07558_/C vssd1 vssd1 vccd1 vccd1 _07558_/X sky130_fd_sc_hd__or3_1
XFILLER_41_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06509_ _06516_/C _06508_/X _06516_/C _06508_/X vssd1 vssd1 vccd1 vccd1 _06509_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_194_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07489_ _07485_/X _07488_/X _07485_/X _07488_/X vssd1 vssd1 vccd1 vccd1 _07496_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09228_ _09447_/A _09229_/B _09343_/A _09354_/D vssd1 vssd1 vccd1 vccd1 _09230_/A
+ sky130_fd_sc_hd__o22a_1
X_09159_ _09159_/A _09159_/B vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__or2_2
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10003_ _08009_/A _08044_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06860_ _10224_/Q vssd1 vssd1 vccd1 vccd1 _07212_/A sky130_fd_sc_hd__inv_2
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05811_ _07415_/A _10253_/Q vssd1 vssd1 vccd1 vccd1 _05811_/Y sky130_fd_sc_hd__nor2_1
X_06791_ _06795_/A _06791_/B vssd1 vssd1 vccd1 vccd1 _06791_/Y sky130_fd_sc_hd__nor2_1
X_08530_ _08533_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__and2_1
X_05742_ _10282_/Q _05741_/X _09644_/X _05732_/X _05737_/X vssd1 vssd1 vccd1 vccd1
+ _10282_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08461_ _08461_/A _10045_/Q vssd1 vssd1 vccd1 vccd1 _08461_/Y sky130_fd_sc_hd__nor2_4
X_05673_ _05673_/A _05673_/B vssd1 vssd1 vccd1 vccd1 _05673_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07412_ _07412_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__or2_1
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08392_ _08392_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08392_/Y sky130_fd_sc_hd__nor2_1
XFILLER_195_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07343_ _07016_/X _07342_/X _07016_/A _07342_/X vssd1 vssd1 vccd1 vccd1 _07343_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07274_ _07266_/Y _07270_/X _07272_/X _07273_/X vssd1 vssd1 vccd1 vccd1 _07274_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06225_ _06225_/A vssd1 vssd1 vccd1 vccd1 _06225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09091_/C _09012_/B _09055_/A vssd1 vssd1 vccd1 vccd1 _09013_/X sky130_fd_sc_hd__a21bo_1
X_06156_ _06156_/A vssd1 vssd1 vccd1 vccd1 _06156_/X sky130_fd_sc_hd__buf_1
XFILLER_208_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06087_ _06102_/A vssd1 vssd1 vccd1 vccd1 _06101_/A sky130_fd_sc_hd__inv_2
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05107_ _10208_/Q vssd1 vssd1 vccd1 vccd1 _05202_/A sky130_fd_sc_hd__buf_2
X_05038_ input19/X vssd1 vssd1 vccd1 vccd1 _05038_/X sky130_fd_sc_hd__buf_4
X_09915_ _08847_/B _07446_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__mux2_2
X_09846_ _08276_/X _10370_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09777_ _09776_/X input46/X _09781_/S vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06989_ _10225_/Q _07219_/B _07311_/A _07311_/B vssd1 vssd1 vccd1 vccd1 _06989_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08728_ _08724_/A _08742_/B _06632_/Y _08727_/Y vssd1 vssd1 vccd1 vccd1 _08728_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ _08130_/X _10046_/Q _08077_/X _10045_/Q _08657_/Y vssd1 vssd1 vccd1 vccd1
+ _08704_/C sky130_fd_sc_hd__a221o_1
XFILLER_202_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06010_ _09873_/X _05998_/X _06271_/A _06002_/X _06005_/X vssd1 vssd1 vccd1 vccd1
+ _10205_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07961_ _07878_/A _07868_/B _07878_/C _07867_/B vssd1 vssd1 vccd1 vccd1 _07961_/X
+ sky130_fd_sc_hd__o22a_1
X_09700_ _06553_/Y input33/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06912_ _07165_/A _06912_/B _06923_/A vssd1 vssd1 vccd1 vccd1 _06913_/A sky130_fd_sc_hd__and3_1
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07892_ _07792_/X _07891_/X _07792_/X _07891_/X vssd1 vssd1 vccd1 vccd1 _07892_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09631_ _06286_/Y _06289_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__mux2_1
X_06843_ _06911_/A vssd1 vssd1 vccd1 vccd1 _06962_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06774_ _10400_/Q _06807_/B _10399_/Q _06806_/B _06773_/Y vssd1 vssd1 vccd1 vccd1
+ _06774_/X sky130_fd_sc_hd__o221a_1
X_09562_ _09561_/X _10355_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09562_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08513_ _10195_/Q _08513_/B vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__nand2_2
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05725_ _10289_/Q _05715_/X _05800_/A _05719_/X _05724_/X vssd1 vssd1 vccd1 vccd1
+ _10289_/D sky130_fd_sc_hd__o221a_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09493_ _09492_/X _06640_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__mux2_2
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08444_ _08444_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08444_/Y sky130_fd_sc_hd__nor2_1
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05656_ _10307_/Q vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__inv_2
XFILLER_63_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08375_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__buf_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05587_ _09984_/X _05577_/X _05689_/A vssd1 vssd1 vccd1 vccd1 _05685_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07326_ _07320_/X _07325_/X _07320_/X _07325_/X vssd1 vssd1 vccd1 vccd1 _07326_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07257_ _07250_/X _07251_/X _07250_/X _07251_/X vssd1 vssd1 vccd1 vccd1 _07303_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06208_ _09696_/X _06203_/X _10097_/Q _06204_/X vssd1 vssd1 vccd1 vccd1 _10097_/D
+ sky130_fd_sc_hd__a22o_1
X_07188_ _07186_/X _07187_/X _07186_/X _07187_/X vssd1 vssd1 vccd1 vccd1 _07188_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06139_ _06157_/A vssd1 vssd1 vccd1 vccd1 _06156_/A sky130_fd_sc_hd__inv_2
XFILLER_2_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _09828_/X input28/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10397_ _10433_/CLK _10397_/D vssd1 vssd1 vccd1 vccd1 _10397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06490_ _08392_/A _06489_/X _06495_/A _06484_/X vssd1 vssd1 vccd1 vccd1 _06490_/Y
+ sky130_fd_sc_hd__o22ai_1
X_05510_ _05510_/A vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05441_ _10321_/Q _05441_/B vssd1 vssd1 vccd1 vccd1 _05441_/Y sky130_fd_sc_hd__nor2_1
X_08160_ _08765_/A vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__buf_2
XFILLER_158_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05372_ _05439_/A vssd1 vssd1 vccd1 vccd1 _05372_/X sky130_fd_sc_hd__clkbuf_2
X_07111_ _07111_/A _07111_/B vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__or2_1
X_08091_ _10376_/Q _08303_/A _06630_/Y _10200_/Q _08090_/X vssd1 vssd1 vccd1 vccd1
+ _08098_/C sky130_fd_sc_hd__o221a_1
XFILLER_173_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07042_ _06942_/X _07041_/X _06942_/X _07041_/X vssd1 vssd1 vccd1 vccd1 _07042_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ _09038_/A _09096_/A _08993_/C vssd1 vssd1 vccd1 vccd1 _08993_/X sky130_fd_sc_hd__or3_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07944_ _07709_/X _07756_/X _07709_/X _07756_/X vssd1 vssd1 vccd1 vccd1 _07944_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _07870_/X _07871_/X _07870_/X _07871_/X vssd1 vssd1 vccd1 vccd1 _07875_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ _06641_/Y _08104_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09614_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06826_ _06826_/A _06826_/B vssd1 vssd1 vccd1 vccd1 _06827_/B sky130_fd_sc_hd__or2_1
XFILLER_55_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06757_ _06757_/A vssd1 vssd1 vccd1 vccd1 _06757_/Y sky130_fd_sc_hd__inv_2
X_09545_ _09544_/X _10113_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06688_ _10376_/Q _08709_/A vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__or2_2
X_09476_ _09472_/X _09475_/Y _09472_/X _09475_/Y vssd1 vssd1 vccd1 vccd1 _09476_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_05708_ _10295_/Q _05701_/X _05786_/A _05705_/X _05660_/X vssd1 vssd1 vccd1 vccd1
+ _10295_/D sky130_fd_sc_hd__o221a_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08427_/Y sky130_fd_sc_hd__nor2_1
X_05639_ _10310_/Q _05467_/X _05637_/X _05638_/Y _05245_/X vssd1 vssd1 vccd1 vccd1
+ _10310_/D sky130_fd_sc_hd__o221a_1
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08358_ _10231_/Q vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__inv_2
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08289_ _08289_/A _08289_/B vssd1 vssd1 vccd1 vccd1 _08294_/B sky130_fd_sc_hd__or2_2
XFILLER_164_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07309_ _07309_/A _07309_/B vssd1 vssd1 vccd1 vccd1 _07309_/X sky130_fd_sc_hd__or2_1
XFILLER_192_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _10330_/CLK _10320_/D vssd1 vssd1 vccd1 vccd1 _10320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _10274_/CLK _10251_/D vssd1 vssd1 vccd1 vccd1 _10251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10182_ _10421_/CLK _10182_/D vssd1 vssd1 vccd1 vccd1 _10182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10449_ _10450_/CLK _10449_/D vssd1 vssd1 vccd1 vccd1 _10449_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05990_ _05990_/A vssd1 vssd1 vccd1 vccd1 _05990_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07660_ _07660_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__or2_2
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06611_ _10386_/Q _10385_/Q _10384_/Q vssd1 vssd1 vccd1 vccd1 _06613_/C sky130_fd_sc_hd__or3_1
X_07591_ _07591_/A _09921_/X vssd1 vssd1 vccd1 vccd1 _07597_/C sky130_fd_sc_hd__nor2_2
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06542_ _06542_/A _06542_/B vssd1 vssd1 vccd1 vccd1 _06543_/A sky130_fd_sc_hd__nand2_1
X_09330_ _09328_/X _09329_/X _09328_/X _09329_/X vssd1 vssd1 vccd1 vccd1 _09331_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__or2_1
XFILLER_178_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08212_ _08211_/A _08211_/B _08188_/X _08215_/B vssd1 vssd1 vccd1 vccd1 _08212_/X
+ sky130_fd_sc_hd__o211a_1
X_06473_ _06447_/X _06450_/X _06471_/X _06455_/X _06472_/X vssd1 vssd1 vccd1 vccd1
+ _06474_/B sky130_fd_sc_hd__o311a_1
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09192_ _09192_/A vssd1 vssd1 vccd1 vccd1 _09192_/Y sky130_fd_sc_hd__inv_2
X_05424_ _05424_/A vssd1 vssd1 vccd1 vccd1 _05424_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08143_ _08143_/A _08143_/B _08143_/C _08143_/D vssd1 vssd1 vccd1 vccd1 _08176_/C
+ sky130_fd_sc_hd__and4_1
X_05355_ _05355_/A vssd1 vssd1 vccd1 vccd1 _05356_/B sky130_fd_sc_hd__inv_2
XFILLER_174_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08074_ _08074_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08074_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05286_ _10341_/Q vssd1 vssd1 vccd1 vccd1 _05305_/A sky130_fd_sc_hd__inv_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07025_ _07021_/X _07024_/Y _07021_/X _07024_/Y vssd1 vssd1 vccd1 vccd1 _07025_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08976_ _08962_/X _08975_/X _08962_/X _08975_/X vssd1 vssd1 vccd1 vccd1 _08976_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07927_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__or2_1
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07858_ _07853_/Y _07857_/Y _07853_/Y _07857_/Y vssd1 vssd1 vccd1 vccd1 _07858_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06809_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07789_ _09908_/X vssd1 vssd1 vccd1 vccd1 _07789_/Y sky130_fd_sc_hd__inv_2
X_09528_ _06643_/Y _08093_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09455_/X _09458_/X _09455_/X _09458_/X vssd1 vssd1 vccd1 vccd1 _09459_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _10422_/CLK _10303_/D vssd1 vssd1 vccd1 vccd1 _10303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10234_ _10414_/CLK _10234_/D vssd1 vssd1 vccd1 vccd1 _10234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10165_ _10343_/CLK _10165_/D vssd1 vssd1 vccd1 vccd1 _10165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10096_ _10176_/CLK _10096_/D vssd1 vssd1 vccd1 vccd1 _10096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05140_ _05157_/A _05140_/B vssd1 vssd1 vccd1 vccd1 _10405_/D sky130_fd_sc_hd__nor2_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05071_ _10429_/Q _05064_/X input28/X _05065_/X _05070_/X vssd1 vssd1 vccd1 vccd1
+ _10429_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08830_ _08079_/X _08723_/Y _08281_/A _08720_/Y _08829_/X vssd1 vssd1 vccd1 vccd1
+ _08831_/B sky130_fd_sc_hd__o221a_1
XFILLER_97_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08761_ _08761_/A _08770_/A vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__or2_1
XFILLER_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05973_ _10216_/Q vssd1 vssd1 vccd1 vccd1 _07483_/A sky130_fd_sc_hd__buf_2
X_08692_ _08169_/X _10069_/Q _08162_/X _10070_/Q vssd1 vssd1 vccd1 vccd1 _08697_/A
+ sky130_fd_sc_hd__o22a_1
X_07712_ _07681_/X _07701_/X _07681_/X _07701_/X vssd1 vssd1 vccd1 vccd1 _07712_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07643_ _07640_/A _07640_/B _07640_/X vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__a21bo_1
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09313_ _09462_/C _09312_/Y _09462_/C _09312_/Y vssd1 vssd1 vccd1 vccd1 _09313_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07574_ _07574_/A vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__inv_2
X_06525_ _10097_/Q vssd1 vssd1 vccd1 vccd1 _08423_/A sky130_fd_sc_hd__inv_2
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ _09244_/A vssd1 vssd1 vccd1 vccd1 _09244_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06456_ _06447_/X _06450_/X _06455_/X vssd1 vssd1 vccd1 vccd1 _06456_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_193_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _09173_/X _09174_/X _09173_/X _09174_/X vssd1 vssd1 vccd1 vccd1 _09176_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05407_ _10328_/Q _05407_/B vssd1 vssd1 vccd1 vccd1 _05407_/Y sky130_fd_sc_hd__nor2_1
X_08126_ _10368_/Q _08269_/A _10364_/Q _08125_/X vssd1 vssd1 vccd1 vccd1 _08126_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06387_ _10140_/Q vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__inv_2
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05338_ _05338_/A vssd1 vssd1 vccd1 vccd1 _10340_/D sky130_fd_sc_hd__inv_2
X_05269_ _10350_/Q vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__buf_2
X_08057_ _10314_/Q _10007_/X vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__or2_2
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07008_ _07008_/A vssd1 vssd1 vccd1 vccd1 _07008_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput59 _09569_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08959_ _08959_/A vssd1 vssd1 vccd1 vccd1 _09001_/C sky130_fd_sc_hd__inv_2
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10217_/CLK _10217_/D vssd1 vssd1 vccd1 vccd1 _10217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10148_ _10330_/CLK _10148_/D vssd1 vssd1 vccd1 vccd1 _10148_/Q sky130_fd_sc_hd__dfxtp_1
X_10079_ _10176_/CLK _10079_/D vssd1 vssd1 vccd1 vccd1 _10079_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06310_ _10239_/Q vssd1 vssd1 vccd1 vccd1 _06311_/A sky130_fd_sc_hd__inv_2
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07290_ _05956_/X _07219_/B _07219_/A _07152_/D _07289_/X vssd1 vssd1 vccd1 vccd1
+ _07290_/X sky130_fd_sc_hd__a41o_1
XFILLER_175_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06241_ _08380_/A vssd1 vssd1 vccd1 vccd1 _09544_/S sky130_fd_sc_hd__buf_2
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06172_ _06175_/A _09671_/X vssd1 vssd1 vccd1 vccd1 _10120_/D sky130_fd_sc_hd__and2_1
XFILLER_190_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05123_ _05116_/X _06614_/C _05122_/Y _05113_/X vssd1 vssd1 vccd1 vccd1 _05124_/B
+ sky130_fd_sc_hd__o22a_1
X_05054_ _10439_/Q _05047_/X input39/X _05048_/X _05053_/X vssd1 vssd1 vccd1 vccd1
+ _10439_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09931_ _09930_/X _07118_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09862_ _08292_/X _10374_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09862_/X sky130_fd_sc_hd__mux2_1
X_08813_ _08160_/X _08766_/A _06254_/A _08756_/A _08769_/X vssd1 vssd1 vccd1 vccd1
+ _08821_/A sky130_fd_sc_hd__a221o_1
X_09793_ _09792_/X input50/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _08521_/A _08739_/Y _08809_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08824_/A
+ sky130_fd_sc_hd__a22o_1
X_05956_ _10222_/Q vssd1 vssd1 vccd1 vccd1 _05956_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08675_ _08172_/X _10061_/Q _08079_/X _10068_/Q vssd1 vssd1 vccd1 vccd1 _08680_/B
+ sky130_fd_sc_hd__a22o_1
X_05887_ _07660_/A vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__buf_2
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10202_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_198_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__nor2_4
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ _07557_/A vssd1 vssd1 vccd1 vccd1 _07558_/C sky130_fd_sc_hd__inv_2
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06508_ _06516_/A _06516_/B _06499_/Y _06507_/X vssd1 vssd1 vccd1 vccd1 _06508_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_194_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_29_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10414_/CLK sky130_fd_sc_hd__clkbuf_16
X_07488_ _07868_/A _07537_/D vssd1 vssd1 vccd1 vccd1 _07488_/X sky130_fd_sc_hd__or2_1
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09227_ _05922_/X _09142_/X _09225_/X _09283_/A vssd1 vssd1 vccd1 vccd1 _09227_/X
+ sky130_fd_sc_hd__a31o_1
X_06439_ _06421_/Y _06438_/X _06445_/A vssd1 vssd1 vccd1 vccd1 _06439_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ _09122_/A _09108_/Y _09043_/A _09109_/X vssd1 vssd1 vccd1 vccd1 _09159_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08109_ _08753_/A _08104_/X _06642_/Y _06254_/A _08108_/X vssd1 vssd1 vccd1 vccd1
+ _08119_/B sky130_fd_sc_hd__o221a_1
X_09089_ _09259_/A _09089_/B vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__or2_2
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10002_ _08015_/A _08054_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _10002_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05810_ _10271_/Q _10254_/Q _07434_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _05810_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06790_ _09717_/S _06790_/B vssd1 vssd1 vccd1 vccd1 _06790_/X sky130_fd_sc_hd__and2_1
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05741_ _05741_/A vssd1 vssd1 vccd1 vccd1 _05741_/X sky130_fd_sc_hd__clkbuf_2
X_08460_ _10046_/Q vssd1 vssd1 vccd1 vccd1 _08460_/Y sky130_fd_sc_hd__inv_2
X_05672_ _05672_/A vssd1 vssd1 vccd1 vccd1 _05672_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ _09629_/X _08391_/B vssd1 vssd1 vccd1 vccd1 _08391_/Y sky130_fd_sc_hd__nor2_1
X_07411_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__or2_1
XFILLER_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07342_ _06923_/A _06923_/B _06924_/B vssd1 vssd1 vccd1 vccd1 _07342_/X sky130_fd_sc_hd__a21bo_1
XFILLER_149_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _07266_/Y _07270_/X _07266_/Y _07270_/X vssd1 vssd1 vccd1 vccd1 _07273_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06224_ _06224_/A vssd1 vssd1 vccd1 vccd1 _06224_/X sky130_fd_sc_hd__clkbuf_2
X_09012_ _09091_/C _09012_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__or2_2
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06155_ _09651_/X _06148_/X _10133_/Q _06149_/X _06154_/X vssd1 vssd1 vccd1 vccd1
+ _10133_/D sky130_fd_sc_hd__o221a_1
X_05106_ _10410_/Q vssd1 vssd1 vccd1 vccd1 _06614_/A sky130_fd_sc_hd__inv_2
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06086_ _06086_/A _09897_/X vssd1 vssd1 vccd1 vccd1 _06102_/A sky130_fd_sc_hd__or2_2
XFILLER_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05037_ _10444_/Q _05012_/A input49/X _05013_/A _05036_/X vssd1 vssd1 vccd1 vccd1
+ _10444_/D sky130_fd_sc_hd__o221a_1
X_09914_ _05852_/X _07444_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09914_/X sky130_fd_sc_hd__mux2_2
X_09845_ _09844_/X input33/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09776_ _09775_/X _08202_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09776_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06988_ _07152_/B vssd1 vssd1 vccd1 vccd1 _07219_/B sky130_fd_sc_hd__clkbuf_2
X_08727_ _08727_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08727_/Y sky130_fd_sc_hd__nor2_1
X_05939_ _10227_/Q vssd1 vssd1 vccd1 vccd1 _05939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08658_ _08116_/X _08456_/X _08554_/A _10047_/Q vssd1 vssd1 vccd1 vccd1 _08658_/X
+ sky130_fd_sc_hd__o22a_1
X_07609_ _07596_/A _07596_/B _07596_/X vssd1 vssd1 vccd1 vccd1 _07610_/B sky130_fd_sc_hd__a21bo_1
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08589_ _08589_/A _08589_/B _08588_/X vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__or3b_1
XFILLER_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07960_ _07956_/X _07957_/X _07956_/X _07957_/X vssd1 vssd1 vccd1 vccd1 _07960_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06911_ _06911_/A _06911_/B vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__or2_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07891_ _07882_/A _07882_/B _07882_/X vssd1 vssd1 vccd1 vccd1 _07891_/X sky130_fd_sc_hd__a21bo_1
XFILLER_82_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09630_ _06278_/X _06279_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__mux2_1
X_06842_ _07125_/A vssd1 vssd1 vccd1 vccd1 _06911_/A sky130_fd_sc_hd__buf_1
X_06773_ _05168_/Y _06718_/A _06616_/D _06713_/A _06772_/Y vssd1 vssd1 vccd1 vccd1
+ _06773_/Y sky130_fd_sc_hd__o221ai_1
X_09561_ _10387_/Q _10184_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09561_/X sky130_fd_sc_hd__mux2_1
X_08512_ _10064_/Q _08482_/B _08511_/Y vssd1 vssd1 vccd1 vccd1 _08513_/B sky130_fd_sc_hd__a21oi_2
X_05724_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05724_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09492_ _06639_/Y _08107_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08443_ _09602_/X _08449_/B vssd1 vssd1 vccd1 vccd1 _08443_/Y sky130_fd_sc_hd__nor2_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05655_ _05655_/A _05655_/B vssd1 vssd1 vccd1 vccd1 _05655_/X sky130_fd_sc_hd__and2_1
XFILLER_211_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08374_ _10233_/Q vssd1 vssd1 vccd1 vccd1 _09258_/A sky130_fd_sc_hd__inv_2
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05586_ _05694_/A _05690_/B vssd1 vssd1 vccd1 vccd1 _05689_/A sky130_fd_sc_hd__or2_1
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07325_ _07321_/X _07322_/X _07323_/X _07324_/X vssd1 vssd1 vccd1 vccd1 _07325_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07256_ _07252_/X _07255_/X _07252_/X _07255_/X vssd1 vssd1 vccd1 vccd1 _07256_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06207_ _09697_/X _06203_/X _10098_/Q _06204_/X vssd1 vssd1 vccd1 vccd1 _10098_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _07137_/A _07137_/B _07138_/B vssd1 vssd1 vccd1 vccd1 _07187_/X sky130_fd_sc_hd__a21bo_1
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06138_ _06083_/A _08319_/A _10266_/Q vssd1 vssd1 vccd1 vccd1 _06157_/A sky130_fd_sc_hd__o21ai_4
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06069_ _06069_/A vssd1 vssd1 vccd1 vccd1 _06069_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09828_ _09827_/X _08256_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ _10348_/Q _09758_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10396_ _10433_/CLK _10396_/D vssd1 vssd1 vccd1 vccd1 _10396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05440_ _05440_/A vssd1 vssd1 vccd1 vccd1 _05441_/B sky130_fd_sc_hd__inv_2
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05371_ _09897_/X _05465_/A vssd1 vssd1 vccd1 vccd1 _05439_/A sky130_fd_sc_hd__or2_1
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07110_ _06887_/A _09889_/X _07112_/A _09890_/X _07109_/Y vssd1 vssd1 vccd1 vccd1
+ _07111_/B sky130_fd_sc_hd__o41a_1
X_08090_ _06699_/Y _10203_/Q _08762_/A _08081_/X vssd1 vssd1 vccd1 vccd1 _08090_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07041_ _07039_/X _07040_/X _07039_/X _07040_/X vssd1 vssd1 vccd1 vccd1 _07041_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _09977_/X vssd1 vssd1 vccd1 vccd1 _09096_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_141_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ _07867_/X _07892_/X _07867_/X _07892_/X vssd1 vssd1 vccd1 vccd1 _07943_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07874_ _07872_/X _07873_/X _07872_/X _07873_/X vssd1 vssd1 vccd1 vccd1 _07874_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09613_ _10426_/Q _09613_/A1 _09899_/S vssd1 vssd1 vccd1 vccd1 _09613_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06825_ _06824_/X _05888_/Y _06820_/B vssd1 vssd1 vccd1 vccd1 _06825_/Y sky130_fd_sc_hd__o21ai_1
X_06756_ _06750_/Y _06755_/Y _06789_/B _06748_/Y _06790_/B vssd1 vssd1 vccd1 vccd1
+ _06757_/A sky130_fd_sc_hd__o32a_1
X_09544_ _10081_/Q _10175_/Q _09544_/S vssd1 vssd1 vccd1 vccd1 _09544_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06687_ _10375_/Q _08711_/A vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__or2_2
X_09475_ _09473_/X _09474_/X _09473_/X _09474_/X vssd1 vssd1 vccd1 vccd1 _09475_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_05707_ _10279_/Q vssd1 vssd1 vccd1 vccd1 _05786_/A sky130_fd_sc_hd__clkbuf_2
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08426_ _09951_/X _08435_/B vssd1 vssd1 vccd1 vccd1 _08426_/X sky130_fd_sc_hd__and2_1
X_05638_ _05549_/X _05605_/X _05549_/X _05605_/X vssd1 vssd1 vccd1 vccd1 _05638_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08357_ _08357_/A _09544_/S vssd1 vssd1 vccd1 vccd1 _08357_/Y sky130_fd_sc_hd__nor2_1
X_05569_ _09974_/X _05568_/X _09974_/X _05568_/X vssd1 vssd1 vccd1 vccd1 _05673_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ _08134_/X _08283_/Y _06269_/B vssd1 vssd1 vccd1 vccd1 _08288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_149_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07308_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07309_/B sky130_fd_sc_hd__or2_1
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07239_ _07239_/A vssd1 vssd1 vccd1 vccd1 _07241_/A sky130_fd_sc_hd__inv_2
XFILLER_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _10274_/CLK _10250_/D vssd1 vssd1 vccd1 vccd1 _10250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10421_/CLK _10181_/D vssd1 vssd1 vccd1 vccd1 _10181_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10448_ _10450_/CLK _10448_/D vssd1 vssd1 vccd1 vccd1 _10448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _10421_/CLK _10379_/D vssd1 vssd1 vccd1 vccd1 _10379_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06610_ _10398_/Q _10397_/Q _10396_/Q _10395_/Q vssd1 vssd1 vccd1 vccd1 _06613_/B
+ sky130_fd_sc_hd__or4_4
X_07590_ _07588_/X _07589_/X _07588_/X _07589_/X vssd1 vssd1 vccd1 vccd1 _07596_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06541_ _08423_/A _06540_/X _08425_/A _06540_/X _06529_/B vssd1 vssd1 vccd1 vccd1
+ _06542_/B sky130_fd_sc_hd__o221a_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _09260_/A vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__inv_2
X_06472_ _08373_/A _06487_/A _08382_/A _06430_/A vssd1 vssd1 vccd1 vccd1 _06472_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__nand2_2
X_05423_ _05423_/A vssd1 vssd1 vccd1 vccd1 _05424_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09191_ _09189_/X _09190_/X _09189_/X _09190_/X vssd1 vssd1 vccd1 vccd1 _09191_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08142_ _10351_/Q _08138_/X _08759_/A _08797_/A _08141_/X vssd1 vssd1 vccd1 vccd1
+ _08143_/D sky130_fd_sc_hd__o221a_1
X_05354_ _05354_/A vssd1 vssd1 vccd1 vccd1 _10336_/D sky130_fd_sc_hd__inv_2
X_08073_ _08073_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08073_/Y sky130_fd_sc_hd__nor2_1
X_05285_ _10342_/Q vssd1 vssd1 vccd1 vccd1 _05306_/A sky130_fd_sc_hd__inv_2
XFILLER_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07024_ _07022_/Y _07023_/X _07022_/Y _07023_/X vssd1 vssd1 vccd1 vccd1 _07024_/Y
+ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08975_ _08943_/A _08943_/B _08974_/A _08943_/Y _08974_/Y vssd1 vssd1 vccd1 vccd1
+ _08975_/X sky130_fd_sc_hd__o32a_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07926_ _07918_/Y _07925_/X _07918_/Y _07925_/X vssd1 vssd1 vccd1 vccd1 _07928_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07857_ _07854_/X _07856_/X _07854_/X _07856_/X vssd1 vssd1 vccd1 vccd1 _07857_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_204_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06808_ _06808_/A _06808_/B vssd1 vssd1 vccd1 vccd1 _06808_/Y sky130_fd_sc_hd__nor2_1
X_07788_ _07878_/D vssd1 vssd1 vccd1 vccd1 _07788_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _09526_/X _06636_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09527_/X sky130_fd_sc_hd__mux2_2
X_06739_ _06739_/A _06740_/A vssd1 vssd1 vccd1 vccd1 _06739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09456_/Y _09457_/Y _09456_/Y _09457_/Y vssd1 vssd1 vccd1 vccd1 _09458_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09389_ _09229_/X _09344_/X _09345_/X _09346_/X vssd1 vssd1 vccd1 vccd1 _09389_/X
+ sky130_fd_sc_hd__o22a_1
X_08409_ _08409_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08409_/X sky130_fd_sc_hd__or2_1
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ _10420_/CLK _10302_/D vssd1 vssd1 vccd1 vccd1 _10302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _10312_/CLK _10233_/D vssd1 vssd1 vccd1 vccd1 _10233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _10334_/CLK _10164_/D vssd1 vssd1 vccd1 vccd1 _10164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10095_ _10176_/CLK _10095_/D vssd1 vssd1 vccd1 vccd1 _10095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05070_ _05189_/A vssd1 vssd1 vccd1 vccd1 _05070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08760_ _08760_/A _08760_/B vssd1 vssd1 vccd1 vccd1 _08770_/A sky130_fd_sc_hd__or2_1
X_05972_ _05966_/X _05970_/X input48/X _05971_/X _05960_/X vssd1 vssd1 vccd1 vccd1
+ _10217_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08691_ _08304_/A _10074_/Q _08297_/A _10073_/Q vssd1 vssd1 vccd1 vccd1 _08694_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07711_ _07581_/X _07652_/X _07581_/X _07652_/X vssd1 vssd1 vccd1 vccd1 _07711_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07642_ _07637_/X _07641_/X _07637_/X _07641_/X vssd1 vssd1 vccd1 vccd1 _07642_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09312_ _09452_/A _09282_/A _09311_/Y vssd1 vssd1 vccd1 vccd1 _09312_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ _07573_/A _07579_/A vssd1 vssd1 vccd1 vccd1 _07573_/Y sky130_fd_sc_hd__nor2_1
X_06524_ _06527_/B _06523_/Y _06527_/B _06523_/Y vssd1 vssd1 vccd1 vccd1 _06524_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09243_ _09208_/X _09209_/X _09210_/X _09211_/X vssd1 vssd1 vccd1 vccd1 _09244_/A
+ sky130_fd_sc_hd__o22a_1
X_06455_ _08357_/A _06430_/A _08365_/A _06430_/A vssd1 vssd1 vccd1 vccd1 _06455_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09174_ _09174_/A _09918_/X _09174_/C vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__or3_1
X_06386_ _06384_/A _06381_/X _06384_/A _06381_/X vssd1 vssd1 vccd1 vccd1 _06386_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_05406_ _05406_/A vssd1 vssd1 vccd1 vccd1 _05407_/B sky130_fd_sc_hd__inv_2
X_08125_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08125_/X sky130_fd_sc_hd__buf_2
XFILLER_147_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05337_ _05330_/B _05333_/X _05335_/Y _05336_/X _05304_/A vssd1 vssd1 vccd1 vccd1
+ _05338_/A sky130_fd_sc_hd__o32a_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05268_ _05028_/X _05263_/X _10351_/Q _05264_/X _05265_/X vssd1 vssd1 vccd1 vccd1
+ _10351_/D sky130_fd_sc_hd__a221o_1
X_08056_ _07921_/A _07878_/A _08001_/X _08014_/A vssd1 vssd1 vccd1 vccd1 _08056_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_134_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05199_ _05193_/X _10387_/Q _05194_/X _09606_/X _05198_/X vssd1 vssd1 vccd1 vccd1
+ _10387_/D sky130_fd_sc_hd__o221a_1
X_07007_ _10225_/Q _07082_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__a21oi_4
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _09128_/A vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__inv_2
XFILLER_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08889_ _08889_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__or2_1
X_07909_ _05966_/X _07516_/B _07913_/A _07780_/Y vssd1 vssd1 vccd1 vccd1 _07909_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10216_ _10217_/CLK _10216_/D vssd1 vssd1 vccd1 vccd1 _10216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10147_ _10330_/CLK _10147_/D vssd1 vssd1 vccd1 vccd1 _10147_/Q sky130_fd_sc_hd__dfxtp_1
X_10078_ _10205_/CLK _10078_/D vssd1 vssd1 vccd1 vccd1 _10078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06240_ _06240_/A vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__inv_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06171_ _06175_/A _09672_/X vssd1 vssd1 vccd1 vccd1 _10121_/D sky130_fd_sc_hd__and2_1
X_05122_ _10440_/Q vssd1 vssd1 vccd1 vccd1 _05122_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05053_ _05189_/A vssd1 vssd1 vccd1 vccd1 _05053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _09929_/X _09451_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09861_ _09860_/X input37/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08812_ _08824_/C _08812_/B vssd1 vssd1 vccd1 vccd1 _08812_/X sky130_fd_sc_hd__or2_1
X_09792_ _09791_/X _08217_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08743_ _06636_/Y _08742_/Y _08738_/Y vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__o21bai_1
X_05955_ _07219_/A _05947_/X _05093_/X _05948_/X _05950_/X vssd1 vssd1 vccd1 vccd1
+ _10223_/D sky130_fd_sc_hd__o221a_1
X_08674_ _08674_/A _08674_/B _08674_/C _08673_/X vssd1 vssd1 vccd1 vccd1 _08680_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05886_ _10252_/Q _05871_/X _05699_/X _06820_/A _05885_/X vssd1 vssd1 vccd1 vccd1
+ _10252_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ _07625_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__or2_4
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07556_ _07811_/A _09935_/X vssd1 vssd1 vccd1 vccd1 _07557_/A sky130_fd_sc_hd__or2_2
XFILLER_194_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06507_ _08403_/A _06496_/X _08407_/A _06496_/X vssd1 vssd1 vccd1 vccd1 _06507_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _09142_/X _09225_/X _09170_/A vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__o21ai_2
X_07487_ _07672_/A vssd1 vssd1 vccd1 vccd1 _07868_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_194_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06438_ _06489_/A vssd1 vssd1 vccd1 vccd1 _06438_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09157_ _09127_/X _09156_/X _09127_/X _09156_/X vssd1 vssd1 vccd1 vccd1 _09159_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06369_ _10245_/Q vssd1 vssd1 vccd1 vccd1 _06370_/A sky130_fd_sc_hd__inv_2
XFILLER_181_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08108_ _06640_/Y _10189_/Q _10360_/Q _08107_/X vssd1 vssd1 vccd1 vccd1 _08108_/X
+ sky130_fd_sc_hd__o22a_1
X_09088_ _09087_/A _09087_/B _09187_/A vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__a21bo_1
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08039_ _07408_/A _07408_/B _07409_/B vssd1 vssd1 vccd1 vccd1 _08039_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10001_ _08053_/Y _07401_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__mux2_2
XFILLER_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05740_ _05581_/X _05728_/X _07594_/C _05732_/X _05737_/X vssd1 vssd1 vccd1 vccd1
+ _10283_/D sky130_fd_sc_hd__o221a_1
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05671_ _05677_/A _05671_/B vssd1 vssd1 vccd1 vccd1 _10304_/D sky130_fd_sc_hd__nor2_1
X_08390_ _08390_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__or2_1
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07410_ _07410_/A _07410_/B vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__or2_1
XFILLER_211_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07341_ _07336_/X _07338_/X _07336_/X _07338_/X vssd1 vssd1 vccd1 vccd1 _07341_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ _05956_/X _07082_/B _07219_/A _07189_/Y _07271_/X vssd1 vssd1 vccd1 vccd1
+ _07272_/X sky130_fd_sc_hd__a41o_1
XFILLER_191_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ _09009_/X _09010_/X _09009_/X _09010_/X vssd1 vssd1 vccd1 vccd1 _09012_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_06223_ _09685_/X _06217_/X _10086_/Q _06218_/X vssd1 vssd1 vccd1 vccd1 _10086_/D
+ sky130_fd_sc_hd__a22o_1
X_06154_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05105_ _05105_/A vssd1 vssd1 vccd1 vccd1 _05133_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06085_ _05322_/X _09943_/S input41/X _06084_/A _05993_/X vssd1 vssd1 vccd1 vccd1
+ _10175_/D sky130_fd_sc_hd__o221a_1
X_09913_ _09485_/X _09484_/Y _09994_/S vssd1 vssd1 vccd1 vccd1 _09913_/X sky130_fd_sc_hd__mux2_2
XFILLER_144_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05036_ _06176_/A vssd1 vssd1 vccd1 vccd1 _05036_/X sky130_fd_sc_hd__buf_2
X_09844_ _09843_/X _08274_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09775_ _10352_/Q _09774_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06987_ _09886_/X vssd1 vssd1 vccd1 vccd1 _07152_/B sky130_fd_sc_hd__inv_2
X_08726_ _08726_/A vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05938_ _10228_/Q _05927_/A _05032_/X _05928_/A _05934_/X vssd1 vssd1 vccd1 vccd1
+ _10228_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08657_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08657_/Y sky130_fd_sc_hd__nor2_1
X_05869_ _05869_/A vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__inv_2
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07608_ _07608_/A _07587_/X vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__or2b_1
XFILLER_186_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08588_ _08545_/A _08545_/B _08545_/Y _08569_/Y _08551_/A vssd1 vssd1 vccd1 vccd1
+ _08588_/X sky130_fd_sc_hd__o2111a_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ _07603_/A _07539_/B _07813_/C _09936_/X vssd1 vssd1 vccd1 vccd1 _07539_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_210_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09209_ _09141_/X _09151_/X _09131_/X _09152_/X vssd1 vssd1 vccd1 vccd1 _09209_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_182_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10436_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06910_ _06897_/X _06898_/X _06897_/X _06898_/X vssd1 vssd1 vccd1 vccd1 _06910_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_07890_ _07886_/X _07887_/X _07886_/X _07887_/X vssd1 vssd1 vccd1 vccd1 _07894_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10300_/CLK sky130_fd_sc_hd__clkbuf_16
X_06841_ _07146_/A vssd1 vssd1 vccd1 vccd1 _07125_/A sky130_fd_sc_hd__buf_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06772_ _10397_/Q _06804_/B _10398_/Q _06805_/B _06771_/X vssd1 vssd1 vccd1 vccd1
+ _06772_/Y sky130_fd_sc_hd__o221ai_1
X_09560_ _08382_/Y _10118_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09560_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _08511_/A vssd1 vssd1 vccd1 vccd1 _08511_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09491_ _10413_/Q _08061_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09491_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05723_ _10273_/Q vssd1 vssd1 vccd1 vccd1 _05800_/A sky130_fd_sc_hd__buf_2
X_08442_ _08442_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05654_ _05654_/A vssd1 vssd1 vccd1 vccd1 _05654_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08373_ _08373_/A _09544_/S vssd1 vssd1 vccd1 vccd1 _08373_/Y sky130_fd_sc_hd__nor2_1
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05585_ _09984_/X _05577_/X _09984_/X _05577_/X vssd1 vssd1 vccd1 vccd1 _05690_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _07308_/A _07308_/B _07309_/B vssd1 vssd1 vccd1 vccd1 _07324_/X sky130_fd_sc_hd__a21bo_1
XFILLER_176_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07255_ _07254_/A _07254_/B _07254_/X vssd1 vssd1 vccd1 vccd1 _07255_/X sky130_fd_sc_hd__a21bo_1
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06206_ _09698_/X _06203_/X _10099_/Q _06204_/X vssd1 vssd1 vccd1 vccd1 _10099_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07186_ _07162_/X _07183_/X _07162_/X _07183_/X vssd1 vssd1 vccd1 vccd1 _07186_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06137_ _06137_/A _06137_/B vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__or2_2
X_06068_ _10182_/Q vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05019_ input52/X vssd1 vssd1 vccd1 vccd1 _05034_/A sky130_fd_sc_hd__inv_2
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _10365_/Q _09826_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09827_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09758_ _08184_/B _10348_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08709_ _08709_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08709_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09689_ _06491_/X input21/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09689_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10395_ _10433_/CLK _10395_/D vssd1 vssd1 vccd1 vccd1 _10395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05370_ _05399_/A vssd1 vssd1 vccd1 vccd1 _05465_/A sky130_fd_sc_hd__inv_2
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07040_ _07056_/A _06868_/Y _05956_/X _06870_/Y _06880_/Y vssd1 vssd1 vccd1 vccd1
+ _07040_/X sky130_fd_sc_hd__a41o_1
XFILLER_141_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08991_ _08912_/X _08966_/X _08967_/X _08968_/Y vssd1 vssd1 vccd1 vccd1 _08991_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07942_ _07913_/A _07913_/B _07913_/Y vssd1 vssd1 vccd1 vccd1 _07942_/Y sky130_fd_sc_hd__o21ai_1
X_07873_ _07483_/A _07800_/X _07885_/A _07864_/Y _07869_/Y vssd1 vssd1 vccd1 vccd1
+ _07873_/X sky130_fd_sc_hd__a41o_1
X_09612_ _10425_/Q _08075_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09612_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06824_ _07234_/B vssd1 vssd1 vccd1 vccd1 _06824_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09543_ _09542_/X _10349_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06755_ _10386_/Q _06755_/B vssd1 vssd1 vccd1 vccd1 _06755_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _10374_/Q _08713_/A vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__or2_2
X_09474_ _09474_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09474_/X sky130_fd_sc_hd__or2_1
X_05706_ _10296_/Q _05701_/X _05704_/X _05705_/X _05660_/X vssd1 vssd1 vccd1 vccd1
+ _10296_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08425_ _08425_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08425_/Y sky130_fd_sc_hd__nor2_1
X_05637_ _05863_/A vssd1 vssd1 vccd1 vccd1 _05637_/X sky130_fd_sc_hd__buf_2
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _09912_/X _08364_/B vssd1 vssd1 vccd1 vccd1 _08356_/Y sky130_fd_sc_hd__nor2_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _07254_/X _07306_/X _07254_/X _07306_/X vssd1 vssd1 vccd1 vccd1 _07308_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_05568_ _05491_/X _05519_/X _05491_/X _05519_/X vssd1 vssd1 vccd1 vccd1 _05568_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08287_ _08162_/X _08285_/B _08193_/X _08286_/Y vssd1 vssd1 vccd1 vccd1 _08287_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05499_ _10218_/Q vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__inv_2
X_07238_ _07224_/X _07225_/X _07224_/X _07225_/X vssd1 vssd1 vccd1 vccd1 _07239_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07169_ _07160_/A _07166_/Y _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07182_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_160_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10180_ _10447_/CLK _10180_/D vssd1 vssd1 vccd1 vccd1 _10180_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ _10447_/CLK _10447_/D vssd1 vssd1 vccd1 vccd1 _10447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10378_ _10442_/CLK _10378_/D vssd1 vssd1 vccd1 vccd1 _10378_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06540_ _06540_/A vssd1 vssd1 vccd1 vccd1 _06540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06471_ _06471_/A _06454_/X vssd1 vssd1 vccd1 vccd1 _06471_/X sky130_fd_sc_hd__or2b_1
X_08210_ _08086_/X _08206_/Y _06251_/B vssd1 vssd1 vccd1 vccd1 _08210_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05422_ _10325_/Q _05422_/B vssd1 vssd1 vccd1 vccd1 _05422_/Y sky130_fd_sc_hd__nor2_1
X_09190_ _09245_/A _09245_/B _09190_/C vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__or3_1
X_08141_ _10369_/Q _08273_/A _06631_/Y _06026_/X vssd1 vssd1 vccd1 vccd1 _08141_/X
+ sky130_fd_sc_hd__o22a_1
X_05353_ _05348_/B _05333_/X _05352_/Y _05336_/X _05300_/A vssd1 vssd1 vccd1 vccd1
+ _05354_/A sky130_fd_sc_hd__o32a_1
XFILLER_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08072_ _08075_/B _10310_/Q vssd1 vssd1 vccd1 vccd1 _08072_/Y sky130_fd_sc_hd__nor2b_1
X_05284_ _10343_/Q vssd1 vssd1 vccd1 vccd1 _05307_/A sky130_fd_sc_hd__inv_2
X_07023_ _07023_/A _07023_/B _07023_/C _10022_/S vssd1 vssd1 vccd1 vccd1 _07023_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_161_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08974_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07925_ _07506_/A _07924_/X _07506_/A _07924_/X vssd1 vssd1 vccd1 vccd1 _07925_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07856_ _07878_/C _09908_/X vssd1 vssd1 vccd1 vccd1 _07856_/X sky130_fd_sc_hd__or2_1
X_06807_ _06808_/A _06807_/B vssd1 vssd1 vccd1 vccd1 _06807_/Y sky130_fd_sc_hd__nor2_1
X_04999_ _06184_/A vssd1 vssd1 vccd1 vccd1 _06083_/A sky130_fd_sc_hd__buf_2
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07787_ _09904_/X vssd1 vssd1 vccd1 vccd1 _07878_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_09526_ _05181_/Y _08172_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__mux2_1
X_06738_ _06661_/X _06737_/X _06661_/X _06737_/X vssd1 vssd1 vccd1 vccd1 _06740_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09457_/A _09457_/B _09457_/C _09994_/S vssd1 vssd1 vccd1 vccd1 _09457_/Y
+ sky130_fd_sc_hd__nor4_2
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _09493_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08408_/Y sky130_fd_sc_hd__nor2_2
X_06669_ _10357_/Q _06669_/B vssd1 vssd1 vccd1 vccd1 _06670_/B sky130_fd_sc_hd__or2_2
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09388_ _09336_/A _09336_/B _09387_/A _09457_/A _09457_/B vssd1 vssd1 vccd1 vccd1
+ _09388_/X sky130_fd_sc_hd__a32o_1
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08339_ _10228_/Q vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__inv_2
XFILLER_137_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _10422_/CLK _10301_/D vssd1 vssd1 vccd1 vccd1 _10301_/Q sky130_fd_sc_hd__dfxtp_1
X_10232_ _10312_/CLK _10232_/D vssd1 vssd1 vccd1 vccd1 _10232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10163_ _10334_/CLK _10163_/D vssd1 vssd1 vccd1 vccd1 _10163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10094_ _10176_/CLK _10094_/D vssd1 vssd1 vccd1 vccd1 _10094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05971_ _05971_/A vssd1 vssd1 vccd1 vccd1 _05971_/X sky130_fd_sc_hd__buf_1
X_07710_ _07703_/X _07704_/X _07703_/X _07704_/X vssd1 vssd1 vccd1 vccd1 _07710_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08690_ _08134_/X _10071_/Q _08162_/X _10070_/Q vssd1 vssd1 vccd1 vccd1 _08697_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07641_ _07638_/X _07640_/X _07638_/X _07640_/X vssd1 vssd1 vccd1 vccd1 _07641_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ _07557_/A _07567_/Y _07564_/X _07568_/X vssd1 vssd1 vccd1 vccd1 _07579_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_179_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09311_ _09311_/A vssd1 vssd1 vccd1 vccd1 _09311_/Y sky130_fd_sc_hd__inv_2
X_06523_ _08418_/A _06438_/X _06527_/A vssd1 vssd1 vccd1 vccd1 _06523_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ _09227_/X _09241_/X _09227_/X _09241_/X vssd1 vssd1 vccd1 vccd1 _09242_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06454_ _10085_/Q _06460_/A _08373_/A _06442_/X vssd1 vssd1 vccd1 vccd1 _06454_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_178_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _09289_/A _09983_/X vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__or2_2
X_05405_ _05396_/A _05401_/Y _05404_/Y _05400_/X vssd1 vssd1 vccd1 vccd1 _10329_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06385_ _06384_/A _06384_/B _06384_/X vssd1 vssd1 vccd1 vccd1 _06385_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ _08249_/A vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05336_ _05336_/A vssd1 vssd1 vccd1 vccd1 _05336_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05267_ _05093_/X _05263_/X _10352_/Q _05264_/X _05265_/X vssd1 vssd1 vccd1 vccd1
+ _10352_/D sky130_fd_sc_hd__a221o_1
X_08055_ _07023_/C _06824_/X _07385_/X _07400_/A vssd1 vssd1 vccd1 vccd1 _08055_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05198_ _05236_/A vssd1 vssd1 vccd1 vccd1 _05198_/X sky130_fd_sc_hd__clkbuf_2
X_07006_ _07056_/C vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08957_ _09938_/X vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__clkbuf_2
X_08888_ _09289_/A _09045_/B _09300_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _08891_/B
+ sky130_fd_sc_hd__o22a_1
X_07908_ _07783_/X _07785_/X _07783_/X _07785_/X vssd1 vssd1 vccd1 vccd1 _07915_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07839_ _07839_/A vssd1 vssd1 vccd1 vccd1 _07839_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09509_ _09508_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__mux2_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10215_ _10217_/CLK _10215_/D vssd1 vssd1 vccd1 vccd1 _10215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10146_ _10330_/CLK _10146_/D vssd1 vssd1 vccd1 vccd1 _10146_/Q sky130_fd_sc_hd__dfxtp_1
X_10077_ _10205_/CLK _10077_/D vssd1 vssd1 vccd1 vccd1 _10077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06170_ _06176_/A vssd1 vssd1 vccd1 vccd1 _06175_/A sky130_fd_sc_hd__buf_1
X_05121_ _10408_/Q vssd1 vssd1 vccd1 vccd1 _06614_/C sky130_fd_sc_hd__inv_2
XFILLER_144_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05052_ _05468_/A vssd1 vssd1 vccd1 vccd1 _05189_/A sky130_fd_sc_hd__clkbuf_4
X_09860_ _09859_/X _08290_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08811_ _08824_/A _08811_/B vssd1 vssd1 vccd1 vccd1 _08812_/B sky130_fd_sc_hd__and2b_1
X_09791_ _10356_/Q _09790_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09791_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08742_ _08742_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08742_/Y sky130_fd_sc_hd__nor2_1
X_05954_ _10223_/Q vssd1 vssd1 vccd1 vccd1 _07219_/A sky130_fd_sc_hd__clkbuf_2
X_08673_ _08172_/X _10061_/Q _08125_/X _10062_/Q vssd1 vssd1 vccd1 vccd1 _08673_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05885_ _05934_/A vssd1 vssd1 vccd1 vccd1 _05885_/X sky130_fd_sc_hd__clkbuf_4
X_07624_ _07597_/C _07593_/X _07597_/C _07593_/X vssd1 vssd1 vccd1 vccd1 _07625_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07555_ _07538_/X _07539_/X _07553_/X _07554_/X vssd1 vssd1 vccd1 vccd1 _07555_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06506_ _08411_/A _06496_/A _10093_/Q _06462_/A vssd1 vssd1 vccd1 vccd1 _06516_/C
+ sky130_fd_sc_hd__a22o_1
X_07486_ _10215_/Q vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__inv_2
X_06437_ _06437_/A vssd1 vssd1 vccd1 vccd1 _06489_/A sky130_fd_sc_hd__buf_1
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09225_ _09225_/A vssd1 vssd1 vccd1 vccd1 _09225_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09156_ _09107_/Y _09155_/X _09107_/Y _09155_/X vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06368_ _06362_/Y _06367_/A _06362_/A _06367_/Y vssd1 vssd1 vccd1 vccd1 _06368_/X
+ sky130_fd_sc_hd__o22a_1
X_08107_ _08804_/A vssd1 vssd1 vccd1 vccd1 _08107_/X sky130_fd_sc_hd__buf_2
X_09087_ _09087_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09187_/A sky130_fd_sc_hd__or2_1
X_05319_ _05319_/A vssd1 vssd1 vccd1 vccd1 _05320_/B sky130_fd_sc_hd__inv_2
X_06299_ _10238_/Q vssd1 vssd1 vccd1 vccd1 _06299_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _08023_/A _08023_/B _08024_/B vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10000_ _09999_/X _07802_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09989_ _08010_/A _08046_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10129_ _10447_/CLK _10129_/D vssd1 vssd1 vccd1 vccd1 _10129_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05670_ _05653_/X _05667_/Y _05668_/Y _08065_/A _05644_/X vssd1 vssd1 vccd1 vccd1
+ _05671_/B sky130_fd_sc_hd__o32a_1
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07340_ _07334_/X _07339_/X _07334_/X _07339_/X vssd1 vssd1 vccd1 vccd1 _07340_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_188_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09010_ _09097_/A _09010_/B _09010_/C vssd1 vssd1 vccd1 vccd1 _09010_/X sky130_fd_sc_hd__or3_1
X_07271_ _06866_/A _07102_/B _07068_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07271_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06222_ _09686_/X _06217_/X _10087_/Q _06218_/X vssd1 vssd1 vccd1 vccd1 _10087_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06153_ _09652_/X _06148_/X _10134_/Q _06149_/X _06146_/X vssd1 vssd1 vccd1 vccd1
+ _10134_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05104_ _06099_/A vssd1 vssd1 vccd1 vccd1 _05105_/A sky130_fd_sc_hd__buf_2
XFILLER_144_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06084_ _06084_/A vssd1 vssd1 vccd1 vccd1 _09943_/S sky130_fd_sc_hd__inv_2
X_05035_ _06119_/A vssd1 vssd1 vccd1 vccd1 _06176_/A sky130_fd_sc_hd__buf_2
X_09912_ _09911_/X _07897_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__mux2_1
X_09843_ _10369_/Q _09842_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _08199_/X _10352_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06986_ _07311_/A _07228_/A _06970_/A _06985_/A vssd1 vssd1 vccd1 vccd1 _06986_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08725_ _08722_/A _08724_/B _06631_/Y _08724_/Y vssd1 vssd1 vccd1 vccd1 _08726_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05937_ _09294_/A _05927_/X _05030_/X _05928_/X _05934_/X vssd1 vssd1 vccd1 vccd1
+ _10229_/D sky130_fd_sc_hd__o221a_1
X_08656_ _08155_/X _10050_/Q _10180_/Q _08467_/A vssd1 vssd1 vccd1 vccd1 _08656_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05868_ _05803_/X _05819_/X _05803_/X _05819_/X vssd1 vssd1 vccd1 vccd1 _05869_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08587_ _08587_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08595_/B sky130_fd_sc_hd__nand2_1
X_07607_ _07613_/B _09919_/X _07667_/A _07587_/D vssd1 vssd1 vccd1 vccd1 _07608_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05799_ _10274_/Q _10257_/Q _05797_/Y _05798_/Y vssd1 vssd1 vccd1 vccd1 _05799_/X
+ sky130_fd_sc_hd__a22o_1
X_07538_ _07538_/A _07537_/X vssd1 vssd1 vccd1 vccd1 _07538_/X sky130_fd_sc_hd__or2b_1
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07469_ _07660_/B vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__buf_1
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _09197_/X _09207_/X _09197_/X _09207_/X vssd1 vssd1 vccd1 vccd1 _09208_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ _09187_/B vssd1 vssd1 vccd1 vccd1 _09139_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_9_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10205_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06840_ _07164_/A vssd1 vssd1 vccd1 vccd1 _07146_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06771_ _10396_/Q _06802_/B _10397_/Q _06804_/B _06770_/X vssd1 vssd1 vccd1 vccd1
+ _06771_/X sky130_fd_sc_hd__a221o_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08510_ _10198_/Q _08504_/B _06263_/A _08509_/Y vssd1 vssd1 vccd1 vccd1 _08597_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09490_ _08435_/B _09583_/S _09600_/S vssd1 vssd1 vccd1 vccd1 _09490_/X sky130_fd_sc_hd__mux2_8
X_05722_ _10290_/Q _05715_/X _08850_/B _05719_/X _05711_/X vssd1 vssd1 vccd1 vccd1
+ _10290_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08441_ _08452_/B vssd1 vssd1 vccd1 vccd1 _08450_/B sky130_fd_sc_hd__clkbuf_2
X_05653_ _05718_/A vssd1 vssd1 vccd1 vccd1 _05653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08372_ _09625_/X _08391_/B vssd1 vssd1 vccd1 vccd1 _08372_/Y sky130_fd_sc_hd__nor2_1
X_05584_ _05695_/A _08899_/C vssd1 vssd1 vccd1 vccd1 _05694_/A sky130_fd_sc_hd__or2_1
XFILLER_176_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ _07321_/X _07322_/X _07321_/X _07322_/X vssd1 vssd1 vccd1 vccd1 _07323_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07254_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07254_/X sky130_fd_sc_hd__or2_1
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06205_ _09699_/X _06203_/X _10100_/Q _06204_/X vssd1 vssd1 vccd1 vccd1 _10100_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07185_ _07142_/X _07184_/X _07142_/X _07184_/X vssd1 vssd1 vccd1 vccd1 _07185_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06136_ _10143_/Q _05623_/X _10315_/Q _06130_/X _06135_/X vssd1 vssd1 vccd1 vccd1
+ _10143_/D sky130_fd_sc_hd__o221a_1
X_06067_ _06067_/A vssd1 vssd1 vccd1 vccd1 _06067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05018_ _10449_/Q vssd1 vssd1 vccd1 vccd1 _05018_/X sky130_fd_sc_hd__buf_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09826_ _08254_/Y _10365_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__mux2_1
X_09757_ _09756_/X input19/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06969_ _06977_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _06970_/A sky130_fd_sc_hd__or2_2
XFILLER_199_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08708_ _06690_/A _08709_/B _06625_/Y _08707_/Y vssd1 vssd1 vccd1 vccd1 _08708_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09688_ _06485_/Y input20/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08724_/B vssd1 vssd1 vccd1 vccd1 _08717_/B sky130_fd_sc_hd__buf_1
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10394_ _10426_/CLK _10394_/D vssd1 vssd1 vccd1 vccd1 _10394_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08990_ _08989_/A _08989_/B _09022_/A vssd1 vssd1 vccd1 vccd1 _08990_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _07937_/X _07938_/X _07937_/X _07938_/X vssd1 vssd1 vccd1 vccd1 _07941_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_205_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _07862_/X _07863_/X _07870_/X _07871_/X vssd1 vssd1 vccd1 vccd1 _07872_/X
+ sky130_fd_sc_hd__o22a_1
X_09611_ _10424_/Q _08074_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09611_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06823_ _06820_/A _06820_/B _06821_/B vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__a21bo_1
X_06754_ _10354_/Q vssd1 vssd1 vccd1 vccd1 _06755_/B sky130_fd_sc_hd__inv_2
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09542_ _10381_/Q _10178_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05705_ _05863_/A vssd1 vssd1 vccd1 vccd1 _05705_/X sky130_fd_sc_hd__clkbuf_2
X_06685_ _10373_/Q _08715_/A vssd1 vssd1 vccd1 vccd1 _08713_/A sky130_fd_sc_hd__or2_2
X_09473_ _09408_/A _09292_/B _09356_/B _09232_/Y _09355_/A vssd1 vssd1 vccd1 vccd1
+ _09473_/X sky130_fd_sc_hd__o32a_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08424_ _09533_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08424_/Y sky130_fd_sc_hd__nor2_1
X_05636_ _05718_/A vssd1 vssd1 vccd1 vccd1 _05863_/A sky130_fd_sc_hd__clkbuf_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05567_ _09987_/X _05566_/X _09987_/X _05566_/X vssd1 vssd1 vccd1 vccd1 _05668_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_08355_ _08355_/A _09748_/S vssd1 vssd1 vccd1 vccd1 _08355_/X sky130_fd_sc_hd__or2_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07306_ _07089_/A _07095_/A _07089_/Y vssd1 vssd1 vccd1 vccd1 _07306_/X sky130_fd_sc_hd__a21o_1
X_08286_ _08289_/B vssd1 vssd1 vccd1 vccd1 _08286_/Y sky130_fd_sc_hd__inv_2
X_05498_ _09988_/X _09996_/X _09988_/X _09996_/X vssd1 vssd1 vccd1 vccd1 _05498_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07237_ _07233_/X _07236_/X _07233_/X _07236_/X vssd1 vssd1 vccd1 vccd1 _07269_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07168_ _07154_/X _07155_/X _07154_/X _07155_/X vssd1 vssd1 vccd1 vccd1 _07168_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06119_ _06119_/A vssd1 vssd1 vccd1 vccd1 _06154_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07099_ _07099_/A vssd1 vssd1 vccd1 vccd1 _07099_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09809_ _09808_/X input23/X _09821_/S vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_2_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10178_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10274_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10446_ _10447_/CLK _10446_/D vssd1 vssd1 vccd1 vccd1 _10446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10377_ _10442_/CLK _10377_/D vssd1 vssd1 vccd1 vccd1 _10377_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06470_ _08385_/A _06487_/A _10087_/Q _06461_/A vssd1 vssd1 vccd1 vccd1 _06474_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05421_ _05421_/A vssd1 vssd1 vccd1 vccd1 _05422_/B sky130_fd_sc_hd__inv_2
X_08140_ _08504_/A vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__inv_2
XFILLER_14_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05352_ _10336_/Q _05352_/B vssd1 vssd1 vccd1 vccd1 _05352_/Y sky130_fd_sc_hd__nor2_1
X_05283_ _10345_/Q vssd1 vssd1 vccd1 vccd1 _05309_/A sky130_fd_sc_hd__inv_2
X_08071_ _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08071_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _06901_/X _06904_/X _06905_/X _06926_/X _06884_/X vssd1 vssd1 vccd1 vccd1
+ _07022_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_142_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08973_ _08972_/A _08995_/B _08972_/Y vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__a21oi_2
X_07924_ _07781_/Y _07923_/X _07781_/Y _07923_/X vssd1 vssd1 vccd1 vccd1 _07924_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07855_ _07855_/A vssd1 vssd1 vccd1 vccd1 _07878_/C sky130_fd_sc_hd__buf_2
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06806_ _06808_/A _06806_/B vssd1 vssd1 vccd1 vccd1 _06806_/Y sky130_fd_sc_hd__nor2_1
X_04998_ input51/X vssd1 vssd1 vccd1 vccd1 _06184_/A sky130_fd_sc_hd__inv_2
X_07786_ _07779_/X _07782_/Y _07783_/X _07785_/X vssd1 vssd1 vccd1 vccd1 _07786_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06737_ _08625_/A _08624_/B _06656_/Y vssd1 vssd1 vccd1 vccd1 _06737_/X sky130_fd_sc_hd__a21o_1
X_09525_ _09524_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09389_/X _09390_/X _09391_/X _09395_/Y _09343_/X vssd1 vssd1 vccd1 vccd1
+ _09456_/Y sky130_fd_sc_hd__o221ai_2
X_06668_ _10356_/Q _06668_/B vssd1 vssd1 vccd1 vccd1 _06669_/B sky130_fd_sc_hd__or2_1
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ _08407_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08407_/Y sky130_fd_sc_hd__nor2_1
X_05619_ _06130_/A vssd1 vssd1 vccd1 vccd1 _05619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06599_ _10382_/Q vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__inv_2
X_09387_ _09387_/A vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__inv_2
XFILLER_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ _09972_/X _08364_/B vssd1 vssd1 vccd1 vccd1 _08338_/Y sky130_fd_sc_hd__nor2_1
X_08269_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08273_/B sky130_fd_sc_hd__or2_1
XFILLER_165_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _10300_/CLK _10300_/D vssd1 vssd1 vccd1 vccd1 _10300_/Q sky130_fd_sc_hd__dfxtp_1
X_10231_ _10312_/CLK _10231_/D vssd1 vssd1 vccd1 vccd1 _10231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ _10334_/CLK _10162_/D vssd1 vssd1 vccd1 vccd1 _10162_/Q sky130_fd_sc_hd__dfxtp_1
X_10093_ _10176_/CLK _10093_/D vssd1 vssd1 vccd1 vccd1 _10093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10429_ _10433_/CLK _10429_/D vssd1 vssd1 vccd1 vccd1 _10429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05970_ _05970_/A vssd1 vssd1 vccd1 vccd1 _05970_/X sky130_fd_sc_hd__buf_1
XFILLER_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07640_ _07640_/A _07640_/B vssd1 vssd1 vccd1 vccd1 _07640_/X sky130_fd_sc_hd__or2_1
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07571_ _07571_/A vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__inv_2
XFILLER_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ _09310_/A _09417_/A vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__or2_2
X_06522_ _10096_/Q _06463_/A _08420_/A _06536_/A vssd1 vssd1 vccd1 vccd1 _06527_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06453_ _10085_/Q vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__inv_2
X_09241_ _09240_/A _09240_/B _09393_/A vssd1 vssd1 vccd1 vccd1 _09241_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _09292_/A _09354_/D vssd1 vssd1 vccd1 vccd1 _09294_/C sky130_fd_sc_hd__or2_2
X_06384_ _06384_/A _06384_/B vssd1 vssd1 vccd1 vccd1 _06384_/X sky130_fd_sc_hd__or2_1
X_05404_ _05404_/A vssd1 vssd1 vccd1 vccd1 _05404_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ _10193_/Q vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__inv_2
XFILLER_159_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05335_ _10340_/Q _05335_/B vssd1 vssd1 vccd1 vccd1 _05335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08054_ _08015_/A _08015_/B _08016_/B vssd1 vssd1 vccd1 vccd1 _08054_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05266_ _05091_/X _05263_/X _10353_/Q _05264_/X _05265_/X vssd1 vssd1 vccd1 vccd1
+ _10353_/D sky130_fd_sc_hd__a221o_1
X_07005_ _07235_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07056_/C sky130_fd_sc_hd__nor2_1
XFILLER_162_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05197_ _05468_/A vssd1 vssd1 vccd1 vccd1 _05236_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08956_ _08955_/A _08955_/B _08989_/A vssd1 vssd1 vccd1 vccd1 _08956_/X sky130_fd_sc_hd__a21bo_1
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08887_ _09010_/B vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__clkbuf_2
X_07907_ _07907_/A _07907_/B vssd1 vssd1 vccd1 vccd1 _07928_/A sky130_fd_sc_hd__or2_1
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07838_ _10213_/Q _07885_/B _07849_/A vssd1 vssd1 vccd1 vccd1 _07839_/A sky130_fd_sc_hd__and3_1
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09508_ _09507_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09508_/X sky130_fd_sc_hd__mux2_1
X_07769_ _07921_/B _07916_/C _07921_/A vssd1 vssd1 vccd1 vccd1 _07769_/X sky130_fd_sc_hd__or3_1
XFILLER_197_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09439_ _09338_/X _09381_/A _09380_/X vssd1 vssd1 vccd1 vccd1 _09439_/X sky130_fd_sc_hd__o21a_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10214_ _10217_/CLK _10214_/D vssd1 vssd1 vccd1 vccd1 _10214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ _10330_/CLK _10145_/D vssd1 vssd1 vccd1 vccd1 _10145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10076_ _10205_/CLK _10076_/D vssd1 vssd1 vccd1 vccd1 _10076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05120_ _05133_/A _05120_/B vssd1 vssd1 vccd1 vccd1 _10409_/D sky130_fd_sc_hd__nor2_1
XFILLER_129_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05051_ _10440_/Q _05047_/X input40/X _05048_/X _05036_/X vssd1 vssd1 vccd1 vccd1
+ _10440_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08810_ _08810_/A _08823_/A vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__or2_1
XFILLER_124_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09790_ _08214_/X _10356_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09790_/X sky130_fd_sc_hd__mux2_1
X_08741_ _08741_/A _08741_/B _08741_/C vssd1 vssd1 vccd1 vccd1 _08824_/C sky130_fd_sc_hd__or3_1
X_05953_ _07056_/A _05947_/X _05091_/X _05948_/X _05950_/X vssd1 vssd1 vccd1 vccd1
+ _10224_/D sky130_fd_sc_hd__o221a_1
X_08672_ _06030_/X _08671_/Y _06035_/X _08524_/Y vssd1 vssd1 vccd1 vccd1 _08674_/C
+ sky130_fd_sc_hd__a22o_1
X_05884_ _06119_/A vssd1 vssd1 vccd1 vccd1 _05934_/A sky130_fd_sc_hd__buf_2
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07623_ _07610_/A _07610_/B _07639_/A vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07554_ _07538_/X _07539_/X _07538_/X _07539_/X vssd1 vssd1 vccd1 vccd1 _07554_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06505_ _10093_/Q vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__inv_2
X_07485_ _07485_/A _07552_/B vssd1 vssd1 vccd1 vccd1 _07485_/X sky130_fd_sc_hd__or2_1
XFILLER_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06436_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06437_/A sky130_fd_sc_hd__buf_1
XFILLER_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _09213_/X _09214_/X _09159_/X _09215_/X vssd1 vssd1 vccd1 vccd1 _09224_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09155_ _09153_/X _09154_/X _09153_/X _09154_/X vssd1 vssd1 vccd1 vccd1 _09155_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06367_ _06367_/A vssd1 vssd1 vccd1 vccd1 _06367_/Y sky130_fd_sc_hd__inv_2
X_08106_ _08232_/A vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05318_ _05309_/B _05312_/B _05317_/X _06086_/A _10344_/Q vssd1 vssd1 vccd1 vccd1
+ _10344_/D sky130_fd_sc_hd__a32o_1
X_09086_ _09085_/A _09084_/Y _09085_/Y _09084_/A vssd1 vssd1 vccd1 vccd1 _09087_/B
+ sky130_fd_sc_hd__a22o_1
X_06298_ _06294_/X _06297_/X _06294_/X _06297_/X vssd1 vssd1 vccd1 vccd1 _06298_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05249_ _10359_/Q vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__buf_2
X_08037_ _07409_/A _07409_/B _07410_/B vssd1 vssd1 vccd1 vccd1 _08037_/X sky130_fd_sc_hd__a21bo_1
XFILLER_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _08001_/X _08056_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _09988_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08939_ _08939_/A _09977_/X _08939_/C vssd1 vssd1 vccd1 vccd1 _08939_/X sky130_fd_sc_hd__or3_1
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _10447_/CLK _10128_/D vssd1 vssd1 vccd1 vccd1 _10128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10059_ _10426_/CLK _10059_/D vssd1 vssd1 vccd1 vccd1 _10059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07270_ _07267_/X _07269_/X _07267_/X _07269_/X vssd1 vssd1 vccd1 vccd1 _07270_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06221_ _09687_/X _06217_/X _10088_/Q _06218_/X vssd1 vssd1 vccd1 vccd1 _10088_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06152_ _09653_/X _06148_/X _10135_/Q _06149_/X _06146_/X vssd1 vssd1 vccd1 vccd1
+ _10135_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05103_ _05038_/X _05047_/X _10411_/Q _05048_/X _05097_/X vssd1 vssd1 vccd1 vccd1
+ _10411_/D sky130_fd_sc_hd__a221o_1
X_06083_ _06083_/A _06240_/A vssd1 vssd1 vccd1 vccd1 _06084_/A sky130_fd_sc_hd__or2_1
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05034_ _05034_/A vssd1 vssd1 vccd1 vccd1 _06119_/A sky130_fd_sc_hd__clkbuf_2
X_09911_ _09910_/X _07031_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09911_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _08272_/Y _10369_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09773_ _09772_/X input45/X _09781_/S vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _08724_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08724_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06985_ _06985_/A vssd1 vssd1 vccd1 vccd1 _07228_/A sky130_fd_sc_hd__inv_2
X_05936_ _10229_/Q vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08655_ _08569_/A _10051_/Q _08121_/X _10052_/Q vssd1 vssd1 vccd1 vccd1 _08655_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05867_ _10257_/Q _05851_/X _05863_/X _06829_/A _05866_/X vssd1 vssd1 vccd1 vccd1
+ _10257_/D sky130_fd_sc_hd__o221a_1
X_08586_ _08586_/A _08586_/B _08586_/C vssd1 vssd1 vccd1 vccd1 _08602_/A sky130_fd_sc_hd__and3_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07606_ _07600_/X _07605_/X _07600_/X _07605_/X vssd1 vssd1 vccd1 vccd1 _07606_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07537_ _07828_/A _07552_/B _07830_/A _07537_/D vssd1 vssd1 vccd1 vccd1 _07537_/X
+ sky130_fd_sc_hd__or4_4
X_05798_ _10257_/Q vssd1 vssd1 vccd1 vccd1 _05798_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _10217_/Q vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__inv_2
X_09207_ _09319_/A _09207_/B vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__or2_1
X_06419_ _10079_/Q _06418_/X _10079_/Q _06418_/X vssd1 vssd1 vccd1 vccd1 _06419_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07399_ _06942_/A _06824_/X _07384_/B vssd1 vssd1 vccd1 vccd1 _07400_/A sky130_fd_sc_hd__o21ai_2
XFILLER_147_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _09136_/Y _09137_/Y _09136_/Y _09137_/Y vssd1 vssd1 vccd1 vccd1 _09187_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_162_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09069_/A _09976_/X vssd1 vssd1 vccd1 vccd1 _09122_/A sky130_fd_sc_hd__or2_2
XFILLER_190_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06770_ _10395_/Q _06801_/B _10396_/Q _06802_/B _06769_/X vssd1 vssd1 vccd1 vccd1
+ _06770_/X sky130_fd_sc_hd__o221a_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05721_ _10274_/Q vssd1 vssd1 vccd1 vccd1 _08850_/B sky130_fd_sc_hd__buf_2
X_08440_ _09967_/X _08449_/B vssd1 vssd1 vccd1 vccd1 _08440_/Y sky130_fd_sc_hd__nor2_1
X_05652_ _05677_/A _05652_/B vssd1 vssd1 vccd1 vccd1 _10308_/D sky130_fd_sc_hd__nor2_1
XFILLER_211_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08371_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08391_/B sky130_fd_sc_hd__buf_1
X_05583_ _08915_/A _08882_/A vssd1 vssd1 vccd1 vccd1 _08899_/C sky130_fd_sc_hd__or2_2
XFILLER_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07322_ _06958_/A _06958_/B _06958_/X vssd1 vssd1 vccd1 vccd1 _07322_/X sky130_fd_sc_hd__a21bo_1
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07253_ _07253_/A _07253_/B vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__nor2_1
XFILLER_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06204_ _06204_/A vssd1 vssd1 vccd1 vccd1 _06204_/X sky130_fd_sc_hd__clkbuf_2
X_07184_ _07158_/X _07161_/X _07162_/X _07183_/X _07144_/X vssd1 vssd1 vccd1 vccd1
+ _07184_/X sky130_fd_sc_hd__o221a_1
XFILLER_191_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06135_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06135_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06066_ _09785_/X _06054_/X _08545_/A _06056_/X _06057_/X vssd1 vssd1 vccd1 vccd1
+ _10183_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05017_ _05016_/A _05016_/B _05016_/Y vssd1 vssd1 vccd1 vccd1 _05017_/Y sky130_fd_sc_hd__a21oi_1
X_09825_ _09824_/X input27/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09756_ _09755_/X _08179_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09756_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06968_ _07217_/B vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__buf_1
X_08707_ _08707_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08707_/Y sky130_fd_sc_hd__nor2_1
X_09687_ _06479_/X input50/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__mux2_1
X_05919_ _10235_/Q _05910_/X _05101_/X _05911_/X _05918_/X vssd1 vssd1 vccd1 vccd1
+ _10235_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08638_ _08742_/B vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__clkbuf_2
X_06899_ _06888_/X _06889_/X _06897_/X _06898_/X vssd1 vssd1 vccd1 vccd1 _06899_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08569_/Y sky130_fd_sc_hd__nand2_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10393_ _10426_/CLK _10393_/D vssd1 vssd1 vccd1 vccd1 _10393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_190_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _07934_/X _07939_/X _07934_/X _07939_/X vssd1 vssd1 vccd1 vccd1 _07940_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _07862_/X _07863_/X _07862_/X _07863_/X vssd1 vssd1 vccd1 vccd1 _07871_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_205_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _10423_/Q _08073_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09610_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06822_ _06821_/A _06821_/B _06826_/B vssd1 vssd1 vccd1 vccd1 _06822_/X sky130_fd_sc_hd__a21bo_1
X_06753_ _06748_/Y _06790_/B _06752_/X vssd1 vssd1 vccd1 vccd1 _06753_/Y sky130_fd_sc_hd__a21oi_1
X_09541_ _09540_/X _10112_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__mux2_1
X_05704_ _08842_/B vssd1 vssd1 vccd1 vccd1 _05704_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06684_ _10372_/Q _08717_/A vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__or2_2
X_09472_ _09468_/Y _09471_/X _09468_/Y _09471_/X vssd1 vssd1 vccd1 vccd1 _09472_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08423_ _08423_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08423_/Y sky130_fd_sc_hd__nor2_1
X_05635_ _05646_/A _05635_/B vssd1 vssd1 vccd1 vccd1 _10311_/D sky130_fd_sc_hd__nor2_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08354_ _09354_/A vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05566_ _05490_/X _05520_/X _05490_/X _05520_/X vssd1 vssd1 vccd1 vccd1 _05566_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_07305_ _07252_/X _07255_/X _07256_/X _07304_/X vssd1 vssd1 vccd1 vccd1 _07308_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08285_ _08285_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08289_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_8_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05497_ _05497_/A _05497_/B vssd1 vssd1 vccd1 vccd1 _05497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07236_ _06991_/Y _07228_/B _07228_/B _07235_/X vssd1 vssd1 vccd1 vccd1 _07236_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_152_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07167_ _07161_/C _07166_/A _07160_/A _07166_/Y vssd1 vssd1 vccd1 vccd1 _07167_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06118_ _10154_/Q _06117_/X _10326_/Q _06113_/X _06111_/X vssd1 vssd1 vccd1 vccd1
+ _10154_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07098_ _07125_/A _09887_/X vssd1 vssd1 vccd1 vccd1 _07099_/A sky130_fd_sc_hd__or2_2
X_06049_ _10190_/Q vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09808_ _09807_/X _08234_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09808_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09739_ _06812_/Y _10404_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10070_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10445_ _10447_/CLK _10445_/D vssd1 vssd1 vccd1 vccd1 _10445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10376_ _10442_/CLK _10376_/D vssd1 vssd1 vccd1 vccd1 _10376_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05420_ _05420_/A vssd1 vssd1 vccd1 vccd1 _10326_/D sky130_fd_sc_hd__inv_2
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05351_ _05351_/A vssd1 vssd1 vccd1 vccd1 _05352_/B sky130_fd_sc_hd__inv_2
XFILLER_201_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05282_ _05333_/A vssd1 vssd1 vccd1 vccd1 _05282_/X sky130_fd_sc_hd__buf_2
X_08070_ _08070_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07021_ _07118_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _07021_/X sky130_fd_sc_hd__or2_2
XFILLER_154_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08972_ _08972_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07923_ _07886_/B _07922_/Y _07886_/B _07922_/Y vssd1 vssd1 vccd1 vccd1 _07923_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07854_ _07854_/A _07854_/B _10282_/Q _07854_/D vssd1 vssd1 vccd1 vccd1 _07854_/X
+ sky130_fd_sc_hd__and4_1
X_06805_ _06808_/A _06805_/B vssd1 vssd1 vccd1 vccd1 _06805_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07785_ _07785_/A vssd1 vssd1 vccd1 vccd1 _07785_/X sky130_fd_sc_hd__buf_1
X_06736_ _06662_/X _06735_/X _06662_/X _06735_/X vssd1 vssd1 vccd1 vccd1 _06736_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09524_ _09523_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__mux2_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09451_/Y _09454_/X _09451_/Y _09454_/X vssd1 vssd1 vccd1 vccd1 _09455_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06667_ _10355_/Q _06667_/B vssd1 vssd1 vccd1 vccd1 _06668_/B sky130_fd_sc_hd__or2_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _09513_/X _08414_/B vssd1 vssd1 vccd1 vccd1 _08406_/Y sky130_fd_sc_hd__nor2_1
X_05618_ _10314_/Q _05467_/X _05468_/X _05617_/X vssd1 vssd1 vccd1 vccd1 _10314_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06598_ _08445_/B vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__buf_2
XFILLER_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _08840_/X _08871_/X _08840_/X _08871_/X vssd1 vssd1 vccd1 vccd1 _09387_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05549_ _09901_/X _05548_/X _09901_/X _05548_/X vssd1 vssd1 vccd1 vccd1 _05549_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08337_ _08397_/A vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__buf_1
XFILLER_192_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08268_ _06030_/X _06263_/B _08267_/Y vssd1 vssd1 vccd1 vccd1 _08268_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07219_ _07219_/A _07219_/B _07293_/A vssd1 vssd1 vccd1 vccd1 _07220_/B sky130_fd_sc_hd__and3_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _06072_/X _06247_/B _08198_/Y vssd1 vssd1 vccd1 vccd1 _08199_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10230_ _10312_/CLK _10230_/D vssd1 vssd1 vccd1 vccd1 _10230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10161_ _10334_/CLK _10161_/D vssd1 vssd1 vccd1 vccd1 _10161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10092_ _10346_/CLK _10092_/D vssd1 vssd1 vccd1 vccd1 _10092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10428_ _10433_/CLK _10428_/D vssd1 vssd1 vccd1 vccd1 _10428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10359_ _10421_/CLK _10359_/D vssd1 vssd1 vccd1 vccd1 _10359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07570_ _07553_/X _07554_/X _07553_/X _07554_/X vssd1 vssd1 vccd1 vccd1 _07571_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06521_ _10096_/Q vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__inv_2
XFILLER_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09240_ _09240_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06452_ _06450_/X _06451_/Y _06450_/X _06451_/Y vssd1 vssd1 vccd1 vccd1 _06452_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09171_/A vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__buf_1
X_05403_ _05403_/A vssd1 vssd1 vccd1 vccd1 _10330_/D sky130_fd_sc_hd__inv_2
X_06383_ _06383_/A vssd1 vssd1 vccd1 vccd1 _06384_/B sky130_fd_sc_hd__inv_2
X_08122_ _10197_/Q vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__inv_2
X_05334_ _05334_/A vssd1 vssd1 vccd1 vccd1 _05335_/B sky130_fd_sc_hd__inv_2
XFILLER_174_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08053_ _07401_/A _07401_/B _07402_/B vssd1 vssd1 vccd1 vccd1 _08053_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05265_ _05274_/A vssd1 vssd1 vccd1 vccd1 _05265_/X sky130_fd_sc_hd__clkbuf_2
X_07004_ _07189_/A vssd1 vssd1 vccd1 vccd1 _07081_/B sky130_fd_sc_hd__clkbuf_2
X_05196_ _05193_/X _10388_/Q _05194_/X _09607_/X _05189_/X vssd1 vssd1 vccd1 vccd1
+ _10388_/D sky130_fd_sc_hd__o221a_1
XFILLER_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10442_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_130_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08955_ _08955_/A _08955_/B vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__or2_1
XFILLER_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07906_ _07906_/A _07906_/B vssd1 vssd1 vccd1 vccd1 _07907_/B sky130_fd_sc_hd__and2_1
X_08886_ _09968_/X vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07837_ _07837_/A _07837_/B vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_26_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10298_/CLK sky130_fd_sc_hd__clkbuf_16
X_07768_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__buf_1
X_06719_ _08738_/A vssd1 vssd1 vccd1 vccd1 _06719_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09507_ _09506_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _07699_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__nor2_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09436_/X _09437_/X _09436_/X _09437_/X vssd1 vssd1 vccd1 vccd1 _09438_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09369_ _09202_/A _09315_/A _09408_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__a211o_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10213_ _10297_/CLK _10213_/D vssd1 vssd1 vccd1 vccd1 _10213_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10144_ _10330_/CLK _10144_/D vssd1 vssd1 vccd1 vccd1 _10144_/Q sky130_fd_sc_hd__dfxtp_1
X_10075_ _10205_/CLK _10075_/D vssd1 vssd1 vccd1 vccd1 _10075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05050_ _10441_/Q _05047_/X input42/X _05048_/X _05036_/X vssd1 vssd1 vccd1 vccd1
+ _10441_/D sky130_fd_sc_hd__o221a_1
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08740_ _08521_/A _08739_/Y _08253_/X _08735_/X vssd1 vssd1 vccd1 vccd1 _08741_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05952_ _10224_/Q vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08671_ _10066_/Q vssd1 vssd1 vccd1 vccd1 _08671_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05883_ _05883_/A vssd1 vssd1 vccd1 vccd1 _06820_/A sky130_fd_sc_hd__inv_2
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _07622_/A vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__inv_2
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07553_ _07540_/X _07542_/X _07550_/X _07552_/X vssd1 vssd1 vccd1 vccd1 _07553_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06504_ _06516_/B _06503_/X _06516_/B _06503_/X vssd1 vssd1 vccd1 vccd1 _06504_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07484_ _07511_/A vssd1 vssd1 vccd1 vccd1 _07484_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06435_ _06435_/A vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09223_ _09222_/A _09222_/B _09280_/A vssd1 vssd1 vccd1 vccd1 _09223_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09154_ _09088_/X _09102_/X _09104_/A _09105_/A vssd1 vssd1 vccd1 vccd1 _09154_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08105_ _10189_/Q vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__inv_2
X_06366_ _10243_/Q _08386_/A _06352_/B _06357_/X vssd1 vssd1 vccd1 vccd1 _06367_/A
+ sky130_fd_sc_hd__o22a_1
X_05317_ _10344_/Q _05317_/B vssd1 vssd1 vccd1 vccd1 _05317_/X sky130_fd_sc_hd__or2_1
X_09085_ _09085_/A vssd1 vssd1 vccd1 vccd1 _09085_/Y sky130_fd_sc_hd__inv_2
X_06297_ _10236_/Q _08343_/A _06285_/A _06288_/A vssd1 vssd1 vccd1 vccd1 _06297_/X
+ sky130_fd_sc_hd__o22a_1
X_05248_ _10360_/Q _05263_/A input23/X _05264_/A _05245_/X vssd1 vssd1 vccd1 vccd1
+ _10360_/D sky130_fd_sc_hd__o221a_1
XFILLER_107_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08036_ _08024_/A _08024_/B _08025_/B vssd1 vssd1 vccd1 vccd1 _08036_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05179_ _05179_/A _05179_/B vssd1 vssd1 vccd1 vccd1 _10396_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09987_ _08986_/X _08984_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09987_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08938_ _08993_/C _08937_/A _09038_/C _08937_/Y vssd1 vssd1 vccd1 vccd1 _08938_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08869_ _10294_/Q _07437_/Y _08845_/Y _08868_/X vssd1 vssd1 vccd1 vccd1 _08869_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _10249_/CLK _10127_/D vssd1 vssd1 vccd1 vccd1 _10127_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10058_ _10426_/CLK _10058_/D vssd1 vssd1 vccd1 vccd1 _10058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06220_ _09688_/X _06217_/X _10089_/Q _06218_/X vssd1 vssd1 vccd1 vccd1 _10089_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06151_ _09654_/X _06148_/X _10136_/Q _06149_/X _06146_/X vssd1 vssd1 vccd1 vccd1
+ _10136_/D sky130_fd_sc_hd__o221a_1
X_06082_ _06183_/A _06082_/B _08324_/B vssd1 vssd1 vccd1 vccd1 _06240_/A sky130_fd_sc_hd__or3_4
X_05102_ _05101_/X _05094_/X _10412_/Q _05095_/X _05097_/X vssd1 vssd1 vccd1 vccd1
+ _10412_/D sky130_fd_sc_hd__a221o_1
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05033_ _10445_/Q _05012_/A _05032_/X _05013_/A _06182_/A vssd1 vssd1 vccd1 vccd1
+ _10445_/D sky130_fd_sc_hd__o221a_1
X_09910_ _09909_/X _09470_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09910_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09841_ _09840_/X input32/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09841_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09772_ _09771_/X _08197_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09772_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06984_ _06984_/A vssd1 vssd1 vccd1 vccd1 _06984_/X sky130_fd_sc_hd__buf_1
X_08723_ _06706_/Y _08722_/Y _08719_/Y vssd1 vssd1 vccd1 vccd1 _08723_/Y sky130_fd_sc_hd__o21bai_1
X_05935_ _05933_/X _05927_/X _05028_/X _05928_/X _05934_/X vssd1 vssd1 vccd1 vccd1
+ _10230_/D sky130_fd_sc_hd__o221a_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _06047_/X _08643_/Y _08644_/X _08653_/X vssd1 vssd1 vccd1 vccd1 _08654_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05866_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05866_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _08597_/C _08585_/B vssd1 vssd1 vccd1 vccd1 _08586_/C sky130_fd_sc_hd__or2_1
X_07605_ _07811_/C _07676_/B _07605_/C vssd1 vssd1 vccd1 vccd1 _07605_/X sky130_fd_sc_hd__or3_1
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05797_ _10274_/Q vssd1 vssd1 vccd1 vccd1 _05797_/Y sky130_fd_sc_hd__inv_2
X_07536_ _07811_/C vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__buf_2
X_09206_ _09310_/A _09259_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09207_/B sky130_fd_sc_hd__o21a_1
X_07467_ _07485_/A vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_194_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06418_ _10080_/Q _06420_/A _10080_/Q _06420_/A vssd1 vssd1 vccd1 vccd1 _06418_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_07398_ _07398_/A vssd1 vssd1 vccd1 vccd1 _07402_/A sky130_fd_sc_hd__inv_2
XFILLER_182_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09137_ _09073_/A _09075_/Y _09076_/X _09081_/X vssd1 vssd1 vccd1 vccd1 _09137_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_108_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06349_ _10243_/Q _08386_/A vssd1 vssd1 vccd1 vccd1 _06352_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _09067_/A _09067_/B _09117_/A vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__or2_1
XFILLER_150_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05720_ _10291_/Q _05715_/X _10275_/Q _05719_/X _05711_/X vssd1 vssd1 vccd1 vccd1
+ _10291_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05651_ _05619_/X _05648_/Y _05649_/Y _08070_/A _05644_/X vssd1 vssd1 vccd1 vccd1
+ _05652_/B sky130_fd_sc_hd__o32a_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _08370_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08370_/X sky130_fd_sc_hd__or2_1
XFILLER_211_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05582_ _05581_/X _05510_/A _10283_/Q _05510_/A vssd1 vssd1 vccd1 vccd1 _08882_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_07321_ _07049_/X _07050_/Y _07049_/X _07050_/Y vssd1 vssd1 vccd1 vccd1 _07321_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07252_ _07208_/X _07249_/X _07250_/X _07251_/X vssd1 vssd1 vccd1 vccd1 _07252_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06203_ _06203_/A vssd1 vssd1 vccd1 vccd1 _06203_/X sky130_fd_sc_hd__clkbuf_2
X_07183_ _07181_/A _07178_/X _07180_/X _07182_/Y vssd1 vssd1 vccd1 vccd1 _07183_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06134_ _10144_/Q _05623_/X _10316_/Q _06130_/X _06128_/X vssd1 vssd1 vccd1 vccd1
+ _10144_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06065_ _08772_/A vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__clkbuf_2
X_05016_ _05016_/A _05016_/B vssd1 vssd1 vccd1 vccd1 _05016_/Y sky130_fd_sc_hd__nor2_1
X_09824_ _09823_/X _08251_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09824_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _10347_/Q _09754_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06967_ _09885_/X vssd1 vssd1 vccd1 vccd1 _07217_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08706_ _08696_/X _08700_/X _08705_/X vssd1 vssd1 vccd1 vccd1 _08706_/Y sky130_fd_sc_hd__o21ai_2
X_09686_ _06475_/Y input49/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05918_ _05934_/A vssd1 vssd1 vccd1 vccd1 _05918_/X sky130_fd_sc_hd__buf_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06898_ _06942_/C _07031_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06898_/X sky130_fd_sc_hd__or3_1
X_08637_ _08738_/B vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__clkbuf_2
X_05849_ _05849_/A vssd1 vssd1 vccd1 vccd1 _06837_/A sky130_fd_sc_hd__inv_2
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08564_/Y _08589_/B _08589_/A vssd1 vssd1 vccd1 vccd1 _08568_/X sky130_fd_sc_hd__o21ba_1
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08499_ _10071_/Q _08489_/B _08490_/B vssd1 vssd1 vccd1 vccd1 _08499_/X sky130_fd_sc_hd__a21bo_1
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07519_ _07514_/X _07518_/X _07514_/X _07518_/X vssd1 vssd1 vccd1 vccd1 _07707_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10392_ _10426_/CLK _10392_/D vssd1 vssd1 vccd1 vccd1 _10392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07870_ _07869_/A _07869_/B _07869_/Y vssd1 vssd1 vccd1 vccd1 _07870_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06821_ _06821_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06826_/B sky130_fd_sc_hd__or2_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06752_ _06750_/Y _06789_/B _06733_/Y _06788_/B vssd1 vssd1 vccd1 vccd1 _06752_/X
+ sky130_fd_sc_hd__a22o_1
X_09540_ _10080_/Q _10040_/Q _09544_/S vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__mux2_1
X_09471_ _09469_/Y _09470_/Y _09469_/Y _09470_/Y vssd1 vssd1 vccd1 vccd1 _09471_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05703_ _10280_/Q vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__clkbuf_2
X_06683_ _10371_/Q _08719_/A vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__or2_1
X_08422_ _09531_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05634_ _05619_/X _05631_/Y _05632_/X _08073_/A _05623_/X vssd1 vssd1 vccd1 vccd1
+ _05635_/B sky130_fd_sc_hd__o32a_1
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ _09070_/A vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__clkbuf_2
X_05565_ _09946_/X _05564_/X _09946_/X _05564_/X vssd1 vssd1 vccd1 vccd1 _05663_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08284_ _06020_/X _06267_/B _08283_/Y vssd1 vssd1 vccd1 vccd1 _08284_/X sky130_fd_sc_hd__a21o_1
X_07304_ _07263_/X _07302_/X _07337_/B vssd1 vssd1 vccd1 vccd1 _07304_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07235_ _07235_/A _07235_/B _07245_/A vssd1 vssd1 vccd1 vccd1 _07235_/X sky130_fd_sc_hd__or3_2
X_05496_ _10001_/X vssd1 vssd1 vccd1 vccd1 _05497_/B sky130_fd_sc_hd__inv_2
XFILLER_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07166_ _07166_/A vssd1 vssd1 vccd1 vccd1 _07166_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06117_ _06126_/A vssd1 vssd1 vccd1 vccd1 _06117_/X sky130_fd_sc_hd__clkbuf_2
X_07097_ _07075_/X _07096_/X _07075_/X _07096_/X vssd1 vssd1 vccd1 vccd1 _07309_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06048_ _09817_/X _06043_/X _06047_/X _06044_/X _06045_/X vssd1 vssd1 vccd1 vccd1
+ _10191_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09807_ _10360_/Q _09806_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07999_ _07878_/A _07777_/B _07425_/A _07878_/C vssd1 vssd1 vccd1 vccd1 _08000_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09738_ _06811_/Y _10403_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10069_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09669_ _10150_/Q _10166_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10444_ _10447_/CLK _10444_/D vssd1 vssd1 vccd1 vccd1 _10444_/Q sky130_fd_sc_hd__dfxtp_1
X_10375_ _10442_/CLK _10375_/D vssd1 vssd1 vccd1 vccd1 _10375_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05350_ _05350_/A vssd1 vssd1 vccd1 vccd1 _10337_/D sky130_fd_sc_hd__inv_2
XFILLER_186_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05281_ _05311_/A vssd1 vssd1 vccd1 vccd1 _05333_/A sky130_fd_sc_hd__clkbuf_2
X_07020_ _07017_/Y _07019_/Y _07017_/Y _07019_/Y vssd1 vssd1 vccd1 vccd1 _07020_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_161_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08971_ _09038_/C _08937_/Y _08938_/X _08940_/X vssd1 vssd1 vccd1 vccd1 _08995_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_142_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07922_ _07920_/Y _07921_/Y _07769_/X vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__o21ai_2
X_07853_ _07827_/X _07830_/X _07831_/X _07852_/X _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07853_/Y sky130_fd_sc_hd__o221ai_2
X_06804_ _06808_/A _06804_/B vssd1 vssd1 vccd1 vccd1 _06804_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07784_ _07921_/B _07916_/A _07910_/C vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__mux2_1
X_06735_ _08624_/A _10351_/Q _06652_/Y vssd1 vssd1 vccd1 vccd1 _06735_/X sky130_fd_sc_hd__a21o_1
X_09523_ _09522_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09523_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ _09452_/X _09453_/X _09452_/X _09453_/X vssd1 vssd1 vccd1 vccd1 _09454_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06666_ _10354_/Q _06666_/B vssd1 vssd1 vccd1 vccd1 _06667_/B sky130_fd_sc_hd__or2_2
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _09384_/A _09384_/B _09442_/A vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__a21bo_1
X_05617_ _05615_/A _05614_/Y _10007_/S _05614_/A _05771_/A vssd1 vssd1 vccd1 vccd1
+ _05617_/X sky130_fd_sc_hd__a221o_1
X_08405_ _08405_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__or2_1
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06597_ _06466_/X _06596_/X _06466_/X _06596_/X vssd1 vssd1 vccd1 vccd1 _06597_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08336_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__inv_2
XFILLER_177_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05548_ _05546_/Y _05547_/Y _05546_/Y _05547_/Y vssd1 vssd1 vccd1 vccd1 _05548_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08267_ _08267_/A vssd1 vssd1 vccd1 vccd1 _08267_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05479_ _10019_/X vssd1 vssd1 vccd1 vccd1 _05481_/A sky130_fd_sc_hd__inv_2
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08198_ _08198_/A vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__inv_2
X_07218_ _07218_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _07293_/A sky130_fd_sc_hd__or2_1
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07149_ _07147_/X _07148_/X _07147_/X _07148_/X vssd1 vssd1 vccd1 vccd1 _07154_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10346_/CLK _10160_/D vssd1 vssd1 vccd1 vccd1 _10160_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10091_ _10346_/CLK _10091_/D vssd1 vssd1 vccd1 vccd1 _10091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10427_ _10433_/CLK _10427_/D vssd1 vssd1 vccd1 vccd1 _10427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10358_ _10421_/CLK _10358_/D vssd1 vssd1 vccd1 vccd1 _10358_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10289_ _10289_/CLK _10289_/D vssd1 vssd1 vccd1 vccd1 _10289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10102_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06520_ _06519_/A _06519_/B _06527_/A vssd1 vssd1 vccd1 vccd1 _06520_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06451_ _08357_/A _06438_/X _06447_/X vssd1 vssd1 vccd1 vccd1 _06451_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_194_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05402_ _10330_/Q _05372_/X _05400_/C _05397_/Y _05401_/Y vssd1 vssd1 vccd1 vccd1
+ _05403_/A sky130_fd_sc_hd__o32a_1
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _09170_/A _09225_/A _09170_/C vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__nand3_1
X_06382_ _06353_/Y _06362_/A _06372_/A _06345_/Y _06381_/X vssd1 vssd1 vccd1 vccd1
+ _06383_/A sky130_fd_sc_hd__a41o_1
X_08121_ _08208_/A vssd1 vssd1 vccd1 vccd1 _08121_/X sky130_fd_sc_hd__buf_2
X_05333_ _05333_/A vssd1 vssd1 vccd1 vccd1 _05333_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05264_ _05264_/A vssd1 vssd1 vccd1 vccd1 _05264_/X sky130_fd_sc_hd__clkbuf_2
X_08052_ _08016_/A _08016_/B _08017_/B vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__a21bo_1
X_07003_ _09890_/X vssd1 vssd1 vccd1 vccd1 _07189_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05195_ _05193_/X _10389_/Q _05194_/X _09608_/X _05189_/X vssd1 vssd1 vccd1 vccd1
+ _10389_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ _08955_/B vssd1 vssd1 vccd1 vccd1 _08954_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07905_ _07906_/A _07906_/B vssd1 vssd1 vccd1 vccd1 _07907_/A sky130_fd_sc_hd__nor2_1
X_08885_ _09069_/A vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07836_ _07823_/X _07824_/X _07823_/X _07824_/X vssd1 vssd1 vccd1 vccd1 _07836_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07767_ _07777_/C _07764_/X _07916_/B vssd1 vssd1 vccd1 vccd1 _07767_/X sky130_fd_sc_hd__mux2_1
X_06718_ _06718_/A vssd1 vssd1 vccd1 vccd1 _06805_/B sky130_fd_sc_hd__inv_2
X_09506_ _08383_/X _06337_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ _07698_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _07699_/B sky130_fd_sc_hd__or2_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09437_ _09360_/X _09361_/X _09362_/X _09376_/X vssd1 vssd1 vccd1 vccd1 _09437_/X
+ sky130_fd_sc_hd__o22a_1
X_06649_ _10351_/Q vssd1 vssd1 vccd1 vccd1 _08632_/A sky130_fd_sc_hd__inv_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _09260_/A _09367_/A _09261_/B _09367_/Y vssd1 vssd1 vccd1 vccd1 _09368_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09299_ _09945_/X vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__clkbuf_2
X_08319_ _08319_/A vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _10217_/CLK _10212_/D vssd1 vssd1 vccd1 vccd1 _10212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _10330_/CLK _10143_/D vssd1 vssd1 vccd1 vccd1 _10143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10074_ _10205_/CLK _10074_/D vssd1 vssd1 vccd1 vccd1 _10074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05951_ _05943_/X _05947_/X _05089_/X _05948_/X _05950_/X vssd1 vssd1 vccd1 vccd1
+ _10225_/D sky130_fd_sc_hd__o221a_1
X_08670_ _08253_/X _10063_/Q _08125_/X _10062_/Q vssd1 vssd1 vccd1 vccd1 _08674_/B
+ sky130_fd_sc_hd__a22o_1
X_05882_ _05815_/A _05881_/Y _05815_/A _05881_/Y vssd1 vssd1 vccd1 vccd1 _05883_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07621_ _07621_/A _07627_/A vssd1 vssd1 vccd1 vccd1 _07621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07552_ _07855_/A _07552_/B _07552_/C vssd1 vssd1 vccd1 vccd1 _07552_/X sky130_fd_sc_hd__or3_1
X_06503_ _10091_/Q _06466_/X _06494_/A _06499_/A vssd1 vssd1 vccd1 vccd1 _06503_/X
+ sky130_fd_sc_hd__a22o_1
X_07483_ _07483_/A _07566_/B _07509_/A vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__and3_1
XFILLER_166_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06434_ _06434_/A vssd1 vssd1 vccd1 vccd1 _06435_/A sky130_fd_sc_hd__clkbuf_2
X_09222_ _09222_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09153_ _09131_/X _09152_/X _09131_/X _09152_/X vssd1 vssd1 vccd1 vccd1 _09153_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06365_ _06362_/Y _06364_/A _06362_/A _06364_/Y vssd1 vssd1 vccd1 vccd1 _06365_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08104_ _08539_/A vssd1 vssd1 vccd1 vccd1 _08104_/X sky130_fd_sc_hd__clkbuf_2
X_05316_ _05309_/A _05313_/X _05309_/B _05313_/B vssd1 vssd1 vccd1 vccd1 _10345_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_174_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09084_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09084_/Y sky130_fd_sc_hd__inv_2
X_06296_ _06294_/X _06295_/Y _06294_/X _06295_/Y vssd1 vssd1 vccd1 vccd1 _06296_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05247_ _10361_/Q _05239_/X input24/X _05240_/X _05245_/X vssd1 vssd1 vccd1 vccd1
+ _10361_/D sky130_fd_sc_hd__o221a_1
X_08035_ _07410_/A _07410_/B _07411_/B vssd1 vssd1 vccd1 vccd1 _08035_/X sky130_fd_sc_hd__a21bo_1
X_05178_ _05193_/A _05176_/Y _05177_/Y _05161_/X vssd1 vssd1 vccd1 vccd1 _05179_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09986_ _08931_/X _08929_/A _09986_/S vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08937_ _08937_/A vssd1 vssd1 vccd1 vccd1 _08937_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08868_ _10293_/Q _05852_/X _08846_/X _08867_/X vssd1 vssd1 vccd1 vccd1 _08868_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _07819_/A _09916_/X vssd1 vssd1 vccd1 vccd1 _07820_/C sky130_fd_sc_hd__or2_2
X_08799_ _08086_/X _08774_/B _08215_/A _08767_/X vssd1 vssd1 vccd1 vccd1 _08820_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _10244_/CLK _10126_/D vssd1 vssd1 vccd1 vccd1 _10126_/Q sky130_fd_sc_hd__dfxtp_1
X_10057_ _10426_/CLK _10057_/D vssd1 vssd1 vccd1 vccd1 _10057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10437_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06150_ _09655_/X _06148_/X _10137_/Q _06149_/X _06146_/X vssd1 vssd1 vccd1 vccd1
+ _10137_/D sky130_fd_sc_hd__o221a_1
XFILLER_129_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05101_ input30/X vssd1 vssd1 vccd1 vccd1 _05101_/X sky130_fd_sc_hd__buf_4
X_06081_ _06081_/A _06081_/B input16/X vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__or3b_4
Xclkbuf_leaf_25_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10217_/CLK sky130_fd_sc_hd__clkbuf_16
X_05032_ input41/X vssd1 vssd1 vccd1 vccd1 _05032_/X sky130_fd_sc_hd__buf_2
XFILLER_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09840_ _09839_/X _08271_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09771_ _10351_/Q _09770_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06983_ _07213_/A _07047_/D _06976_/A vssd1 vssd1 vccd1 vccd1 _06984_/A sky130_fd_sc_hd__o21ai_1
X_08722_ _08722_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08722_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05934_ _05934_/A vssd1 vssd1 vccd1 vccd1 _05934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08653_ _08666_/A _08651_/Y _08652_/Y vssd1 vssd1 vccd1 vccd1 _08653_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05865_ _05865_/A vssd1 vssd1 vccd1 vccd1 _06829_/A sky130_fd_sc_hd__inv_2
XFILLER_54_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08584_ _08523_/X _08596_/A _08583_/X vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__o21ba_1
X_07604_ _07604_/A vssd1 vssd1 vccd1 vccd1 _07605_/C sky130_fd_sc_hd__inv_2
X_05796_ _10275_/Q _10258_/Q _07445_/A _05795_/Y vssd1 vssd1 vccd1 vccd1 _05796_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07535_ _07811_/A _07552_/B _07811_/C _07537_/D vssd1 vssd1 vccd1 vccd1 _07538_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07466_ _07663_/A vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__buf_1
X_06417_ _06233_/Y _10039_/Q _10036_/D _06236_/Y vssd1 vssd1 vccd1 vccd1 _06420_/A
+ sky130_fd_sc_hd__o22a_1
X_09205_ _09452_/A _09282_/A _09205_/C vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__nor3_4
XFILLER_139_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _07397_/A vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__inv_2
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09136_ _09134_/X _09135_/X _09134_/X _09135_/X vssd1 vssd1 vccd1 vccd1 _09136_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
X_06348_ _10136_/Q vssd1 vssd1 vccd1 vccd1 _08386_/A sky130_fd_sc_hd__inv_2
XFILLER_147_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ _09067_/A _09067_/B vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__or2_1
X_06279_ _05770_/A _10127_/Q _06277_/A _05771_/C _06277_/Y vssd1 vssd1 vccd1 vccd1
+ _06279_/X sky130_fd_sc_hd__o32a_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08018_ _08018_/A _08018_/B vssd1 vssd1 vccd1 vccd1 _08019_/B sky130_fd_sc_hd__or2_1
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09969_ _08335_/X _06275_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09969_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10109_ _10205_/CLK _10109_/D vssd1 vssd1 vccd1 vccd1 _10109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05650_ _10308_/Q vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__inv_2
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05581_ _10283_/Q vssd1 vssd1 vccd1 vccd1 _05581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07320_ _07316_/X _07319_/X _07316_/X _07319_/X vssd1 vssd1 vccd1 vccd1 _07320_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07251_ _07208_/X _07249_/X _07208_/X _07249_/X vssd1 vssd1 vccd1 vccd1 _07251_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06202_ _09700_/X _06196_/X _10101_/Q _06197_/X vssd1 vssd1 vccd1 vccd1 _10101_/D
+ sky130_fd_sc_hd__a22o_1
X_07182_ _07182_/A _07182_/B vssd1 vssd1 vccd1 vccd1 _07182_/Y sky130_fd_sc_hd__nor2_1
X_06133_ _10145_/Q _06126_/X _10317_/Q _06130_/X _06128_/X vssd1 vssd1 vccd1 vccd1
+ _10145_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06064_ _10183_/Q vssd1 vssd1 vccd1 vccd1 _08772_/A sky130_fd_sc_hd__clkbuf_2
X_05015_ input46/X vssd1 vssd1 vccd1 vccd1 _05016_/B sky130_fd_sc_hd__inv_2
X_09823_ _10364_/Q _09822_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _08077_/X _10347_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09754_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06966_ _10225_/Q vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__inv_2
XFILLER_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08705_ _08705_/A _08705_/B _08705_/C _08705_/D vssd1 vssd1 vccd1 vccd1 _08705_/X
+ sky130_fd_sc_hd__or4_4
X_09685_ _06468_/X input48/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__mux2_1
X_05917_ _05032_/X _05896_/X _10236_/Q _05897_/X _05274_/X vssd1 vssd1 vccd1 vccd1
+ _10236_/D sky130_fd_sc_hd__a221o_1
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06897_ _06897_/A _06897_/B vssd1 vssd1 vccd1 vccd1 _06897_/X sky130_fd_sc_hd__or2_1
XFILLER_54_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08636_ _08738_/B vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05848_ _05826_/A _05847_/Y _05826_/A _05847_/Y vssd1 vssd1 vccd1 vccd1 _05849_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08155_/X _08549_/X _08782_/A _08565_/Y vssd1 vssd1 vccd1 vccd1 _08589_/A
+ sky130_fd_sc_hd__a22o_1
X_05779_ _06083_/A _05777_/A input19/X _05468_/X _05778_/X vssd1 vssd1 vccd1 vccd1
+ _10266_/D sky130_fd_sc_hd__o311a_1
XFILLER_210_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08498_ _10072_/Q _08490_/B _08491_/B vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__a21bo_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07518_ _07506_/B _07517_/A _07505_/A _07517_/Y vssd1 vssd1 vccd1 vccd1 _07518_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _07613_/B vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09119_ _09045_/B _09042_/B _09168_/A _09043_/Y _08377_/A vssd1 vssd1 vccd1 vccd1
+ _09119_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10391_ _10426_/CLK _10391_/D vssd1 vssd1 vccd1 vccd1 _10391_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_190_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06820_ _06820_/A _06820_/B vssd1 vssd1 vccd1 vccd1 _06821_/B sky130_fd_sc_hd__or2_1
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06751_ _10353_/Q _06665_/B _06666_/B vssd1 vssd1 vccd1 vccd1 _06789_/B sky130_fd_sc_hd__a21bo_1
X_06682_ _10370_/Q _08722_/A vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__or2_2
X_09470_ _09470_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05702_ _10297_/Q _05701_/X _10281_/Q _05699_/X _05660_/X vssd1 vssd1 vccd1 vccd1
+ _10297_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08421_ _08453_/B vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__buf_1
XFILLER_91_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05633_ _10311_/Q vssd1 vssd1 vccd1 vccd1 _08073_/A sky130_fd_sc_hd__inv_2
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08352_ _10230_/Q vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__inv_2
X_05564_ _05562_/Y _05563_/Y _05562_/Y _05563_/Y vssd1 vssd1 vccd1 vccd1 _05564_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_08283_ _08283_/A vssd1 vssd1 vccd1 vccd1 _08283_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07303_ _07303_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__or2_1
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05495_ _10002_/X vssd1 vssd1 vccd1 vccd1 _05497_/A sky130_fd_sc_hd__inv_2
XFILLER_137_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07234_ _07234_/A _07234_/B vssd1 vssd1 vccd1 vccd1 _07245_/A sky130_fd_sc_hd__nor2_2
XFILLER_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07165_ _07165_/A _07219_/B _07176_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__and3_1
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06116_ _10155_/Q _05891_/X _10327_/Q _06113_/X _06111_/X vssd1 vssd1 vccd1 vccd1
+ _10155_/D sky130_fd_sc_hd__o221a_1
X_07096_ _07090_/A _07254_/A _07089_/Y _07087_/A _07095_/Y vssd1 vssd1 vccd1 vccd1
+ _07096_/X sky130_fd_sc_hd__o32a_1
X_06047_ _10191_/Q vssd1 vssd1 vccd1 vccd1 _06047_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09806_ _08231_/X _10360_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07998_ _07625_/A _07625_/B _07626_/B vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__a21bo_1
X_09737_ _06810_/Y _10402_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10068_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06949_ _07031_/A _06960_/B _07028_/A _06949_/D vssd1 vssd1 vccd1 vccd1 _06949_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ _06850_/X _05861_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__mux2_1
X_09599_ _08451_/Y _08450_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09599_/X sky130_fd_sc_hd__mux2_2
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08619_ _08623_/A _09944_/X vssd1 vssd1 vccd1 vccd1 _10041_/D sky130_fd_sc_hd__or2_1
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10443_ _10447_/CLK _10443_/D vssd1 vssd1 vccd1 vccd1 _10443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10374_ _10437_/CLK _10374_/D vssd1 vssd1 vccd1 vccd1 _10374_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05280_ _06086_/A _06185_/A vssd1 vssd1 vccd1 vccd1 _05311_/A sky130_fd_sc_hd__or2_1
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _08970_/A vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__inv_2
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07921_ _07921_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07852_ _07846_/A _07882_/A _07845_/Y _07843_/A _07851_/Y vssd1 vssd1 vccd1 vccd1
+ _07852_/X sky130_fd_sc_hd__o32a_1
Xinput1 io_QEI_ChA vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_06803_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06808_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07783_ _07779_/X _07782_/Y _07779_/X _07782_/Y vssd1 vssd1 vccd1 vccd1 _07783_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09522_ _08386_/X _06351_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__mux2_1
X_06734_ _06664_/A _06664_/B _06665_/B vssd1 vssd1 vccd1 vccd1 _06788_/B sky130_fd_sc_hd__o21ai_2
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09453_ _09411_/X _09412_/X _09359_/X _09413_/X vssd1 vssd1 vccd1 vccd1 _09453_/X
+ sky130_fd_sc_hd__o22a_1
X_06665_ _10353_/Q _06665_/B vssd1 vssd1 vccd1 vccd1 _06666_/B sky130_fd_sc_hd__or2_1
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09384_ _09384_/A _09384_/B vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__or2_1
X_08404_ _09615_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08404_/Y sky130_fd_sc_hd__nor2_2
X_05616_ _05718_/A vssd1 vssd1 vccd1 vccd1 _05771_/A sky130_fd_sc_hd__buf_1
X_06596_ _08452_/A _06595_/X _08452_/A _06595_/X vssd1 vssd1 vccd1 vccd1 _06596_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08335_ _08335_/A _09748_/S vssd1 vssd1 vccd1 vccd1 _08335_/X sky130_fd_sc_hd__or2_1
X_05547_ _05478_/A _05478_/B _05478_/Y vssd1 vssd1 vccd1 vccd1 _05547_/Y sky130_fd_sc_hd__a21oi_2
X_08266_ _06035_/X _08261_/Y _08264_/X _08269_/B vssd1 vssd1 vccd1 vccd1 _08266_/X
+ sky130_fd_sc_hd__o211a_1
X_05478_ _05478_/A _05478_/B vssd1 vssd1 vccd1 vccd1 _05478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08197_ _10180_/Q _08192_/Y _08200_/B _08188_/X vssd1 vssd1 vccd1 vccd1 _08197_/X
+ sky130_fd_sc_hd__o211a_1
X_07217_ _07218_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07223_/C sky130_fd_sc_hd__nor2_1
XFILLER_192_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07148_ _07155_/A _09885_/X vssd1 vssd1 vccd1 vccd1 _07148_/X sky130_fd_sc_hd__or2_1
XFILLER_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ _07079_/A _07079_/B vssd1 vssd1 vccd1 vccd1 _07090_/A sky130_fd_sc_hd__or2_1
XINSDIODE3_0 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10090_ _10346_/CLK _10090_/D vssd1 vssd1 vccd1 vccd1 _10090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10426_ _10426_/CLK _10426_/D vssd1 vssd1 vccd1 vccd1 _10426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10357_ _10421_/CLK _10357_/D vssd1 vssd1 vccd1 vccd1 _10357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10288_ _10289_/CLK _10288_/D vssd1 vssd1 vccd1 vccd1 _10288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06450_ _10084_/Q _06460_/A _08365_/A _06430_/A vssd1 vssd1 vccd1 vccd1 _06450_/X
+ sky130_fd_sc_hd__a22o_1
X_05401_ _09897_/X _06130_/A _05400_/X vssd1 vssd1 vccd1 vccd1 _05401_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_194_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06381_ _10245_/Q _08396_/A _06370_/Y _06375_/X vssd1 vssd1 vccd1 vccd1 _06381_/X
+ sky130_fd_sc_hd__o22a_1
X_08120_ _10183_/Q vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__inv_2
XFILLER_119_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05332_ _05332_/A vssd1 vssd1 vccd1 vccd1 _10341_/D sky130_fd_sc_hd__inv_2
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05263_ _05263_/A vssd1 vssd1 vccd1 vccd1 _05263_/X sky130_fd_sc_hd__clkbuf_2
X_08051_ _07402_/A _07402_/B _07403_/B vssd1 vssd1 vccd1 vccd1 _08051_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07002_ _07126_/B vssd1 vssd1 vccd1 vccd1 _07082_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05194_ _05203_/A vssd1 vssd1 vccd1 vccd1 _05194_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ _08862_/Y _08952_/X _08862_/Y _08952_/X vssd1 vssd1 vccd1 vccd1 _08955_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07904_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07906_/B sky130_fd_sc_hd__and2_1
X_08884_ _08915_/A vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__buf_1
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ _07835_/A _07835_/B vssd1 vssd1 vccd1 vccd1 _07846_/A sky130_fd_sc_hd__or2_1
X_07766_ _07766_/A _07777_/B _07770_/A vssd1 vssd1 vccd1 vccd1 _07916_/B sky130_fd_sc_hd__or3_4
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06717_ _10365_/Q _08734_/A _06715_/Y vssd1 vssd1 vccd1 vccd1 _06804_/B sky130_fd_sc_hd__a21oi_2
X_09505_ _09504_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09505_/X sky130_fd_sc_hd__mux2_1
X_09436_ _09426_/X _09435_/X _09426_/X _09435_/X vssd1 vssd1 vccd1 vccd1 _09436_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07697_ _07672_/C _07669_/B _07669_/Y vssd1 vssd1 vccd1 vccd1 _07698_/B sky130_fd_sc_hd__o21ai_1
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06648_ _10352_/Q vssd1 vssd1 vccd1 vccd1 _06664_/A sky130_fd_sc_hd__inv_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06579_ _10107_/Q _06466_/A _08446_/A _06437_/A vssd1 vssd1 vccd1 vccd1 _06583_/A
+ sky130_fd_sc_hd__a22o_1
X_09367_ _09367_/A vssd1 vssd1 vccd1 vccd1 _09367_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09298_ _09298_/A vssd1 vssd1 vccd1 vccd1 _09298_/Y sky130_fd_sc_hd__inv_2
X_08318_ _08318_/A vssd1 vssd1 vccd1 vccd1 _10000_/S sky130_fd_sc_hd__clkinv_8
X_08249_ _08249_/A _08249_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__or2_1
XFILLER_192_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _10289_/CLK _10211_/D vssd1 vssd1 vccd1 vccd1 _10211_/Q sky130_fd_sc_hd__dfxtp_1
X_10142_ _10244_/CLK _10142_/D vssd1 vssd1 vccd1 vccd1 _10142_/Q sky130_fd_sc_hd__dfxtp_1
X_10073_ _10205_/CLK _10073_/D vssd1 vssd1 vccd1 vccd1 _10073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10409_ _10442_/CLK _10409_/D vssd1 vssd1 vccd1 vccd1 _10409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05950_ _06111_/A vssd1 vssd1 vccd1 vccd1 _05950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05881_ _10269_/Q _10252_/Q _05812_/Y vssd1 vssd1 vccd1 vccd1 _05881_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _07604_/A _07615_/Y _07611_/X _07616_/X vssd1 vssd1 vccd1 vccd1 _07627_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07551_ _07815_/A vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__buf_1
X_06502_ _10092_/Q _06462_/A _08407_/A _06432_/A vssd1 vssd1 vccd1 vccd1 _06516_/B
+ sky130_fd_sc_hd__a22o_1
X_07482_ _07676_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__nor2_1
X_06433_ _06536_/A vssd1 vssd1 vccd1 vccd1 _06434_/A sky130_fd_sc_hd__clkbuf_2
X_09221_ _08868_/X _09220_/X _08868_/X _09220_/X vssd1 vssd1 vccd1 vccd1 _09222_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_61_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09152_ _09141_/X _09151_/X _09141_/X _09151_/X vssd1 vssd1 vccd1 vccd1 _09152_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06364_ _06364_/A vssd1 vssd1 vccd1 vccd1 _06364_/Y sky130_fd_sc_hd__inv_2
X_08103_ _08228_/A vssd1 vssd1 vccd1 vccd1 _08539_/A sky130_fd_sc_hd__clkbuf_2
X_05315_ _05315_/A vssd1 vssd1 vccd1 vccd1 _10346_/D sky130_fd_sc_hd__inv_2
XFILLER_174_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09083_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__or2_1
XFILLER_107_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06295_ _06281_/Y _10129_/Q _06285_/X vssd1 vssd1 vccd1 vccd1 _06295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05246_ _10362_/Q _05239_/X input25/X _05240_/X _05245_/X vssd1 vssd1 vccd1 vccd1
+ _10362_/D sky130_fd_sc_hd__o221a_1
X_08034_ _08025_/A _08025_/B _08026_/B vssd1 vssd1 vccd1 vccd1 _08034_/X sky130_fd_sc_hd__a21bo_1
X_05177_ _10428_/Q vssd1 vssd1 vccd1 vccd1 _05177_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _08896_/Y _08893_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09985_/X sky130_fd_sc_hd__mux2_2
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08936_ _10229_/Q _08978_/A _08936_/C vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__and3_1
XFILLER_123_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08867_ _08847_/Y _08866_/Y _10292_/Q _08847_/B vssd1 vssd1 vccd1 vccd1 _08867_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07818_ _09915_/X vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__inv_2
X_08798_ _08772_/A _08772_/B _08817_/A _08796_/Y _08797_/X vssd1 vssd1 vccd1 vccd1
+ _08798_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07749_ _07739_/X _07740_/X _07741_/X _07748_/X vssd1 vssd1 vccd1 vccd1 _07750_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _08377_/A _09282_/A _08377_/A _09417_/A _09311_/A vssd1 vssd1 vccd1 vccd1
+ _09464_/A sky130_fd_sc_hd__o221a_1
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10346_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _10330_/CLK _10125_/D vssd1 vssd1 vccd1 vccd1 _10125_/Q sky130_fd_sc_hd__dfxtp_1
X_10056_ _10421_/CLK _10056_/D vssd1 vssd1 vccd1 vccd1 _10056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06080_ _09757_/X _06028_/A _08179_/A _06031_/A _06032_/A vssd1 vssd1 vccd1 vccd1
+ _10176_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05100_ _05032_/X _05094_/X _10413_/Q _05095_/X _05097_/X vssd1 vssd1 vccd1 vccd1
+ _10413_/D sky130_fd_sc_hd__a221o_1
X_05031_ _10446_/Q _09940_/S _05030_/X _05013_/X _06182_/A vssd1 vssd1 vccd1 vccd1
+ _10446_/D sky130_fd_sc_hd__o221a_1
XFILLER_171_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09770_ _08195_/Y _10351_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__mux2_1
X_06982_ _07235_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07047_/D sky130_fd_sc_hd__nor2_4
X_08721_ _06020_/X _08718_/X _08281_/A _08720_/Y vssd1 vssd1 vccd1 vccd1 _08831_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_05933_ _10230_/Q vssd1 vssd1 vccd1 vccd1 _05933_/X sky130_fd_sc_hd__clkbuf_2
X_08652_ _08166_/X _10059_/Q _08107_/X _10058_/Q vssd1 vssd1 vccd1 vccd1 _08652_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07603_ _07603_/A _07677_/A vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__or2_4
X_05864_ _05799_/X _05820_/X _05799_/X _05820_/X vssd1 vssd1 vccd1 vccd1 _05865_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08583_ _08597_/A _08582_/X vssd1 vssd1 vccd1 vccd1 _08583_/X sky130_fd_sc_hd__or2b_1
X_05795_ _10258_/Q vssd1 vssd1 vccd1 vccd1 _05795_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07534_ _07813_/C vssd1 vssd1 vccd1 vccd1 _07811_/C sky130_fd_sc_hd__clkbuf_2
X_07465_ _07667_/B vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__buf_1
XFILLER_194_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ _09202_/A _09203_/A _09316_/C _09203_/Y vssd1 vssd1 vccd1 vccd1 _09205_/C
+ sky130_fd_sc_hd__a22o_1
X_06416_ _10079_/Q vssd1 vssd1 vccd1 vccd1 _06416_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _07396_/A vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__inv_2
XFILLER_182_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _09000_/X _09078_/A _09174_/A _09247_/A vssd1 vssd1 vccd1 vccd1 _09135_/X
+ sky130_fd_sc_hd__a211o_1
X_06347_ _06344_/A _06341_/X _06344_/A _06341_/X vssd1 vssd1 vccd1 vccd1 _06347_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_135_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09066_ _09066_/A vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__inv_2
X_06278_ _10234_/Q _05768_/B _06277_/A _05771_/B _06277_/Y vssd1 vssd1 vccd1 vccd1
+ _06278_/X sky130_fd_sc_hd__o32a_1
X_05229_ _10371_/Q _05221_/X input35/X _05223_/X _05227_/X vssd1 vssd1 vccd1 vccd1
+ _10371_/D sky130_fd_sc_hd__o221a_1
XFILLER_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08017_ _08017_/A _08017_/B vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__or2_1
XFILLER_150_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09968_ _08880_/Y _08876_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08919_ _08918_/A _08918_/B _08918_/Y vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__a21o_1
X_09899_ _10416_/Q _08065_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10108_ _10205_/CLK _10108_/D vssd1 vssd1 vccd1 vccd1 _10108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _10176_/CLK _10039_/D vssd1 vssd1 vccd1 vccd1 _10039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05580_ _10226_/Q vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__inv_2
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07250_ _07094_/A _07094_/B _07253_/B vssd1 vssd1 vccd1 vccd1 _07250_/X sky130_fd_sc_hd__a21o_1
X_06201_ _09701_/X _06196_/X _10102_/Q _06197_/X vssd1 vssd1 vccd1 vccd1 _10102_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07181_ _07181_/A vssd1 vssd1 vccd1 vccd1 _07182_/A sky130_fd_sc_hd__inv_2
X_06132_ _10146_/Q _06126_/X _10318_/Q _06130_/X _06128_/X vssd1 vssd1 vccd1 vccd1
+ _10146_/D sky130_fd_sc_hd__o221a_1
X_06063_ _09789_/X _06054_/X _08211_/A _06056_/X _06057_/X vssd1 vssd1 vccd1 vccd1
+ _10184_/D sky130_fd_sc_hd__o221a_1
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05014_ input47/X vssd1 vssd1 vccd1 vccd1 _05016_/A sky130_fd_sc_hd__inv_2
X_09822_ _08248_/X _10364_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09822_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09753_ _10417_/Q _08066_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09753_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08704_ _08704_/A _08704_/B _08704_/C _08703_/X vssd1 vssd1 vccd1 vccd1 _08705_/D
+ sky130_fd_sc_hd__or4b_4
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06965_ _06959_/Y _06964_/Y _06959_/Y _06964_/Y vssd1 vssd1 vccd1 vccd1 _06965_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09684_ _06457_/X input47/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05916_ _10237_/Q _05910_/X _05030_/X _05911_/X _05908_/X vssd1 vssd1 vccd1 vccd1
+ _10237_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06896_ _06931_/A _09893_/X _06942_/C _09668_/X _06895_/Y vssd1 vssd1 vccd1 vccd1
+ _06897_/B sky130_fd_sc_hd__o41a_1
X_08635_ _08745_/B vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__clkbuf_2
X_05847_ _07437_/A _10261_/Q _05787_/Y vssd1 vssd1 vccd1 vccd1 _05847_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08566_ _08783_/A _08562_/X _08138_/X _08565_/Y vssd1 vssd1 vccd1 vccd1 _08589_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05778_ input51/X _08321_/A _10266_/Q vssd1 vssd1 vccd1 vccd1 _05778_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ _07517_/A vssd1 vssd1 vccd1 vccd1 _07517_/Y sky130_fd_sc_hd__inv_2
X_08497_ _10073_/Q _08491_/B _08492_/B vssd1 vssd1 vccd1 vccd1 _08497_/X sky130_fd_sc_hd__a21bo_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ _10212_/Q vssd1 vssd1 vccd1 vccd1 _07613_/B sky130_fd_sc_hd__inv_2
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07379_ _07291_/X _07293_/X _07291_/X _07293_/X vssd1 vssd1 vccd1 vccd1 _07396_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_182_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09118_ _09117_/A _09117_/B _09166_/A vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__a21bo_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _10426_/CLK _10390_/D vssd1 vssd1 vccd1 vccd1 _10390_/Q sky130_fd_sc_hd__dfxtp_1
X_09049_ _05931_/X _09168_/B _09048_/X vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06750_ _10385_/Q vssd1 vssd1 vccd1 vccd1 _06750_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06681_ _10369_/Q _08724_/A vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__or2_2
X_05701_ _05741_/A vssd1 vssd1 vccd1 vccd1 _05701_/X sky130_fd_sc_hd__clkbuf_2
X_08420_ _08420_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08420_/Y sky130_fd_sc_hd__nor2_1
X_05632_ _05632_/A _05632_/B vssd1 vssd1 vccd1 vccd1 _05632_/X sky130_fd_sc_hd__and2_1
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08351_ _08351_/A _09544_/S vssd1 vssd1 vccd1 vccd1 _08351_/Y sky130_fd_sc_hd__nor2_1
X_05563_ _05489_/A _05489_/B _05489_/Y vssd1 vssd1 vccd1 vccd1 _05563_/Y sky130_fd_sc_hd__a21oi_1
X_08282_ _10200_/Q _08278_/Y _08264_/X _08285_/B vssd1 vssd1 vccd1 vccd1 _08282_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07302_ _07264_/X _07274_/X _07300_/X _07301_/X vssd1 vssd1 vccd1 vccd1 _07302_/X
+ sky130_fd_sc_hd__o22a_1
X_05494_ _05494_/A _05494_/B vssd1 vssd1 vccd1 vccd1 _05494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07233_ _07222_/X _07223_/X _07222_/X _07223_/X vssd1 vssd1 vccd1 vccd1 _07233_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_164_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07164_ _07164_/A _07164_/B vssd1 vssd1 vccd1 vccd1 _07176_/A sky130_fd_sc_hd__or2_1
XFILLER_160_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06115_ _10156_/Q _05891_/X _10328_/Q _06113_/X _06111_/X vssd1 vssd1 vccd1 vccd1
+ _10156_/D sky130_fd_sc_hd__o221a_1
X_07095_ _07095_/A _07253_/B vssd1 vssd1 vccd1 vccd1 _07095_/Y sky130_fd_sc_hd__nor2_1
X_06046_ _09821_/X _06043_/X _10192_/Q _06044_/X _06045_/X vssd1 vssd1 vccd1 vccd1
+ _10192_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09805_ _09804_/X input22/X _09821_/S vssd1 vssd1 vccd1 vccd1 _09805_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07997_ _08016_/A vssd1 vssd1 vccd1 vccd1 _07997_/Y sky130_fd_sc_hd__inv_2
X_09736_ _06808_/Y _10401_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10067_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06948_ _06866_/A _06960_/B _07028_/A _06949_/D vssd1 vssd1 vccd1 vccd1 _06950_/A
+ sky130_fd_sc_hd__o22a_1
X_09667_ _10149_/Q _10165_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09667_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08618_ _08618_/A _09942_/X vssd1 vssd1 vccd1 vccd1 _10040_/D sky130_fd_sc_hd__or2_1
XFILLER_82_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06879_ _07028_/A _06960_/B _06878_/X vssd1 vssd1 vccd1 vccd1 _06880_/B sky130_fd_sc_hd__or3b_1
XFILLER_202_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09598_ _08449_/Y _08448_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09598_/X sky130_fd_sc_hd__mux2_2
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _10050_/Q _08468_/B _08469_/B vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__a21bo_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10442_ _10442_/CLK _10442_/D vssd1 vssd1 vccd1 vccd1 _10442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10437_/CLK _10373_/D vssd1 vssd1 vccd1 vccd1 _10373_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07920_ _07919_/X _07776_/X _07919_/X _07776_/X vssd1 vssd1 vccd1 vccd1 _07920_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _07851_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07851_/Y sky130_fd_sc_hd__nor2_1
Xinput2 io_QEI_ChB vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_06802_ _06802_/A _06802_/B vssd1 vssd1 vccd1 vccd1 _06802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07782_ _07777_/A _07504_/B _07780_/Y _07781_/Y vssd1 vssd1 vccd1 vccd1 _07782_/Y
+ sky130_fd_sc_hd__o31ai_2
X_06733_ _10384_/Q vssd1 vssd1 vccd1 vccd1 _06733_/Y sky130_fd_sc_hd__inv_2
X_09521_ _09520_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09521_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__or2_1
X_06664_ _06664_/A _06664_/B vssd1 vssd1 vccd1 vccd1 _06665_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06595_ _08450_/A _06489_/A _06590_/X _06592_/X vssd1 vssd1 vccd1 vccd1 _06595_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09383_ _09384_/B vssd1 vssd1 vccd1 vccd1 _09383_/Y sky130_fd_sc_hd__inv_2
X_08403_ _08403_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08403_/Y sky130_fd_sc_hd__nor2_1
X_05615_ _05615_/A vssd1 vssd1 vccd1 vccd1 _10007_/S sky130_fd_sc_hd__inv_2
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08334_ _09300_/A vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__buf_2
X_05546_ _05546_/A vssd1 vssd1 vccd1 vccd1 _05546_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08265_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08269_/B sky130_fd_sc_hd__or2_1
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05477_ _10008_/X vssd1 vssd1 vccd1 vccd1 _05478_/B sky130_fd_sc_hd__inv_2
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08196_ _08782_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__or2_2
X_07216_ _07214_/X _07215_/X _07214_/X _07215_/X vssd1 vssd1 vccd1 vccd1 _07222_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07147_ _07147_/A _09884_/X vssd1 vssd1 vccd1 vccd1 _07147_/X sky130_fd_sc_hd__or2_1
XFILLER_173_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07078_ _07067_/A _07067_/B _07067_/X vssd1 vssd1 vccd1 vccd1 _07079_/B sky130_fd_sc_hd__a21bo_1
X_06029_ _10197_/Q vssd1 vssd1 vccd1 vccd1 _06263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE3_1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09719_ _06788_/X _10384_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10050_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10425_ _10426_/CLK _10425_/D vssd1 vssd1 vccd1 vccd1 _10425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _10421_/CLK _10356_/D vssd1 vssd1 vccd1 vccd1 _10356_/Q sky130_fd_sc_hd__dfxtp_2
X_10287_ _10289_/CLK _10287_/D vssd1 vssd1 vccd1 vccd1 _10287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05400_ _06185_/A _05718_/A _05400_/C vssd1 vssd1 vccd1 vccd1 _05400_/X sky130_fd_sc_hd__and3_1
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06380_ _10138_/Q vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__inv_2
XFILLER_202_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05331_ _05326_/B _05282_/X _05330_/Y _05322_/X _05305_/A vssd1 vssd1 vccd1 vccd1
+ _05332_/A sky130_fd_sc_hd__o32a_1
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05262_ _05089_/X _05251_/X _08760_/A _05252_/X _05253_/X vssd1 vssd1 vccd1 vccd1
+ _10354_/D sky130_fd_sc_hd__a221o_1
X_08050_ _08017_/A _08017_/B _08018_/B vssd1 vssd1 vccd1 vccd1 _08050_/X sky130_fd_sc_hd__a21bo_1
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07001_ _07108_/B vssd1 vssd1 vccd1 vccd1 _07126_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05193_ _05193_/A vssd1 vssd1 vccd1 vccd1 _05193_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ _10288_/Q _08852_/B _08852_/Y vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08883_ _10226_/Q _08978_/A _10227_/Q _09168_/C vssd1 vssd1 vccd1 vccd1 _08889_/A
+ sky130_fd_sc_hd__and4_1
X_07903_ _07903_/A _07903_/B vssd1 vssd1 vccd1 vccd1 _07904_/B sky130_fd_sc_hd__or2_1
XFILLER_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07834_ _07823_/A _07823_/B _07823_/X vssd1 vssd1 vccd1 vccd1 _07835_/B sky130_fd_sc_hd__a21bo_1
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07765_ _07765_/A vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06716_ _06714_/Y _06715_/Y _08729_/A vssd1 vssd1 vccd1 vccd1 _06718_/A sky130_fd_sc_hd__o21ai_1
XFILLER_112_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09504_ _09503_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07696_ _07684_/A _07684_/B _07721_/A vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__a21o_1
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09435_ _09434_/A _09434_/B _09434_/X vssd1 vssd1 vccd1 vccd1 _09435_/X sky130_fd_sc_hd__a21bo_1
X_06647_ _06647_/A vssd1 vssd1 vccd1 vccd1 _06647_/Y sky130_fd_sc_hd__inv_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06578_ _10107_/Q vssd1 vssd1 vccd1 vccd1 _08446_/A sky130_fd_sc_hd__inv_2
X_09366_ _09170_/A _09251_/X _09428_/C _09365_/X vssd1 vssd1 vccd1 vccd1 _09367_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _09297_/A _09235_/X vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__or2b_1
X_08317_ _08317_/A vssd1 vssd1 vccd1 vccd1 _09999_/S sky130_fd_sc_hd__clkinv_8
X_05529_ _10011_/X _10015_/X _05472_/Y _05538_/A vssd1 vssd1 vccd1 vccd1 _05529_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08248_ _10193_/Q _06259_/B _08247_/Y vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08179_ _08179_/A _08184_/A vssd1 vssd1 vccd1 vccd1 _08179_/Y sky130_fd_sc_hd__nor2_1
X_10210_ _10217_/CLK _10210_/D vssd1 vssd1 vccd1 vccd1 _10210_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10141_ _10330_/CLK _10141_/D vssd1 vssd1 vccd1 vccd1 _10141_/Q sky130_fd_sc_hd__dfxtp_1
X_10072_ _10437_/CLK _10072_/D vssd1 vssd1 vccd1 vccd1 _10072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10408_ _10442_/CLK _10408_/D vssd1 vssd1 vccd1 vccd1 _10408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10339_ _10343_/CLK _10339_/D vssd1 vssd1 vccd1 vccd1 _10339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05880_ _10253_/Q _05871_/X _05863_/X _06821_/A _05866_/X vssd1 vssd1 vccd1 vccd1
+ _10253_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07550_ _07550_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _07550_/X sky130_fd_sc_hd__or2_1
X_06501_ _10092_/Q vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__inv_2
X_09220_ _08845_/A _08845_/B _08845_/Y vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__a21o_1
X_07481_ _07634_/A vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__clkbuf_2
X_06432_ _06432_/A vssd1 vssd1 vccd1 vccd1 _06536_/A sky130_fd_sc_hd__clkbuf_2
X_09151_ _09192_/A _09101_/B _09150_/Y _09101_/Y _09150_/A vssd1 vssd1 vccd1 vccd1
+ _09151_/X sky130_fd_sc_hd__o32a_1
X_06363_ _06351_/A _10136_/Q _06352_/A _06355_/Y vssd1 vssd1 vccd1 vccd1 _06364_/A
+ sky130_fd_sc_hd__o22a_1
X_08102_ _10188_/Q vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__inv_2
X_05314_ _10346_/Q _05282_/X _05312_/A _05310_/Y _05313_/X vssd1 vssd1 vccd1 vccd1
+ _05315_/A sky130_fd_sc_hd__o32a_1
X_09082_ _09076_/X _09081_/X _09076_/X _09081_/X vssd1 vssd1 vccd1 vccd1 _09085_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06294_ _06294_/A _06294_/B vssd1 vssd1 vccd1 vccd1 _06294_/X sky130_fd_sc_hd__or2_1
X_08033_ _07411_/A _07411_/B _07412_/B vssd1 vssd1 vccd1 vccd1 _08033_/X sky130_fd_sc_hd__a21bo_1
X_05245_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05245_/X sky130_fd_sc_hd__buf_2
X_05176_ _10396_/Q vssd1 vssd1 vccd1 vccd1 _05176_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _08892_/Y _08890_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__mux2_1
X_08935_ _09038_/C vssd1 vssd1 vccd1 vccd1 _08993_/C sky130_fd_sc_hd__inv_2
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08866_ _10291_/Q _07445_/X _08848_/X _08865_/X vssd1 vssd1 vccd1 vccd1 _08866_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08797_ _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08797_/X sky130_fd_sc_hd__or2_1
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07817_ _07819_/A _09914_/X vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__nor2_1
XFILLER_72_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07748_ _07742_/X _07744_/X _07745_/X _07747_/X vssd1 vssd1 vccd1 vccd1 _07748_/X
+ sky130_fd_sc_hd__o22a_1
X_07679_ _07679_/A vssd1 vssd1 vccd1 vccd1 _07680_/B sky130_fd_sc_hd__inv_2
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09418_ _09418_/A _09418_/B vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__or2_1
XFILLER_40_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _09347_/Y _09393_/B _09347_/Y _09393_/B vssd1 vssd1 vccd1 vccd1 _09350_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10244_/CLK _10124_/D vssd1 vssd1 vccd1 vccd1 _10124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10055_ _10421_/CLK _10055_/D vssd1 vssd1 vccd1 vccd1 _10055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05030_ input44/X vssd1 vssd1 vccd1 vccd1 _05030_/X sky130_fd_sc_hd__buf_2
XFILLER_152_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06981_ _06992_/A vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__inv_2
X_08720_ _06630_/Y _08719_/Y _08717_/Y vssd1 vssd1 vccd1 vccd1 _08720_/Y sky130_fd_sc_hd__o21bai_1
X_05932_ _05931_/X _05927_/X _05093_/X _05928_/X _05918_/X vssd1 vssd1 vccd1 vccd1
+ _10231_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08651_ _08646_/X _08649_/X _08664_/B vssd1 vssd1 vccd1 vccd1 _08651_/Y sky130_fd_sc_hd__a21oi_1
X_05863_ _05863_/A vssd1 vssd1 vccd1 vccd1 _05863_/X sky130_fd_sc_hd__clkbuf_2
X_07602_ _09921_/X vssd1 vssd1 vccd1 vccd1 _07677_/A sky130_fd_sc_hd__clkbuf_2
X_08582_ _08596_/A _08596_/B _08596_/C _08582_/D vssd1 vssd1 vccd1 vccd1 _08582_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05794_ _10275_/Q vssd1 vssd1 vccd1 vccd1 _07445_/A sky130_fd_sc_hd__inv_2
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07533_ _07587_/D vssd1 vssd1 vccd1 vccd1 _07813_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07464_ _10214_/Q vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__inv_2
XFILLER_179_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _09203_/A vssd1 vssd1 vccd1 vccd1 _09203_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06415_ _06856_/A vssd1 vssd1 vccd1 vccd1 _06415_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09134_ _09026_/X _09133_/X _09026_/X _09133_/X vssd1 vssd1 vccd1 vccd1 _09134_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_07395_ _07395_/A vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__inv_2
XFILLER_22_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06346_ _06344_/A _06344_/B _06345_/Y vssd1 vssd1 vccd1 vccd1 _06346_/Y sky130_fd_sc_hd__a21oi_1
X_09065_ _08848_/X _08865_/X _08848_/X _08865_/X vssd1 vssd1 vccd1 vccd1 _09066_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06277_ _06277_/A vssd1 vssd1 vccd1 vccd1 _06277_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05228_ _10372_/Q _05221_/X input36/X _05223_/X _05227_/X vssd1 vssd1 vccd1 vccd1
+ _10372_/D sky130_fd_sc_hd__o221a_1
X_08016_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08017_/B sky130_fd_sc_hd__or2_1
XFILLER_116_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05159_ _10400_/Q vssd1 vssd1 vccd1 vccd1 _06616_/C sky130_fd_sc_hd__inv_2
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _09966_/X _06629_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09967_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08918_ _08918_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08918_/Y sky130_fd_sc_hd__nor2_2
X_09898_ _10415_/Q _08063_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08849_ _10290_/Q vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__inv_2
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ _10207_/CLK _10107_/D vssd1 vssd1 vccd1 vccd1 _10107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10038_ _10205_/CLK _10038_/D vssd1 vssd1 vccd1 vccd1 _10039_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_209_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06200_ _09702_/X _06196_/X _10103_/Q _06197_/X vssd1 vssd1 vccd1 vccd1 _10103_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07180_ _07180_/A _07180_/B vssd1 vssd1 vccd1 vccd1 _07180_/X sky130_fd_sc_hd__or2_1
XFILLER_184_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06131_ _10147_/Q _06126_/X _10319_/Q _06130_/X _06128_/X vssd1 vssd1 vccd1 vccd1
+ _10147_/D sky130_fd_sc_hd__o221a_1
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06062_ _10184_/Q vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__buf_2
X_05013_ _05013_/A vssd1 vssd1 vccd1 vccd1 _05013_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09821_ _09820_/X input26/X _09821_/S vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09752_ _09751_/X _10210_/Q _10000_/S vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__mux2_1
X_08703_ _08077_/X _10045_/Q _08702_/Y _08658_/X _08655_/X vssd1 vssd1 vccd1 vccd1
+ _08703_/X sky130_fd_sc_hd__o2111a_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06964_ _06960_/X _06963_/X _06960_/X _06963_/X vssd1 vssd1 vccd1 vccd1 _06964_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_09683_ _06452_/X input46/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__mux2_1
X_05915_ _05028_/X _05896_/X _10238_/Q _05897_/X _05274_/X vssd1 vssd1 vccd1 vccd1
+ _10238_/D sky130_fd_sc_hd__a221o_1
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06895_ _06898_/C _06895_/B vssd1 vssd1 vccd1 vccd1 _06895_/Y sky130_fd_sc_hd__nand2_1
X_08634_ _08752_/B vssd1 vssd1 vccd1 vccd1 _08745_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_5_clock clkbuf_2_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10176_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05846_ _10262_/Q _05780_/X _05842_/X _06855_/A _05845_/X vssd1 vssd1 vccd1 vccd1
+ _10262_/D sky130_fd_sc_hd__o221a_1
XFILLER_199_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08565_ _08467_/A _08467_/B _08468_/B vssd1 vssd1 vccd1 vccd1 _08565_/Y sky130_fd_sc_hd__o21ai_1
X_05777_ _05777_/A vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__inv_2
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ _10217_/Q _07516_/B _07527_/A vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__and3_1
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08496_ _10074_/Q _08492_/B _08493_/Y vssd1 vssd1 vccd1 vccd1 _08496_/Y sky130_fd_sc_hd__a21oi_1
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07447_ _07445_/X _07431_/Y _07439_/B vssd1 vssd1 vccd1 vccd1 _07447_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07378_ _07287_/X _07294_/X _07287_/X _07294_/X vssd1 vssd1 vccd1 vccd1 _07395_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _09117_/A _09117_/B vssd1 vssd1 vccd1 vccd1 _09166_/A sky130_fd_sc_hd__or2_2
X_06329_ _10241_/Q vssd1 vssd1 vccd1 vccd1 _06330_/A sky130_fd_sc_hd__inv_2
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09048_ _09070_/A _09096_/A vssd1 vssd1 vccd1 vccd1 _09048_/X sky130_fd_sc_hd__or2_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06680_ _10368_/Q _08727_/A vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__or2_2
X_05700_ _10298_/Q _05467_/X _10282_/Q _05699_/X _05660_/X vssd1 vssd1 vccd1 vccd1
+ _10298_/D sky130_fd_sc_hd__o221a_1
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05631_ _05631_/A vssd1 vssd1 vccd1 vccd1 _05631_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _09932_/X _08364_/B vssd1 vssd1 vccd1 vccd1 _08350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _07264_/X _07274_/X _07264_/X _07274_/X vssd1 vssd1 vccd1 vccd1 _07301_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05562_ _05562_/A vssd1 vssd1 vccd1 vccd1 _05562_/Y sky130_fd_sc_hd__inv_2
X_08281_ _08281_/A _08281_/B vssd1 vssd1 vccd1 vccd1 _08285_/B sky130_fd_sc_hd__or2_2
XFILLER_177_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05493_ _10005_/X vssd1 vssd1 vccd1 vccd1 _05494_/B sky130_fd_sc_hd__inv_2
XFILLER_177_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07232_ _07232_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__or2_1
XFILLER_192_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07163_ _07156_/X _07157_/X _07156_/X _07157_/X vssd1 vssd1 vccd1 vccd1 _07181_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06114_ _10157_/Q _05891_/X _10329_/Q _06113_/X _06111_/X vssd1 vssd1 vccd1 vccd1
+ _10157_/D sky130_fd_sc_hd__o221a_1
XFILLER_172_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07094_ _07094_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _07253_/B sky130_fd_sc_hd__nor2_2
X_06045_ _06070_/A vssd1 vssd1 vccd1 vccd1 _06045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09803_/X _08229_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07996_ _07626_/A _07626_/B _07639_/B vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__a21oi_4
X_09735_ _06807_/Y _10400_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10066_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06947_ _06944_/X _06946_/X _06944_/X _06946_/X vssd1 vssd1 vccd1 vccd1 _06947_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09666_ _10148_/Q _10164_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ _08617_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _10078_/D sky130_fd_sc_hd__nand2_1
XFILLER_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06878_ _07031_/A _06949_/D vssd1 vssd1 vccd1 vccd1 _06878_/X sky130_fd_sc_hd__or2_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09597_ _08447_/Y _08446_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05829_ _05704_/X _10263_/Q _05785_/Y _05828_/X vssd1 vssd1 vccd1 vccd1 _05829_/X
+ sky130_fd_sc_hd__o2bb2a_2
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _10051_/Q _08469_/B _08470_/B vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__a21bo_1
X_08479_ _10061_/Q _08479_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__or2_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _10442_/CLK _10441_/D vssd1 vssd1 vccd1 vccd1 _10441_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10372_ _10436_/CLK _10372_/D vssd1 vssd1 vccd1 vccd1 _10372_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07850_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__nor2_2
X_06801_ _06802_/A _06801_/B vssd1 vssd1 vccd1 vccd1 _06801_/Y sky130_fd_sc_hd__nor2_1
X_07781_ _07777_/A _07504_/B _07780_/Y vssd1 vssd1 vccd1 vccd1 _07781_/Y sky130_fd_sc_hd__o21ai_1
Xinput3 io_clo_test vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
XFILLER_209_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06732_ _08761_/A _06667_/B _06668_/B vssd1 vssd1 vccd1 vccd1 _06791_/B sky130_fd_sc_hd__a21boi_4
XFILLER_83_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09520_ _09519_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09520_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _09451_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09451_/Y sky130_fd_sc_hd__nor2_1
X_06663_ _06606_/X _08632_/A _06652_/Y _06662_/X vssd1 vssd1 vccd1 vccd1 _06664_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06594_ _10110_/Q vssd1 vssd1 vccd1 vccd1 _08452_/A sky130_fd_sc_hd__inv_2
X_09382_ _09338_/X _09381_/X _09338_/X _09381_/X vssd1 vssd1 vccd1 vccd1 _09384_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _09517_/X _08414_/B vssd1 vssd1 vccd1 vccd1 _08402_/Y sky130_fd_sc_hd__nor2_1
X_05614_ _05614_/A vssd1 vssd1 vccd1 vccd1 _05614_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05545_ _09902_/X _05544_/X _09902_/X _05544_/X vssd1 vssd1 vccd1 vccd1 _05632_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08333_ _09174_/A vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__buf_1
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08264_ _08264_/A vssd1 vssd1 vccd1 vccd1 _08264_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05476_ _10016_/X vssd1 vssd1 vccd1 vccd1 _05478_/A sky130_fd_sc_hd__inv_2
X_08195_ _08138_/X _06246_/B _06247_/B vssd1 vssd1 vccd1 vccd1 _08195_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07215_ _07223_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07215_/X sky130_fd_sc_hd__or2_1
X_07146_ _07146_/A _07212_/B _07146_/C _07164_/B vssd1 vssd1 vccd1 vccd1 _07146_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_105_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10289_/CLK sky130_fd_sc_hd__clkbuf_16
X_07077_ _07077_/A _07077_/B vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__or2_1
X_06028_ _06028_/A vssd1 vssd1 vccd1 vccd1 _06028_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE3_2 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09718_ _09717_/X _10383_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10049_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _07977_/Y _07978_/X _07977_/Y _07978_/X vssd1 vssd1 vccd1 vccd1 _07979_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_19_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _10115_/Q input45/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10424_ _10426_/CLK _10424_/D vssd1 vssd1 vccd1 vccd1 _10424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10355_ _10421_/CLK _10355_/D vssd1 vssd1 vccd1 vccd1 _10355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10286_ _10289_/CLK _10286_/D vssd1 vssd1 vccd1 vccd1 _10286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05330_ _10341_/Q _05330_/B vssd1 vssd1 vccd1 vccd1 _05330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05261_ _10354_/Q vssd1 vssd1 vccd1 vccd1 _08760_/A sky130_fd_sc_hd__buf_2
XFILLER_127_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05192_ _05185_/X _10390_/Q _05186_/X _09609_/X _05189_/X vssd1 vssd1 vccd1 vccd1
+ _10390_/D sky130_fd_sc_hd__o221a_1
X_07000_ _09889_/X vssd1 vssd1 vccd1 vccd1 _07108_/B sky130_fd_sc_hd__inv_2
XFILLER_170_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ _08950_/A _08950_/B _08985_/A vssd1 vssd1 vccd1 vccd1 _08951_/X sky130_fd_sc_hd__a21bo_1
XFILLER_102_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08882_ _08882_/A vssd1 vssd1 vccd1 vccd1 _09168_/C sky130_fd_sc_hd__inv_2
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07902_ _07903_/A _07903_/B vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07833_ _07833_/A _07813_/X vssd1 vssd1 vccd1 vccd1 _07835_/A sky130_fd_sc_hd__or2b_1
XFILLER_110_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07764_ _07916_/A _07916_/C vssd1 vssd1 vccd1 vccd1 _07764_/X sky130_fd_sc_hd__or2_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06715_ _08731_/A vssd1 vssd1 vccd1 vccd1 _06715_/Y sky130_fd_sc_hd__inv_2
X_09503_ _09502_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09503_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07695_ _07695_/A vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__inv_2
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _09434_/A _09434_/B vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__or2_1
X_06646_ _08626_/A _05273_/X _06645_/Y vssd1 vssd1 vccd1 vccd1 _06647_/A sky130_fd_sc_hd__a21oi_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06577_ _06580_/A _06576_/X _06580_/A _06576_/X vssd1 vssd1 vccd1 vccd1 _06577_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09365_ _09245_/A _09417_/A _09310_/A _09247_/A vssd1 vssd1 vccd1 vccd1 _09365_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09296_ _09390_/C _09295_/A _09343_/C _09295_/Y vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__a22o_1
X_08316_ _08316_/A vssd1 vssd1 vccd1 vccd1 _09998_/S sky130_fd_sc_hd__clkinv_8
X_05528_ _10010_/X _10020_/X _05475_/Y _05542_/A vssd1 vssd1 vccd1 vccd1 _05538_/A
+ sky130_fd_sc_hd__o22a_1
X_08247_ _08247_/A vssd1 vssd1 vccd1 vccd1 _08247_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05459_ _05456_/Y _05457_/Y _05458_/Y vssd1 vssd1 vccd1 vccd1 _05459_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08178_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__buf_4
XFILLER_137_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ _07124_/X _07128_/X _07124_/X _07128_/X vssd1 vssd1 vccd1 vccd1 _07129_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ _10330_/CLK _10140_/D vssd1 vssd1 vccd1 vccd1 _10140_/Q sky130_fd_sc_hd__dfxtp_1
X_10071_ _10437_/CLK _10071_/D vssd1 vssd1 vccd1 vccd1 _10071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _10442_/CLK _10407_/D vssd1 vssd1 vccd1 vccd1 _10407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ _10343_/CLK _10338_/D vssd1 vssd1 vccd1 vccd1 _10338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10269_ _10298_/CLK _10269_/D vssd1 vssd1 vccd1 vccd1 _10269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06500_ _06516_/A _06499_/Y _06494_/A _06499_/A vssd1 vssd1 vccd1 vccd1 _06500_/X
+ sky130_fd_sc_hd__o22a_1
X_07480_ _09936_/X vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06431_ _06487_/A vssd1 vssd1 vccd1 vccd1 _06432_/A sky130_fd_sc_hd__clkbuf_2
X_09150_ _09150_/A vssd1 vssd1 vccd1 vccd1 _09150_/Y sky130_fd_sc_hd__inv_2
X_06362_ _06362_/A vssd1 vssd1 vccd1 vccd1 _06362_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ _06625_/Y _10206_/Q _10377_/Q _08307_/A _08100_/X vssd1 vssd1 vccd1 vccd1
+ _08119_/A sky130_fd_sc_hd__o221a_1
XFILLER_159_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05313_ _10175_/Q _05313_/B vssd1 vssd1 vccd1 vccd1 _05313_/X sky130_fd_sc_hd__and2_1
X_09081_ _09078_/Y _09080_/X _09078_/Y _09080_/X vssd1 vssd1 vccd1 vccd1 _09081_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06293_ _06293_/A _10130_/Q vssd1 vssd1 vccd1 vccd1 _06294_/B sky130_fd_sc_hd__nor2_1
X_05244_ _05468_/A vssd1 vssd1 vccd1 vccd1 _05737_/A sky130_fd_sc_hd__clkbuf_2
X_08032_ _08026_/A _08026_/B _08027_/B vssd1 vssd1 vccd1 vccd1 _08032_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 io_wb_dat_i[9] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_4
X_05175_ _05179_/A _05175_/B vssd1 vssd1 vccd1 vccd1 _10397_/D sky130_fd_sc_hd__nor2_1
XFILLER_115_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _09167_/X _09165_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09983_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _08934_/A _09985_/X vssd1 vssd1 vccd1 vccd1 _09038_/C sky130_fd_sc_hd__or2_4
XFILLER_130_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _10290_/Q _05797_/Y _08850_/Y _08864_/X vssd1 vssd1 vccd1 vccd1 _08865_/X
+ sky130_fd_sc_hd__o22a_1
X_08796_ _08780_/X _08818_/A _08794_/X _08819_/C vssd1 vssd1 vccd1 vccd1 _08796_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07816_ _07814_/X _07815_/X _07814_/X _07815_/X vssd1 vssd1 vccd1 vccd1 _07823_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07747_/X sky130_fd_sc_hd__or2_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _07678_/A _07777_/C vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__or2_2
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06629_ _10372_/Q vssd1 vssd1 vccd1 vccd1 _06629_/Y sky130_fd_sc_hd__inv_2
X_09417_ _09417_/A vssd1 vssd1 vccd1 vccd1 _09417_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _09343_/C _09295_/Y _09296_/X _09301_/X vssd1 vssd1 vccd1 vccd1 _09393_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09279_/A vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__inv_2
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _10330_/CLK _10123_/D vssd1 vssd1 vccd1 vccd1 _10123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10054_ _10421_/CLK _10054_/D vssd1 vssd1 vccd1 vccd1 _10054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06980_ _07311_/A _07311_/B _06985_/A _06970_/A _06976_/A vssd1 vssd1 vccd1 vccd1
+ _06980_/X sky130_fd_sc_hd__o32a_1
X_05931_ _10231_/Q vssd1 vssd1 vccd1 vccd1 _05931_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _08160_/X _10056_/Q _08104_/X _10057_/Q vssd1 vssd1 vccd1 vccd1 _08664_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05862_ _10258_/Q _05851_/X _05842_/X _06834_/A _05845_/X vssd1 vssd1 vccd1 vccd1
+ _10258_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07601_ _09920_/X vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__clkbuf_2
X_08581_ _08594_/B _08581_/B vssd1 vssd1 vccd1 vccd1 _08582_/D sky130_fd_sc_hd__nor2_4
XFILLER_81_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05793_ _05790_/A _10259_/Q _05791_/A _05792_/Y vssd1 vssd1 vccd1 vccd1 _05793_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07532_ _10213_/Q vssd1 vssd1 vccd1 vccd1 _07587_/D sky130_fd_sc_hd__inv_2
XFILLER_179_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07463_ _07678_/A vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_210_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09202_ _09202_/A vssd1 vssd1 vccd1 vccd1 _09316_/C sky130_fd_sc_hd__inv_2
X_06414_ _06855_/A vssd1 vssd1 vccd1 vccd1 _06414_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _09294_/A _09251_/A _09180_/C _09132_/X vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07394_ _07394_/A vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__inv_2
X_06345_ _06345_/A vssd1 vssd1 vccd1 vccd1 _06345_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09064_ _09063_/A _09063_/B _09112_/A vssd1 vssd1 vccd1 vccd1 _09064_/X sky130_fd_sc_hd__a21bo_1
X_06276_ _10235_/Q _08335_/A _06275_/Y _10128_/Q vssd1 vssd1 vccd1 vccd1 _06277_/A
+ sky130_fd_sc_hd__o22a_1
X_05227_ _05236_/A vssd1 vssd1 vccd1 vccd1 _05227_/X sky130_fd_sc_hd__clkbuf_2
X_08015_ _08015_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__nand2_1
X_05158_ _05678_/A vssd1 vssd1 vccd1 vccd1 _05179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _06615_/C _08162_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05089_ input48/X vssd1 vssd1 vccd1 vccd1 _05089_/X sky130_fd_sc_hd__buf_4
X_09897_ _06239_/X _06235_/A _10041_/Q vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__mux2_4
X_08917_ _08915_/X _08916_/Y _08915_/X _08916_/Y vssd1 vssd1 vccd1 vccd1 _08918_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08848_ _10291_/Q _07445_/X _10291_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _08848_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08779_ _08630_/X _08778_/X _08630_/X _08778_/X vssd1 vssd1 vccd1 vccd1 _08783_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10106_ _10207_/CLK _10106_/D vssd1 vssd1 vccd1 vccd1 _10106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10037_ _10205_/CLK input2/X vssd1 vssd1 vccd1 vccd1 _10038_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06130_ _06130_/A vssd1 vssd1 vccd1 vccd1 _06130_/X sky130_fd_sc_hd__buf_1
XFILLER_172_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06061_ _09793_/X _06054_/X _10185_/Q _06056_/X _06057_/X vssd1 vssd1 vccd1 vccd1
+ _10185_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05012_ _05012_/A vssd1 vssd1 vccd1 vccd1 _09940_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09820_ _09819_/X _08246_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09751_ _09750_/X _10218_/Q _09999_/S vssd1 vssd1 vccd1 vccd1 _09751_/X sky130_fd_sc_hd__mux2_1
X_06963_ _06961_/Y _06962_/X _06961_/Y _06962_/X vssd1 vssd1 vccd1 vccd1 _06963_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_08702_ _10177_/Q _08460_/Y _08121_/X _10052_/Q vssd1 vssd1 vccd1 vccd1 _08702_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05914_ _10239_/Q _05910_/X _05093_/X _05911_/X _05908_/X vssd1 vssd1 vccd1 vccd1
+ _10239_/D sky130_fd_sc_hd__o221a_1
X_09682_ _06448_/Y input45/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__mux2_1
X_06894_ _07108_/A _06912_/B _06894_/C vssd1 vssd1 vccd1 vccd1 _06895_/B sky130_fd_sc_hd__and3_1
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08633_ _08758_/B vssd1 vssd1 vccd1 vccd1 _08752_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05845_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05845_/X sky130_fd_sc_hd__clkbuf_2
X_08564_ _08554_/X _08560_/X _08591_/A vssd1 vssd1 vccd1 vccd1 _08564_/Y sky130_fd_sc_hd__a21oi_1
X_05776_ _05944_/B _06137_/A vssd1 vssd1 vccd1 vccd1 _05777_/A sky130_fd_sc_hd__or2_2
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07515_ _07678_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__or2_1
X_08495_ _08454_/Y _08493_/Y _08494_/X vssd1 vssd1 vccd1 vccd1 _08495_/Y sky130_fd_sc_hd__o21ai_1
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07446_ _05790_/A _07439_/B _07440_/B vssd1 vssd1 vccd1 vccd1 _07446_/X sky130_fd_sc_hd__a21bo_1
XFILLER_195_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07377_ _07296_/A _07296_/B _07296_/Y vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__o21ai_2
XFILLER_182_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _09117_/B vssd1 vssd1 vccd1 vccd1 _09116_/Y sky130_fd_sc_hd__inv_2
X_06328_ _06322_/Y _06327_/A _06322_/A _06327_/Y vssd1 vssd1 vccd1 vccd1 _06328_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _09089_/B vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__inv_2
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06259_ _10193_/Q _06259_/B vssd1 vssd1 vccd1 vccd1 _08247_/A sky130_fd_sc_hd__or2_1
XFILLER_163_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09023_/Y _09022_/B _09986_/S vssd1 vssd1 vccd1 vccd1 _09949_/X sky130_fd_sc_hd__mux2_2
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05630_ _05646_/A _05630_/B vssd1 vssd1 vccd1 vccd1 _10312_/D sky130_fd_sc_hd__nor2_1
XFILLER_17_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05561_ _09975_/X _05560_/X _09975_/X _05560_/X vssd1 vssd1 vccd1 vccd1 _05561_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07300_ _07275_/X _07279_/X _07280_/X _07299_/Y vssd1 vssd1 vccd1 vccd1 _07300_/X
+ sky130_fd_sc_hd__o22a_1
X_08280_ _08169_/X _08275_/Y _06267_/B vssd1 vssd1 vccd1 vccd1 _08280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05492_ _09993_/X vssd1 vssd1 vccd1 vccd1 _05494_/A sky130_fd_sc_hd__inv_2
XFILLER_192_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07231_ _07222_/A _07222_/B _07222_/X vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__a21bo_1
XFILLER_192_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07162_ _07158_/X _07161_/X _07158_/X _07161_/X vssd1 vssd1 vccd1 vccd1 _07162_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_145_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06113_ _06130_/A vssd1 vssd1 vccd1 vccd1 _06113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07093_ _07093_/A _07093_/B vssd1 vssd1 vccd1 vccd1 _07094_/B sky130_fd_sc_hd__or2_1
XFILLER_172_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06044_ _06069_/A vssd1 vssd1 vccd1 vccd1 _06044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _10359_/Q _09802_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _07747_/A _07747_/B _07747_/X vssd1 vssd1 vccd1 vccd1 _08012_/A sky130_fd_sc_hd__a21bo_1
X_09734_ _06806_/Y _10399_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10065_/D sky130_fd_sc_hd__mux2_1
X_06946_ _06946_/A _06946_/B vssd1 vssd1 vccd1 vccd1 _06946_/X sky130_fd_sc_hd__or2_1
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09665_ _10147_/Q _10163_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06877_ _09893_/X vssd1 vssd1 vccd1 vccd1 _06960_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _08616_/A _08616_/B vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__nand2_1
X_05828_ _05786_/A _10262_/Q _05786_/Y _05827_/X vssd1 vssd1 vccd1 vccd1 _05828_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09596_ _08445_/X _08444_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09596_/X sky130_fd_sc_hd__mux2_2
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08774_/A _08547_/B vssd1 vssd1 vccd1 vccd1 _08547_/X sky130_fd_sc_hd__or2_1
X_05759_ _05871_/A vssd1 vssd1 vccd1 vccd1 _05759_/X sky130_fd_sc_hd__buf_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ _10060_/Q _08478_/B vssd1 vssd1 vccd1 vccd1 _08479_/B sky130_fd_sc_hd__or2_2
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07429_ _10273_/Q _07429_/B vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__or2_1
X_10440_ _10442_/CLK _10440_/D vssd1 vssd1 vccd1 vccd1 _10440_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10436_/CLK _10371_/D vssd1 vssd1 vccd1 vccd1 _10371_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10450_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06800_ _06802_/A _06800_/B vssd1 vssd1 vccd1 vccd1 _06800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07780_ _05966_/X _07516_/B _07913_/A vssd1 vssd1 vccd1 vccd1 _07780_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 io_pwm_test vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
X_06731_ _10356_/Q _06668_/B _06669_/B vssd1 vssd1 vccd1 vccd1 _06792_/B sky130_fd_sc_hd__a21boi_4
XFILLER_209_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09450_ _09446_/X _09449_/X _09446_/X _09449_/X vssd1 vssd1 vccd1 vccd1 _09450_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06662_ _05018_/X _06653_/Y _06656_/Y _06661_/X vssd1 vssd1 vccd1 vccd1 _06662_/X
+ sky130_fd_sc_hd__o22a_1
X_08401_ _08401_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06593_ _06590_/X _06592_/X _06590_/X _06592_/X vssd1 vssd1 vccd1 vccd1 _06593_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_09381_ _09381_/A _09380_/X vssd1 vssd1 vccd1 vccd1 _09381_/X sky130_fd_sc_hd__or2b_1
X_05613_ _09913_/X _05612_/Y _09913_/X _05612_/Y vssd1 vssd1 vccd1 vccd1 _05614_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_08332_ _09029_/A vssd1 vssd1 vccd1 vccd1 _09174_/A sky130_fd_sc_hd__buf_1
X_05544_ _05542_/Y _05543_/Y _05542_/Y _05543_/Y vssd1 vssd1 vccd1 vccd1 _05544_/X
+ sky130_fd_sc_hd__a2bb2o_4
X_08263_ _08265_/A _08257_/Y _06263_/B vssd1 vssd1 vccd1 vccd1 _08263_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05475_ _05475_/A _05475_/B vssd1 vssd1 vccd1 vccd1 _05475_/Y sky130_fd_sc_hd__nor2_1
X_07214_ _07218_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07214_/X sky130_fd_sc_hd__or2_1
X_08194_ _08116_/X _08191_/B _08192_/Y _08193_/X vssd1 vssd1 vccd1 vccd1 _08194_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07145_ _07145_/A _07144_/X vssd1 vssd1 vccd1 vccd1 _07145_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07076_ _07056_/A _07082_/B _07050_/A vssd1 vssd1 vccd1 vccd1 _07077_/B sky130_fd_sc_hd__a21oi_1
X_06027_ _09845_/X _06015_/X _06026_/X _06017_/X _06018_/X vssd1 vssd1 vccd1 vccd1
+ _10198_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07978_ _07501_/X _07506_/X _07507_/X _07530_/X _07476_/X vssd1 vssd1 vccd1 vccd1
+ _07978_/X sky130_fd_sc_hd__o221a_1
XFILLER_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09717_ _10450_/Q _06736_/X _09717_/S vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06929_ _07021_/B vssd1 vssd1 vccd1 vccd1 _06929_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _10114_/Q input44/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _08411_/Y _10125_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09579_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10423_ _10426_/CLK _10423_/D vssd1 vssd1 vccd1 vccd1 _10423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _10421_/CLK _10354_/D vssd1 vssd1 vccd1 vccd1 _10354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10285_ _10297_/CLK _10285_/D vssd1 vssd1 vccd1 vccd1 _10285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05260_ input49/X _05251_/X _08761_/A _05252_/X _05253_/X vssd1 vssd1 vccd1 vccd1
+ _10355_/D sky130_fd_sc_hd__a221o_1
XFILLER_162_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05191_ _05185_/X _10391_/Q _05186_/X _09610_/X _05189_/X vssd1 vssd1 vccd1 vccd1
+ _10391_/D sky130_fd_sc_hd__o221a_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__or2_1
XFILLER_142_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08881_ _09968_/X vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__inv_2
X_07901_ _07804_/X _07900_/X _07804_/X _07900_/X vssd1 vssd1 vccd1 vccd1 _07903_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07832_ _07837_/A _09915_/X _07813_/C _07837_/B vssd1 vssd1 vccd1 vccd1 _07833_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09502_ _08409_/X _06397_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__mux2_1
X_07763_ _07773_/A vssd1 vssd1 vccd1 vccd1 _07916_/C sky130_fd_sc_hd__buf_1
X_06714_ _10366_/Q vssd1 vssd1 vccd1 vccd1 _06714_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07694_ _07694_/A _07700_/A vssd1 vssd1 vccd1 vccd1 _07694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ _09429_/X _09432_/Y _09429_/X _09432_/Y vssd1 vssd1 vccd1 vccd1 _09434_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_06645_ _08626_/A _10348_/Q vssd1 vssd1 vccd1 vccd1 _06645_/Y sky130_fd_sc_hd__nor2_4
XFILLER_197_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ _09462_/C vssd1 vssd1 vccd1 vccd1 _09428_/C sky130_fd_sc_hd__inv_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06576_ _10105_/Q _06466_/A _06570_/X _06572_/Y vssd1 vssd1 vccd1 vccd1 _06576_/X
+ sky130_fd_sc_hd__a22o_1
X_08315_ _08315_/A vssd1 vssd1 vccd1 vccd1 _09997_/S sky130_fd_sc_hd__clkinv_8
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ _09295_/A vssd1 vssd1 vccd1 vccd1 _09295_/Y sky130_fd_sc_hd__inv_2
X_05527_ _10016_/X _10008_/X _05478_/Y _05546_/A vssd1 vssd1 vccd1 vccd1 _05542_/A
+ sky130_fd_sc_hd__o22a_1
X_08246_ _10192_/Q _08242_/Y _08219_/X _08249_/B vssd1 vssd1 vccd1 vccd1 _08246_/X
+ sky130_fd_sc_hd__o211a_1
X_05458_ _10317_/Q vssd1 vssd1 vccd1 vccd1 _05458_/Y sky130_fd_sc_hd__inv_2
X_08177_ _08176_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__nand2b_4
XFILLER_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05389_ _05389_/A _05435_/A vssd1 vssd1 vccd1 vccd1 _05431_/A sky130_fd_sc_hd__or2_1
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07128_ _07118_/C _07127_/A _07117_/A _07127_/Y vssd1 vssd1 vccd1 vccd1 _07128_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07059_ _07223_/A _07072_/B vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__or2_1
X_10070_ _10202_/CLK _10070_/D vssd1 vssd1 vccd1 vccd1 _10070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10406_ _10442_/CLK _10406_/D vssd1 vssd1 vccd1 vccd1 _10406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ _10343_/CLK _10337_/D vssd1 vssd1 vccd1 vccd1 _10337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10268_ _10298_/CLK _10268_/D vssd1 vssd1 vccd1 vccd1 _10268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _10202_/CLK _10199_/D vssd1 vssd1 vccd1 vccd1 _10199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10420_/CLK sky130_fd_sc_hd__clkbuf_16
X_06430_ _06430_/A vssd1 vssd1 vccd1 vccd1 _06487_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06361_ _10244_/Q _08390_/A _06360_/Y _10137_/Q vssd1 vssd1 vccd1 vccd1 _06362_/A
+ sky130_fd_sc_hd__o22a_2
X_08100_ _06628_/Y _10202_/Q _06621_/A _08077_/X vssd1 vssd1 vccd1 vccd1 _08100_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05312_ _05312_/A _05312_/B vssd1 vssd1 vccd1 vccd1 _05313_/B sky130_fd_sc_hd__nand2_1
X_09080_ _09174_/A _09247_/A _09000_/X vssd1 vssd1 vccd1 vccd1 _09080_/X sky130_fd_sc_hd__or3b_1
X_06292_ _10237_/Q vssd1 vssd1 vccd1 vccd1 _06293_/A sky130_fd_sc_hd__inv_2
Xinput40 io_wb_dat_i[29] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_4
X_05243_ _10363_/Q _05239_/X input26/X _05240_/X _05236_/X vssd1 vssd1 vccd1 vccd1
+ _10363_/D sky130_fd_sc_hd__o221a_1
X_08031_ _07412_/A _07412_/B _07413_/B vssd1 vssd1 vccd1 vccd1 _08031_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput51 io_wb_we_i vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
X_05174_ _05153_/X _05172_/Y _05173_/Y _05161_/X vssd1 vssd1 vccd1 vccd1 _05175_/B
+ sky130_fd_sc_hd__o22a_1
X_09982_ _09981_/X _06630_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08933_ _09069_/A _09986_/X vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__or2_2
XFILLER_130_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _10289_/Q _05801_/X _08851_/X _08863_/X vssd1 vssd1 vccd1 vccd1 _08864_/X
+ sky130_fd_sc_hd__o22a_1
X_08795_ _06072_/X _08775_/Y _08782_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _08819_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07815_ _07815_/A _09914_/X vssd1 vssd1 vccd1 vccd1 _07815_/X sky130_fd_sc_hd__or2_1
X_07746_ _07644_/A _07644_/B _07644_/X vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__a21bo_1
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _09474_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09416_/X sky130_fd_sc_hd__or2_1
X_07677_ _07677_/A vssd1 vssd1 vccd1 vccd1 _07777_/C sky130_fd_sc_hd__clkbuf_2
X_06628_ _10373_/Q vssd1 vssd1 vccd1 vccd1 _06628_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06559_ _10103_/Q _06465_/A _08436_/A _06435_/A vssd1 vssd1 vccd1 vccd1 _06563_/A
+ sky130_fd_sc_hd__a22o_1
X_09347_ _09345_/X _09346_/X _09345_/X _09346_/X vssd1 vssd1 vccd1 vccd1 _09347_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _08843_/X _08869_/X _08843_/X _08869_/X vssd1 vssd1 vccd1 vccd1 _09279_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08229_ _06254_/A _08225_/Y _08219_/X _08232_/B vssd1 vssd1 vccd1 vccd1 _08229_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10122_ _10244_/CLK _10122_/D vssd1 vssd1 vccd1 vccd1 _10122_/Q sky130_fd_sc_hd__dfxtp_1
X_10053_ _10178_/CLK _10053_/D vssd1 vssd1 vccd1 vccd1 _10053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05930_ _10232_/Q _05927_/X _05091_/X _05928_/X _05918_/X vssd1 vssd1 vccd1 vccd1
+ _10232_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05861_ _05861_/A vssd1 vssd1 vccd1 vccd1 _06834_/A sky130_fd_sc_hd__inv_2
X_08580_ _08587_/A _08580_/B _08580_/C vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__and3_1
XFILLER_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07600_ _07585_/X _07587_/X _07598_/X _07599_/X vssd1 vssd1 vccd1 vccd1 _07600_/X
+ sky130_fd_sc_hd__o22a_1
X_07531_ _07507_/X _07530_/X _07507_/X _07530_/X vssd1 vssd1 vccd1 vccd1 _07761_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05792_ _10259_/Q vssd1 vssd1 vccd1 vccd1 _05792_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07462_ _07686_/B vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_210_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09201_ _09252_/A _09258_/B _09201_/C vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__or3_4
X_07393_ _07393_/A vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__inv_2
X_06413_ _06836_/A vssd1 vssd1 vccd1 vccd1 _06413_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09132_ _09292_/A _09949_/X _09038_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09132_/X
+ sky130_fd_sc_hd__o22a_1
X_06344_ _06344_/A _06344_/B vssd1 vssd1 vccd1 vccd1 _06345_/A sky130_fd_sc_hd__or2_2
XFILLER_175_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__or2_1
X_06275_ _10235_/Q vssd1 vssd1 vccd1 vccd1 _06275_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05226_ _10373_/Q _05221_/X input37/X _05223_/X _05218_/X vssd1 vssd1 vccd1 vccd1
+ _10373_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08014_ _08014_/A vssd1 vssd1 vccd1 vccd1 _08015_/B sky130_fd_sc_hd__inv_2
X_05157_ _05157_/A _05157_/B vssd1 vssd1 vccd1 vccd1 _10401_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09965_ _09964_/X _10374_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09965_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05088_ input49/X _05082_/X _10419_/Q _05083_/X _05086_/X vssd1 vssd1 vccd1 vccd1
+ _10419_/D sky130_fd_sc_hd__a221o_1
XFILLER_134_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08916_ _08939_/A _09985_/X vssd1 vssd1 vccd1 vccd1 _08916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09896_ _06859_/X _05837_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09896_/X sky130_fd_sc_hd__mux2_2
X_08847_ _10292_/Q _08847_/B vssd1 vssd1 vccd1 vccd1 _08847_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _08624_/A _08624_/B _08624_/Y vssd1 vssd1 vccd1 vccd1 _08778_/X sky130_fd_sc_hd__a21o_1
XFILLER_150_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07729_ _07725_/X _07726_/X _07725_/X _07726_/X vssd1 vssd1 vccd1 vccd1 _07729_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10105_ _10207_/CLK _10105_/D vssd1 vssd1 vccd1 vccd1 _10105_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10036_ _10176_/CLK _10036_/D vssd1 vssd1 vccd1 vccd1 _10036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06060_ _09797_/X _06054_/X _08801_/A _06056_/X _06057_/X vssd1 vssd1 vccd1 vccd1
+ _10186_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05011_ _05013_/A vssd1 vssd1 vccd1 vccd1 _05012_/A sky130_fd_sc_hd__inv_2
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ _09749_/X _10226_/Q _09998_/S vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__mux2_1
X_06962_ _06962_/A _09894_/X vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__or2_1
X_08701_ _08138_/X _10049_/Q _08116_/X _08456_/X _08656_/X vssd1 vssd1 vccd1 vccd1
+ _08704_/B sky130_fd_sc_hd__a221o_1
X_09681_ _06440_/X input44/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05913_ _10240_/Q _05910_/X _05091_/X _05911_/X _05908_/X vssd1 vssd1 vccd1 vccd1
+ _10240_/D sky130_fd_sc_hd__o221a_1
X_08632_ _08632_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06893_ _06931_/A _09668_/X vssd1 vssd1 vccd1 vccd1 _06894_/C sky130_fd_sc_hd__or2_2
X_05844_ _05827_/X _05843_/X _05827_/X _05843_/X vssd1 vssd1 vccd1 vccd1 _06855_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_08563_ _08783_/A _08562_/X _08554_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _08591_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05775_ _05775_/A input11/X input12/X vssd1 vssd1 vccd1 vccd1 _06137_/A sky130_fd_sc_hd__or3b_1
XFILLER_207_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08494_ _10075_/Q _08494_/B vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__or2_1
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07514_ _07496_/X _07498_/X _07496_/X _07498_/X vssd1 vssd1 vccd1 vccd1 _07514_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07445_ _07445_/A vssd1 vssd1 vccd1 vccd1 _07445_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _06993_/B _07356_/X _06993_/B _07356_/X vssd1 vssd1 vccd1 vccd1 _07393_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09115_ _08866_/Y _09114_/X _08866_/Y _09114_/X vssd1 vssd1 vccd1 vccd1 _09117_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_06327_ _06327_/A vssd1 vssd1 vccd1 vccd1 _06327_/Y sky130_fd_sc_hd__inv_2
X_06258_ _10192_/Q _08238_/A vssd1 vssd1 vccd1 vccd1 _06259_/B sky130_fd_sc_hd__or2_1
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09046_ _09043_/Y _09044_/Y _09045_/X vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__o21ai_1
XFILLER_135_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05209_ _05202_/X _10380_/Q _05203_/X _09747_/X _05206_/X vssd1 vssd1 vccd1 vccd1
+ _10380_/D sky130_fd_sc_hd__o221a_1
XFILLER_150_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06189_ _06225_/A vssd1 vssd1 vccd1 vccd1 _06204_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _08990_/X _08988_/A _09986_/S vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_20 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _10378_/Q _09878_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10019_ _08006_/A _08038_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05560_ _05558_/Y _05559_/Y _05558_/Y _05559_/Y vssd1 vssd1 vccd1 vccd1 _05560_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05491_ _10014_/X _10017_/X _10014_/X _10017_/X vssd1 vssd1 vccd1 vccd1 _05491_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07230_ _07213_/A _07213_/B _07213_/Y vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__o21ai_1
XFILLER_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _07161_/A _07223_/B _07161_/C vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__or3_1
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06112_ _10158_/Q _05891_/X _10330_/Q _05761_/X _06111_/X vssd1 vssd1 vccd1 vccd1
+ _10158_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07092_ _07068_/C _07065_/B _07065_/Y vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06043_ _06067_/A vssd1 vssd1 vccd1 vccd1 _06043_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09802_ _08227_/Y _10359_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09802_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07994_ _07745_/X _07747_/X _07745_/X _07747_/X vssd1 vssd1 vccd1 vccd1 _08011_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09733_ _06805_/Y _10398_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10064_/D sky130_fd_sc_hd__mux2_1
X_06945_ _06945_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _06946_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09664_ _10146_/Q _10162_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__mux2_1
X_06876_ _07068_/A vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08615_ _08616_/A _08616_/B _08614_/X vssd1 vssd1 vccd1 vccd1 _08617_/A sky130_fd_sc_hd__o21ai_1
X_09595_ _08443_/Y _08442_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09595_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05827_ _07437_/A _10261_/Q _05787_/Y _05826_/Y vssd1 vssd1 vccd1 vccd1 _05827_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _10053_/Q _08471_/B _08472_/B vssd1 vssd1 vccd1 vccd1 _08547_/B sky130_fd_sc_hd__a21bo_1
X_05758_ _05800_/A _05751_/X _09635_/X _05753_/X _05756_/X vssd1 vssd1 vccd1 vccd1
+ _10273_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08477_ _10059_/Q _08477_/B vssd1 vssd1 vccd1 vccd1 _08478_/B sky130_fd_sc_hd__or2_1
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05689_ _05689_/A vssd1 vssd1 vccd1 vccd1 _05689_/Y sky130_fd_sc_hd__inv_2
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07428_ _10272_/Q _07428_/B vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__or2_1
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07359_ _07347_/X _07352_/X _07353_/X _07358_/X vssd1 vssd1 vccd1 vccd1 _07359_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10370_ _10436_/CLK _10370_/D vssd1 vssd1 vccd1 vccd1 _10370_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09029_ _09029_/A _09948_/X vssd1 vssd1 vccd1 vccd1 _09029_/X sky130_fd_sc_hd__or2_1
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 io_sync_in vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
X_06730_ _10357_/Q _06669_/B _06670_/B vssd1 vssd1 vccd1 vccd1 _06793_/B sky130_fd_sc_hd__a21bo_1
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ _05024_/A _06657_/Y _06645_/Y _06660_/Y vssd1 vssd1 vccd1 vccd1 _06661_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05612_ _09907_/X _05536_/X _05620_/A vssd1 vssd1 vccd1 vccd1 _05612_/Y sky130_fd_sc_hd__o21ai_1
X_08400_ _09495_/X _08435_/B vssd1 vssd1 vccd1 vccd1 _08400_/X sky130_fd_sc_hd__and2_1
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06592_ _08446_/A _06489_/A _08448_/A _06437_/A _06591_/X vssd1 vssd1 vccd1 vccd1
+ _06592_/X sky130_fd_sc_hd__o221a_1
X_09380_ _09380_/A _09380_/B vssd1 vssd1 vccd1 vccd1 _09380_/X sky130_fd_sc_hd__or2_1
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08939_/A vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__buf_1
X_05543_ _05475_/A _05475_/B _05475_/Y vssd1 vssd1 vccd1 vccd1 _05543_/Y sky130_fd_sc_hd__a21oi_2
X_08262_ _08260_/A _08260_/B _08240_/X _08261_/Y vssd1 vssd1 vccd1 vccd1 _08262_/Y
+ sky130_fd_sc_hd__a211oi_2
X_05474_ _10020_/X vssd1 vssd1 vccd1 vccd1 _05475_/B sky130_fd_sc_hd__inv_2
XFILLER_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07213_ _07213_/A _07213_/B vssd1 vssd1 vccd1 vccd1 _07213_/Y sky130_fd_sc_hd__nand2_1
X_08193_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08193_/X sky130_fd_sc_hd__buf_6
XFILLER_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07144_ _07146_/A _09884_/X _07161_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07144_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07075_ _07071_/X _07074_/X _07071_/X _07074_/X vssd1 vssd1 vccd1 vccd1 _07075_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06026_ _08504_/A vssd1 vssd1 vccd1 vccd1 _06026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07977_ _07931_/X _07932_/X _07930_/X _07933_/X vssd1 vssd1 vccd1 vccd1 _07977_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09716_ _09715_/X _10382_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10048_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06928_ _09895_/X vssd1 vssd1 vccd1 vccd1 _07021_/B sky130_fd_sc_hd__buf_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09647_ _10113_/Q input41/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09647_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06859_ _07023_/A _07023_/B _07023_/A _07023_/B vssd1 vssd1 vccd1 vccd1 _06859_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _08408_/Y _09577_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09578_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _10060_/Q _08478_/B _08479_/B vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__a21bo_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10422_ _10422_/CLK _10422_/D vssd1 vssd1 vccd1 vccd1 _10422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10353_ _10414_/CLK _10353_/D vssd1 vssd1 vccd1 vccd1 _10353_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10284_ _10297_/CLK _10284_/D vssd1 vssd1 vccd1 vccd1 _10284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05190_ _05185_/X _10392_/Q _05186_/X _09611_/X _05189_/X vssd1 vssd1 vccd1 vccd1
+ _10392_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08880_ _09042_/B _08876_/X _08895_/B vssd1 vssd1 vccd1 vccd1 _08880_/Y sky130_fd_sc_hd__o21ai_1
X_07900_ _07861_/Y _07899_/X _07861_/Y _07899_/X vssd1 vssd1 vccd1 vccd1 _07900_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07831_ _07827_/X _07830_/X _07827_/X _07830_/X vssd1 vssd1 vccd1 vccd1 _07831_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09501_ _09500_/X _06638_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07762_ _07777_/C vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__inv_2
X_06713_ _06713_/A vssd1 vssd1 vccd1 vccd1 _06806_/B sky130_fd_sc_hd__inv_2
XFILLER_112_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07693_ _07679_/A _07688_/Y _07685_/X _07689_/X vssd1 vssd1 vccd1 vccd1 _07700_/A
+ sky130_fd_sc_hd__o22ai_4
X_09432_ _09432_/A vssd1 vssd1 vccd1 vccd1 _09432_/Y sky130_fd_sc_hd__inv_2
X_06644_ _08763_/A vssd1 vssd1 vccd1 vccd1 _06644_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06575_ _10106_/Q _06465_/A _08444_/A _06435_/A vssd1 vssd1 vccd1 vccd1 _06580_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09363_ _09309_/X _09322_/Y _09323_/X _09324_/X vssd1 vssd1 vccd1 vccd1 _09375_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08314_ _06273_/A _08313_/Y _08616_/A _08313_/A _08188_/X vssd1 vssd1 vccd1 vccd1
+ _08314_/X sky130_fd_sc_hd__o221a_1
X_05526_ _10019_/X _10013_/X _05481_/Y _05550_/A vssd1 vssd1 vccd1 vccd1 _05546_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09294_ _09294_/A _09294_/B _09294_/C vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__and3_1
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08249_/B sky130_fd_sc_hd__or2_2
XFILLER_165_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05457_ _10315_/Q vssd1 vssd1 vccd1 vccd1 _05457_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _08176_/A _08176_/B _08176_/C _08176_/D vssd1 vssd1 vccd1 vccd1 _08176_/X
+ sky130_fd_sc_hd__and4_1
X_05388_ _05388_/A _05440_/A vssd1 vssd1 vccd1 vccd1 _05435_/A sky130_fd_sc_hd__or2_1
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07127_ _07127_/A vssd1 vssd1 vccd1 vccd1 _07127_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07058_ _07063_/A _09887_/X vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__or2_1
X_06009_ _10205_/Q vssd1 vssd1 vccd1 vccd1 _06271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10244_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10405_ _10437_/CLK _10405_/D vssd1 vssd1 vccd1 vccd1 _10405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10336_ _10346_/CLK _10336_/D vssd1 vssd1 vccd1 vccd1 _10336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10267_ _10300_/CLK _10267_/D vssd1 vssd1 vccd1 vccd1 _10267_/Q sky130_fd_sc_hd__dfxtp_1
X_10198_ _10202_/CLK _10198_/D vssd1 vssd1 vccd1 vccd1 _10198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06360_ _10244_/Q vssd1 vssd1 vccd1 vccd1 _06360_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05311_ _05311_/A vssd1 vssd1 vccd1 vccd1 _05312_/B sky130_fd_sc_hd__inv_2
X_06291_ _10237_/Q _08349_/A vssd1 vssd1 vccd1 vccd1 _06294_/A sky130_fd_sc_hd__nor2_1
X_05242_ _10364_/Q _05239_/X input27/X _05240_/X _05236_/X vssd1 vssd1 vccd1 vccd1
+ _10364_/D sky130_fd_sc_hd__o221a_1
Xinput30 io_wb_dat_i[1] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_4
X_08030_ _08027_/A _08027_/B _08027_/Y vssd1 vssd1 vccd1 vccd1 _08030_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput41 io_wb_dat_i[2] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_6
Xinput52 reset vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_4
X_05173_ _10429_/Q vssd1 vssd1 vccd1 vccd1 _05173_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _06615_/D _08169_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__mux2_1
X_08932_ _09070_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__or2_2
XFILLER_96_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ _08852_/Y _08862_/Y _10288_/Q _08852_/B vssd1 vssd1 vccd1 vccd1 _08863_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08794_ _08815_/A _08815_/B _08794_/C vssd1 vssd1 vccd1 vccd1 _08794_/X sky130_fd_sc_hd__or3_1
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07814_ _07814_/A _09917_/X vssd1 vssd1 vccd1 vccd1 _07814_/X sky130_fd_sc_hd__or2_1
XFILLER_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07745_ _07742_/X _07744_/X _07742_/X _07744_/X vssd1 vssd1 vccd1 vccd1 _07745_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09415_ _09245_/B _09225_/X _09170_/C vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__o21a_1
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07773_/A sky130_fd_sc_hd__or2_2
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06627_ _10375_/Q vssd1 vssd1 vccd1 vccd1 _06627_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06558_ _10103_/Q vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__inv_2
X_09346_ _09173_/X _09298_/A _09300_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09346_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06489_ _06489_/A vssd1 vssd1 vccd1 vccd1 _06489_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _09276_/A _09276_/B _09332_/A vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__a21bo_1
X_05509_ _07218_/B vssd1 vssd1 vccd1 vccd1 _07234_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_193_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08228_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__or2_2
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08159_ _10187_/Q vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__inv_2
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10121_ _10244_/CLK _10121_/D vssd1 vssd1 vccd1 vccd1 _10121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _10421_/CLK _10052_/D vssd1 vssd1 vccd1 vccd1 _10052_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10319_ _10343_/CLK _10319_/D vssd1 vssd1 vccd1 vccd1 _10319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05860_ _05796_/X _05821_/X _05796_/X _05821_/X vssd1 vssd1 vccd1 vccd1 _05861_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05791_ _05791_/A vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__buf_2
XFILLER_207_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07530_ _07524_/A _07707_/A _07523_/Y _07521_/A _07529_/Y vssd1 vssd1 vccd1 vccd1
+ _07530_/X sky130_fd_sc_hd__o32a_1
XFILLER_207_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07461_ _10216_/Q vssd1 vssd1 vccd1 vccd1 _07686_/B sky130_fd_sc_hd__inv_2
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ _09354_/A _09417_/A vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__or2_2
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06412_ _06821_/A vssd1 vssd1 vccd1 vccd1 _06412_/Y sky130_fd_sc_hd__inv_2
X_07392_ _07392_/A vssd1 vssd1 vccd1 vccd1 _07408_/A sky130_fd_sc_hd__inv_2
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09131_ _05931_/X _09418_/B _09201_/C _09130_/X vssd1 vssd1 vccd1 vccd1 _09131_/X
+ sky130_fd_sc_hd__a31o_1
X_06343_ _06343_/A vssd1 vssd1 vccd1 vccd1 _06344_/B sky130_fd_sc_hd__inv_2
XFILLER_175_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _09063_/B vssd1 vssd1 vccd1 vccd1 _09062_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06274_ _10128_/Q vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__inv_2
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05225_ _10374_/Q _05221_/X input38/X _05223_/X _05218_/X vssd1 vssd1 vccd1 vccd1
+ _10374_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08013_ _07425_/A _07878_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__o21ai_1
X_05156_ _05153_/X _06616_/B _05155_/Y _05138_/X vssd1 vssd1 vccd1 vccd1 _05157_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09964_ _10406_/Q _10203_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05087_ input50/X _05082_/X _10420_/Q _05083_/X _05086_/X vssd1 vssd1 vccd1 vccd1
+ _10420_/D sky130_fd_sc_hd__a221o_1
XFILLER_103_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08915_ _08915_/A _09977_/X vssd1 vssd1 vccd1 vccd1 _08915_/X sky130_fd_sc_hd__or2_1
X_09895_ _06858_/X _06414_/Y _10022_/S vssd1 vssd1 vccd1 vccd1 _09895_/X sky130_fd_sc_hd__mux2_1
X_08846_ _10293_/Q _05852_/X _10293_/Q _05852_/X vssd1 vssd1 vccd1 vccd1 _08846_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08777_ _06072_/X _08775_/Y _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08817_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05989_ _10445_/Q _06126_/A vssd1 vssd1 vccd1 vccd1 _05989_/X sky130_fd_sc_hd__and2_1
XFILLER_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07728_ _07717_/X _07727_/X _07717_/X _07727_/X vssd1 vssd1 vccd1 vccd1 _07728_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07659_ _07910_/A _07658_/B _07658_/Y vssd1 vssd1 vccd1 vccd1 _07659_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09329_ _09271_/X _09272_/X _09224_/X _09273_/X vssd1 vssd1 vccd1 vccd1 _09329_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10422_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10207_/CLK _10104_/D vssd1 vssd1 vccd1 vccd1 _10104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10035_ _10205_/CLK _10035_/D vssd1 vssd1 vccd1 vccd1 _10036_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_191_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05010_ _06083_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _05013_/A sky130_fd_sc_hd__or2_2
XFILLER_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06961_ _06961_/A _09896_/X vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__nor2_1
X_08700_ _06000_/A _08613_/Y _08695_/A _08699_/X vssd1 vssd1 vccd1 vccd1 _08700_/X
+ sky130_fd_sc_hd__o22a_1
X_09680_ _06426_/X input41/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09680_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05912_ _10241_/Q _05910_/X _05089_/X _05911_/X _05908_/X vssd1 vssd1 vccd1 vccd1
+ _10241_/D sky130_fd_sc_hd__o221a_1
X_08631_ _06606_/X _06653_/Y _08624_/Y _08630_/X vssd1 vssd1 vccd1 vccd1 _08632_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06892_ _09893_/X vssd1 vssd1 vccd1 vccd1 _06912_/B sky130_fd_sc_hd__inv_2
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05843_ _05786_/A _10262_/Q _05786_/Y vssd1 vssd1 vccd1 vccd1 _05843_/X sky130_fd_sc_hd__a21o_1
X_08562_ _08465_/X _08561_/X _08465_/X _08561_/X vssd1 vssd1 vccd1 vccd1 _08562_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_05774_ _08324_/A _05923_/B vssd1 vssd1 vccd1 vccd1 _05944_/B sky130_fd_sc_hd__or2_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08493_ _08494_/B vssd1 vssd1 vccd1 vccd1 _08493_/Y sky130_fd_sc_hd__inv_2
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07513_ _07513_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _07524_/A sky130_fd_sc_hd__or2_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07444_ _05788_/A _07440_/B _07441_/B vssd1 vssd1 vccd1 vccd1 _07444_/X sky130_fd_sc_hd__a21bo_1
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07375_ _07353_/X _07358_/X _07353_/X _07358_/X vssd1 vssd1 vccd1 vccd1 _07390_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09114_ _10292_/Q _08847_/B _08847_/Y vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__a21o_1
X_06326_ _10239_/Q _08363_/A _06312_/B _06317_/X vssd1 vssd1 vccd1 vccd1 _06327_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06257_ _10191_/Q _06257_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__or2_1
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09045_ _09258_/A _09045_/B _09091_/C vssd1 vssd1 vccd1 vccd1 _09045_/X sky130_fd_sc_hd__or3_4
X_05208_ _05202_/X _10381_/Q _05203_/X _09491_/X _05206_/X vssd1 vssd1 vccd1 vccd1
+ _10381_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06188_ _06224_/A vssd1 vssd1 vccd1 vccd1 _06225_/A sky130_fd_sc_hd__inv_2
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05139_ _05129_/X _06615_/B _05137_/Y _05138_/X vssd1 vssd1 vccd1 vccd1 _05140_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09947_ _09113_/X _09111_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09947_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_10 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _08311_/X _10378_/Q _09878_/S vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__mux2_1
XINSDIODE2_21 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08829_ _08273_/A _08726_/Y _08600_/A _08723_/Y _08828_/Y vssd1 vssd1 vccd1 vccd1
+ _08829_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _08002_/A _08030_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10018_/X sky130_fd_sc_hd__mux2_2
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05490_ _10012_/X _09990_/X _10012_/X _09990_/X vssd1 vssd1 vccd1 vccd1 _05490_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07160_ _07160_/A vssd1 vssd1 vccd1 vccd1 _07161_/C sky130_fd_sc_hd__inv_2
XFILLER_172_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06111_ _06111_/A vssd1 vssd1 vccd1 vccd1 _06111_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07091_ _07079_/A _07079_/B _07253_/A vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__a21o_1
X_06042_ _09825_/X _06028_/X _10193_/Q _06031_/X _06032_/X vssd1 vssd1 vccd1 vccd1
+ _10193_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09800_/X input21/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09732_ _06804_/Y _10397_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10063_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07993_ _07741_/X _07748_/X _07741_/X _07748_/X vssd1 vssd1 vccd1 vccd1 _08010_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06944_ _06919_/A _06925_/A _06919_/Y vssd1 vssd1 vccd1 vccd1 _06944_/X sky130_fd_sc_hd__a21o_1
X_09663_ _10145_/Q _10161_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06875_ _07223_/A vssd1 vssd1 vccd1 vccd1 _07068_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ _08454_/Y _08493_/Y _08613_/Y _10076_/Q _08494_/X vssd1 vssd1 vccd1 vccd1
+ _08614_/X sky130_fd_sc_hd__a32o_1
X_09594_ _08440_/Y _08439_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05826_ _05826_/A vssd1 vssd1 vccd1 vccd1 _05826_/Y sky130_fd_sc_hd__inv_2
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08545_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05757_ _08850_/B _05751_/X _09636_/X _05753_/X _05756_/X vssd1 vssd1 vccd1 vccd1
+ _10274_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08476_ _10058_/Q _08476_/B vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__or2_1
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05688_ _08618_/A _05688_/B vssd1 vssd1 vccd1 vccd1 _10301_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07427_ _10271_/Q _07427_/B vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__or2_1
XFILLER_195_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _07358_/A _07358_/B vssd1 vssd1 vccd1 vccd1 _07358_/X sky130_fd_sc_hd__or2_1
XFILLER_50_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06309_ _10239_/Q _08363_/A vssd1 vssd1 vccd1 vccd1 _06312_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07289_ _06866_/A _07235_/B _07068_/A _06824_/X vssd1 vssd1 vccd1 vccd1 _07289_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _09949_/X vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__inv_2
XFILLER_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 io_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06660_ _06660_/A vssd1 vssd1 vccd1 vccd1 _06660_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05611_ _05621_/A _05621_/B vssd1 vssd1 vccd1 vccd1 _05620_/A sky130_fd_sc_hd__nand2_1
X_06591_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06591_/X sky130_fd_sc_hd__or2_1
X_08330_ _10227_/Q vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__inv_2
X_05542_ _05542_/A vssd1 vssd1 vccd1 vccd1 _05542_/Y sky130_fd_sc_hd__inv_2
X_08261_ _08265_/B vssd1 vssd1 vccd1 vccd1 _08261_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05473_ _10010_/X vssd1 vssd1 vccd1 vccd1 _05475_/A sky130_fd_sc_hd__inv_2
X_07212_ _07212_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07213_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08192_ _08196_/B vssd1 vssd1 vccd1 vccd1 _08192_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07143_ _07146_/A _09884_/X _07146_/C _07217_/B vssd1 vssd1 vccd1 vccd1 _07145_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07074_ _07074_/A _07074_/B vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__or2_1
X_06025_ _10198_/Q vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07976_ _07934_/X _07939_/X _07940_/X _07975_/X vssd1 vssd1 vccd1 vccd1 _07976_/Y
+ sky130_fd_sc_hd__o22ai_1
X_09715_ _10449_/Q _06740_/A _09717_/S vssd1 vssd1 vccd1 vccd1 _09715_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06927_ _06905_/X _06926_/X _06905_/X _06926_/X vssd1 vssd1 vccd1 vccd1 _06927_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09646_ _10112_/Q input30/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09646_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06858_ _06855_/A _06855_/B _06856_/B vssd1 vssd1 vccd1 vccd1 _06858_/X sky130_fd_sc_hd__a21bo_1
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06789_ _09717_/S _06789_/B vssd1 vssd1 vccd1 vccd1 _06789_/X sky130_fd_sc_hd__and2_1
X_09577_ _08406_/Y _09576_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09577_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05809_ _10254_/Q vssd1 vssd1 vccd1 vccd1 _05809_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08528_ _08809_/A _08519_/X _08520_/Y vssd1 vssd1 vccd1 vccd1 _08596_/B sky130_fd_sc_hd__o21ai_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _08459_/A _10047_/Q vssd1 vssd1 vccd1 vccd1 _08459_/Y sky130_fd_sc_hd__nor2_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10421_ _10421_/CLK _10421_/D vssd1 vssd1 vccd1 vccd1 _10421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10352_ _10414_/CLK _10352_/D vssd1 vssd1 vccd1 vccd1 _10352_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_164_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10283_ _10297_/CLK _10283_/D vssd1 vssd1 vccd1 vccd1 _10283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07830_ _07830_/A _07897_/B _07830_/C vssd1 vssd1 vccd1 vccd1 _07830_/X sky130_fd_sc_hd__or3_1
XFILLER_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07906_/A sky130_fd_sc_hd__or2_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06712_ _06633_/A _08729_/A _08727_/A vssd1 vssd1 vccd1 vccd1 _06713_/A sky130_fd_sc_hd__a21bo_1
X_09500_ _06637_/Y _08166_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07692_ _07692_/A vssd1 vssd1 vccd1 vccd1 _07694_/A sky130_fd_sc_hd__inv_2
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _09320_/A _09321_/A _09373_/Y _09370_/Y _09430_/X vssd1 vssd1 vccd1 vccd1
+ _09432_/A sky130_fd_sc_hd__a32o_1
X_06643_ _10389_/Q vssd1 vssd1 vccd1 vccd1 _06643_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06574_ _10106_/Q vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__inv_2
X_09362_ _09360_/X _09361_/X _09360_/X _09361_/X vssd1 vssd1 vccd1 vccd1 _09362_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08313_ _08313_/A vssd1 vssd1 vccd1 vccd1 _08313_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05525_ _10023_/X _10022_/X _05482_/X _05524_/X vssd1 vssd1 vccd1 vccd1 _05550_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _09343_/C vssd1 vssd1 vccd1 vccd1 _09390_/C sky130_fd_sc_hd__inv_2
XFILLER_20_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08244_ _08172_/X _08238_/Y _06259_/B vssd1 vssd1 vccd1 vccd1 _08244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_165_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05456_ _10316_/Q vssd1 vssd1 vccd1 vccd1 _05456_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _08175_/A _08175_/B _08175_/C _08175_/D vssd1 vssd1 vccd1 vccd1 _08176_/D
+ sky130_fd_sc_hd__and4_1
X_05387_ _05387_/A _05444_/A vssd1 vssd1 vccd1 vccd1 _05440_/A sky130_fd_sc_hd__or2_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ _07165_/A _07126_/B _07137_/A vssd1 vssd1 vccd1 vccd1 _07127_/A sky130_fd_sc_hd__and3_1
XFILLER_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07057_ _07077_/A vssd1 vssd1 vccd1 vccd1 _07057_/Y sky130_fd_sc_hd__inv_2
X_06008_ _09877_/X _05998_/X _06272_/A _06002_/X _06005_/X vssd1 vssd1 vccd1 vccd1
+ _10206_/D sky130_fd_sc_hd__o221a_1
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07959_ _07954_/X _07958_/X _07954_/X _07958_/X vssd1 vssd1 vccd1 vccd1 _07959_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09629_ _09628_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09629_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10404_ _10437_/CLK _10404_/D vssd1 vssd1 vccd1 vccd1 _10404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ _10346_/CLK _10335_/D vssd1 vssd1 vccd1 vccd1 _10335_/Q sky130_fd_sc_hd__dfxtp_1
X_10266_ _10447_/CLK _10266_/D vssd1 vssd1 vccd1 vccd1 _10266_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10197_ _10202_/CLK _10197_/D vssd1 vssd1 vccd1 vccd1 _10197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05310_ _10346_/Q vssd1 vssd1 vccd1 vccd1 _05310_/Y sky130_fd_sc_hd__inv_2
X_06290_ _10130_/Q vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__inv_2
X_05241_ _10365_/Q _05239_/X input28/X _05240_/X _05236_/X vssd1 vssd1 vccd1 vccd1
+ _10365_/D sky130_fd_sc_hd__o221a_1
Xinput31 io_wb_dat_i[20] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 io_wb_dat_i[10] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
Xinput42 io_wb_dat_i[30] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05172_ _10397_/Q vssd1 vssd1 vccd1 vccd1 _05172_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09980_ _09979_/X _06626_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09980_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08931_ _08930_/A _08930_/B _08955_/A vssd1 vssd1 vccd1 vccd1 _08931_/X sky130_fd_sc_hd__a21bo_1
XFILLER_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _10287_/Q _07434_/X _08853_/X _08861_/X vssd1 vssd1 vccd1 vccd1 _08862_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_96_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07813_ _07837_/A _07868_/B _07813_/C _07837_/B vssd1 vssd1 vccd1 vccd1 _07813_/X
+ sky130_fd_sc_hd__or4_4
X_08793_ _08130_/X _08791_/B _08788_/X _08788_/X _08792_/X vssd1 vssd1 vccd1 vccd1
+ _08794_/C sky130_fd_sc_hd__a32o_1
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07744_ _10214_/Q _07687_/B _07594_/C _07885_/C _07743_/X vssd1 vssd1 vccd1 vccd1
+ _07744_/X sky130_fd_sc_hd__a41o_1
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07675_ _07659_/Y _07662_/X _07673_/X _07674_/X vssd1 vssd1 vccd1 vccd1 _07675_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06626_ _10376_/Q vssd1 vssd1 vccd1 vccd1 _06626_/Y sky130_fd_sc_hd__inv_2
X_09414_ _09359_/X _09413_/X _09359_/X _09413_/X vssd1 vssd1 vccd1 vccd1 _09414_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ _06560_/D _06556_/Y _06560_/D _06556_/Y vssd1 vssd1 vccd1 vccd1 _06557_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09345_ _09229_/X _09344_/X _09229_/X _09344_/X vssd1 vssd1 vccd1 vccd1 _09345_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09276_ _09276_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__or2_1
X_06488_ _08399_/A _06496_/A _10090_/Q _06462_/A vssd1 vssd1 vccd1 vccd1 _06495_/B
+ sky130_fd_sc_hd__a22o_1
X_05508_ _07164_/B vssd1 vssd1 vccd1 vccd1 _07218_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08227_ _08104_/X _08222_/Y _06255_/B vssd1 vssd1 vccd1 vccd1 _08227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05439_ _05439_/A vssd1 vssd1 vccd1 vccd1 _05439_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08158_ _06632_/Y _06030_/X _08153_/Y _08211_/A _08157_/X vssd1 vssd1 vccd1 vccd1
+ _08175_/B sky130_fd_sc_hd__o221a_1
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08089_ _10205_/Q vssd1 vssd1 vccd1 vccd1 _08303_/A sky130_fd_sc_hd__inv_2
X_07109_ _07112_/C _07109_/B vssd1 vssd1 vccd1 vccd1 _07109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10120_ _10244_/CLK _10120_/D vssd1 vssd1 vccd1 vccd1 _10120_/Q sky130_fd_sc_hd__dfxtp_1
X_10051_ _10447_/CLK _10051_/D vssd1 vssd1 vccd1 vccd1 _10051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10318_ _10343_/CLK _10318_/D vssd1 vssd1 vccd1 vccd1 _10318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10249_ _10249_/CLK _10249_/D vssd1 vssd1 vccd1 vccd1 _10249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05790_ _05790_/A vssd1 vssd1 vccd1 vccd1 _05791_/A sky130_fd_sc_hd__inv_2
XFILLER_207_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07460_ _05782_/X _07854_/B _10281_/Q _07456_/A vssd1 vssd1 vccd1 vccd1 _07460_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07391_ _07358_/A _07358_/B _07358_/X vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__a21bo_1
X_06411_ _06819_/B vssd1 vssd1 vccd1 vccd1 _06411_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09130_ _09354_/A _09258_/B _09354_/C _09259_/B vssd1 vssd1 vccd1 vccd1 _09130_/X
+ sky130_fd_sc_hd__o22a_1
X_06342_ _06313_/Y _06322_/A _06332_/A _06305_/Y _06341_/X vssd1 vssd1 vccd1 vccd1
+ _06343_/A sky130_fd_sc_hd__a41o_1
XFILLER_147_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09061_ _09060_/A _09060_/B _09060_/Y vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__a21oi_4
X_06273_ _06273_/A _06273_/B vssd1 vssd1 vccd1 vccd1 _09878_/S sky130_fd_sc_hd__nor2_4
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08012_ _08012_/A vssd1 vssd1 vccd1 vccd1 _08017_/A sky130_fd_sc_hd__inv_2
XFILLER_175_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05224_ _10375_/Q _05221_/X input39/X _05223_/X _05218_/X vssd1 vssd1 vccd1 vccd1
+ _10375_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05155_ _10433_/Q vssd1 vssd1 vccd1 vccd1 _05155_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _09962_/X _06625_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_2_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10334_/CLK sky130_fd_sc_hd__clkbuf_16
X_05086_ _05274_/A vssd1 vssd1 vccd1 vccd1 _05086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08914_ _08939_/C _08899_/X _08889_/A vssd1 vssd1 vccd1 vccd1 _08918_/A sky130_fd_sc_hd__a21oi_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09894_ _06857_/X _06415_/Y _10022_/S vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__mux2_2
XFILLER_111_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08845_ _08845_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _08845_/Y sky130_fd_sc_hd__nor2_1
X_08776_ _08759_/A _08759_/B _08760_/B vssd1 vssd1 vccd1 vccd1 _08797_/B sky130_fd_sc_hd__o21a_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05988_ _09781_/S _10043_/D vssd1 vssd1 vccd1 vccd1 _05990_/A sky130_fd_sc_hd__or2b_2
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07727_ _07719_/Y _07723_/X _07725_/X _07726_/X vssd1 vssd1 vccd1 vccd1 _07727_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07658_ _07910_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06609_ _10394_/Q _10393_/Q _10392_/Q _10391_/Q vssd1 vssd1 vccd1 vccd1 _06613_/A
+ sky130_fd_sc_hd__or4_4
X_07589_ _07597_/A _09921_/X vssd1 vssd1 vccd1 vccd1 _07589_/X sky130_fd_sc_hd__or2_1
X_09328_ _09326_/X _09327_/X _09326_/X _09327_/X vssd1 vssd1 vccd1 vccd1 _09328_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09259_ _09259_/A _09259_/B _09311_/A vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__or3_4
XFILLER_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10103_ _10207_/CLK _10103_/D vssd1 vssd1 vccd1 vccd1 _10103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10034_ _10205_/CLK input1/X vssd1 vssd1 vccd1 vccd1 _10035_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_191_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06960_ _07054_/C _06960_/B vssd1 vssd1 vccd1 vccd1 _06960_/X sky130_fd_sc_hd__or2_1
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05911_ _05911_/A vssd1 vssd1 vccd1 vccd1 _05911_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06891_ _06931_/A _09892_/X vssd1 vssd1 vccd1 vccd1 _06898_/C sky130_fd_sc_hd__nor2_2
X_08630_ _05018_/X _06657_/Y _08625_/Y _08629_/X vssd1 vssd1 vccd1 vccd1 _08630_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05842_ _05863_/A vssd1 vssd1 vccd1 vccd1 _05842_/X sky130_fd_sc_hd__clkbuf_2
X_08561_ _08624_/A _08456_/X _08457_/Y vssd1 vssd1 vccd1 vccd1 _08561_/X sky130_fd_sc_hd__a21o_1
X_05773_ input16/X _06081_/B _05773_/C input17/X vssd1 vssd1 vccd1 vccd1 _05923_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08492_ _10074_/Q _08492_/B vssd1 vssd1 vccd1 vccd1 _08494_/B sky130_fd_sc_hd__or2_1
X_07512_ _07496_/A _07496_/B _07496_/X vssd1 vssd1 vccd1 vccd1 _07513_/B sky130_fd_sc_hd__a21bo_1
XFILLER_35_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07443_ _08845_/B _07441_/B _07442_/Y vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__a21o_1
XFILLER_210_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _09112_/A _09112_/B _09162_/A vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__a21bo_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07374_ _07346_/X _07359_/X _07346_/X _07359_/X vssd1 vssd1 vccd1 vccd1 _07389_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_175_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06325_ _06322_/Y _06324_/A _06322_/A _06324_/Y vssd1 vssd1 vccd1 vccd1 _06325_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06256_ _10190_/Q _08230_/A vssd1 vssd1 vccd1 vccd1 _06257_/B sky130_fd_sc_hd__or2_2
X_09044_ _09259_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _09044_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05207_ _05202_/X _10382_/Q _05203_/X _09882_/X _05206_/X vssd1 vssd1 vccd1 vccd1
+ _10382_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06187_ _06203_/A vssd1 vssd1 vccd1 vccd1 _06187_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05138_ _05161_/A vssd1 vssd1 vccd1 vccd1 _05138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05069_ _10430_/Q _05064_/X input29/X _05065_/X _05062_/X vssd1 vssd1 vccd1 vccd1
+ _10430_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ _09019_/X _09017_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09946_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_22 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09876_/X input42/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _08504_/A _08726_/A _06263_/A _08728_/X _08827_/X vssd1 vssd1 vccd1 vccd1
+ _08828_/Y sky130_fd_sc_hd__a221oi_2
X_08759_ _08759_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10017_ _08049_/X _07397_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10017_/X sky130_fd_sc_hd__mux2_2
XFILLER_95_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06110_ _10331_/Q _06088_/X _10159_/Q _06089_/X _05105_/A vssd1 vssd1 vccd1 vccd1
+ _10159_/D sky130_fd_sc_hd__a221o_1
X_07090_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07253_/A sky130_fd_sc_hd__inv_2
X_06041_ _09829_/X _06028_/X _06260_/A _06031_/X _06032_/X vssd1 vssd1 vccd1 vccd1
+ _10194_/D sky130_fd_sc_hd__o221a_1
XFILLER_145_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09800_ _09799_/X _08226_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09800_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ _07750_/A _07750_/B _07750_/Y vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__o21ai_2
X_09731_ _06802_/Y _10396_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10062_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06943_ _06943_/A _06942_/X vssd1 vssd1 vccd1 vccd1 _06943_/X sky130_fd_sc_hd__or2b_1
X_09662_ _10144_/Q _10160_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09662_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06874_ _10223_/Q vssd1 vssd1 vccd1 vccd1 _07223_/A sky130_fd_sc_hd__inv_2
X_08613_ _10076_/Q vssd1 vssd1 vccd1 vccd1 _08613_/Y sky130_fd_sc_hd__inv_2
X_09593_ _08438_/Y _08436_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05825_ _05853_/A _05853_/B _05824_/Y vssd1 vssd1 vccd1 vccd1 _05826_/A sky130_fd_sc_hd__o21ai_2
X_08544_ _10052_/Q _08470_/B _08471_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__a21boi_2
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05756_ _05866_/A vssd1 vssd1 vccd1 vccd1 _05756_/X sky130_fd_sc_hd__buf_1
XFILLER_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08475_ _10057_/Q _08475_/B vssd1 vssd1 vccd1 vccd1 _08476_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_20_clock clkbuf_2_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10421_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05687_ _05771_/A _05684_/Y _05685_/Y _08061_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05688_/B sky130_fd_sc_hd__o32a_1
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ _07423_/Y _07921_/A _07417_/B vssd1 vssd1 vccd1 vccd1 _07426_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_23_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07357_ _06894_/C _07355_/X _06993_/B _07356_/X vssd1 vssd1 vccd1 vccd1 _07358_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06308_ _10132_/Q vssd1 vssd1 vccd1 vccd1 _08363_/A sky130_fd_sc_hd__inv_2
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _09027_/A _09026_/X vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__or2b_1
X_07288_ _07197_/X _07198_/X _07197_/X _07198_/X vssd1 vssd1 vccd1 vccd1 _07288_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06239_ _06235_/Y _06238_/X _06235_/Y _06238_/X vssd1 vssd1 vccd1 vccd1 _06239_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09929_ _08349_/X _06293_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 io_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05610_ _09994_/X _05540_/X _05626_/A vssd1 vssd1 vccd1 vccd1 _05621_/B sky130_fd_sc_hd__o21ai_1
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06590_ _10109_/Q _06466_/A _08450_/A _06489_/A vssd1 vssd1 vccd1 vccd1 _06590_/X
+ sky130_fd_sc_hd__a22o_1
X_05541_ _09994_/X _05540_/X _09994_/X _05540_/X vssd1 vssd1 vccd1 vccd1 _05627_/A
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08260_ _08260_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__or2_1
XFILLER_189_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05472_ _05472_/A _05472_/B vssd1 vssd1 vccd1 vccd1 _05472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _08191_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__or2_1
X_07211_ _07210_/A _07210_/B _07210_/Y vssd1 vssd1 vccd1 vccd1 _07211_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_158_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07142_ _07138_/A _07138_/B _07202_/B vssd1 vssd1 vccd1 vccd1 _07142_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07073_ _07073_/A vssd1 vssd1 vccd1 vccd1 _07074_/B sky130_fd_sc_hd__inv_2
X_06024_ _09849_/X _06015_/X _06265_/A _06017_/X _06018_/X vssd1 vssd1 vccd1 vccd1
+ _10199_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07975_ _07941_/X _07946_/X _07947_/X _07974_/X vssd1 vssd1 vccd1 vccd1 _07975_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09714_ _09713_/X _10381_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10047_/D sky130_fd_sc_hd__mux2_1
X_06926_ _06920_/A _06946_/A _06919_/Y _06917_/A _06925_/Y vssd1 vssd1 vccd1 vccd1
+ _06926_/X sky130_fd_sc_hd__o32a_2
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09645_ _10111_/Q input19/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__mux2_1
X_06857_ _06856_/A _06856_/B _07023_/B vssd1 vssd1 vccd1 vccd1 _06857_/X sky130_fd_sc_hd__a21bo_1
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05808_ _10271_/Q vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__inv_2
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06788_ _09717_/S _06788_/B vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__and2_1
X_09576_ _08407_/Y _10124_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08527_ _08269_/A _08509_/A _08265_/A _08526_/B vssd1 vssd1 vccd1 vccd1 _08597_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05739_ _10267_/Q vssd1 vssd1 vccd1 vccd1 _07594_/C sky130_fd_sc_hd__buf_2
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _10047_/Q vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__inv_2
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07410_/B sky130_fd_sc_hd__or2_1
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10420_ _10420_/CLK _10420_/D vssd1 vssd1 vccd1 vccd1 _10420_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08389_ _08413_/B vssd1 vssd1 vccd1 vccd1 _08409_/B sky130_fd_sc_hd__buf_1
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _10447_/CLK _10351_/D vssd1 vssd1 vccd1 vccd1 _10351_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10282_ _10297_/CLK _10282_/D vssd1 vssd1 vccd1 vccd1 _10282_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07760_ _07760_/A _07760_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__or2_1
XFILLER_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06711_ _10368_/Q _08727_/A _08724_/A vssd1 vssd1 vccd1 vccd1 _06807_/B sky130_fd_sc_hd__a21boi_4
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09430_ _09430_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _09430_/X sky130_fd_sc_hd__or2_1
X_07691_ _07673_/X _07674_/X _07673_/X _07674_/X vssd1 vssd1 vccd1 vccd1 _07692_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06642_ _08753_/A vssd1 vssd1 vccd1 vccd1 _06642_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06573_ _06570_/X _06572_/Y _06570_/X _06572_/Y vssd1 vssd1 vccd1 vccd1 _06573_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09361_ _09311_/Y _09285_/A _09311_/A _09285_/Y vssd1 vssd1 vccd1 vccd1 _09361_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08312_ _08312_/A vssd1 vssd1 vccd1 vccd1 _08616_/A sky130_fd_sc_hd__clkbuf_2
X_09292_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09343_/C sky130_fd_sc_hd__or2_2
X_05524_ _09992_/X _10021_/X _05483_/X _05523_/X vssd1 vssd1 vccd1 vccd1 _05524_/X
+ sky130_fd_sc_hd__o22a_1
X_08243_ _08533_/A _08241_/B _08240_/X _08242_/Y vssd1 vssd1 vccd1 vccd1 _08243_/Y
+ sky130_fd_sc_hd__a211oi_2
X_05455_ _05455_/A vssd1 vssd1 vccd1 vccd1 _10318_/D sky130_fd_sc_hd__inv_2
XFILLER_177_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08174_ _10361_/Q _08166_/X _10371_/Q _08169_/X _08173_/X vssd1 vssd1 vccd1 vccd1
+ _08175_/D sky130_fd_sc_hd__o221a_1
X_05386_ _05386_/A _05448_/A vssd1 vssd1 vccd1 vccd1 _05444_/A sky130_fd_sc_hd__or2_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ _07125_/A _07189_/A vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__or2_1
XFILLER_161_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07056_ _07056_/A _07126_/B _07056_/C vssd1 vssd1 vccd1 vccd1 _07077_/A sky130_fd_sc_hd__and3_1
X_06007_ _10206_/Q vssd1 vssd1 vccd1 vccd1 _06272_/A sky130_fd_sc_hd__buf_1
XFILLER_161_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07958_ _07785_/X _07955_/X _07956_/X _07957_/X vssd1 vssd1 vccd1 vccd1 _07958_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07889_ _07875_/X _07888_/X _07875_/X _07888_/X vssd1 vssd1 vccd1 vccd1 _07889_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06909_ _06909_/A _06909_/B vssd1 vssd1 vccd1 vccd1 _06920_/A sky130_fd_sc_hd__or2_1
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09628_ _09627_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09559_ _09558_/X _10354_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09559_/X sky130_fd_sc_hd__mux2_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10403_ _10436_/CLK _10403_/D vssd1 vssd1 vccd1 vccd1 _10403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10334_ _10334_/CLK _10334_/D vssd1 vssd1 vccd1 vccd1 _10334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10265_ _10298_/CLK _10265_/D vssd1 vssd1 vccd1 vccd1 _10265_/Q sky130_fd_sc_hd__dfxtp_1
X_10196_ _10202_/CLK _10196_/D vssd1 vssd1 vccd1 vccd1 _10196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05240_ _05240_/A vssd1 vssd1 vccd1 vccd1 _05240_/X sky130_fd_sc_hd__clkbuf_2
Xinput21 io_wb_dat_i[11] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_4
Xinput10 io_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
Xinput43 io_wb_dat_i[31] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_4
X_05171_ _05179_/A _05171_/B vssd1 vssd1 vccd1 vccd1 _10398_/D sky130_fd_sc_hd__nor2_1
Xinput32 io_wb_dat_i[21] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_143_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08930_ _08930_/A _08930_/B vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__or2_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ _10286_/Q _07415_/Y _08855_/Y _08860_/X vssd1 vssd1 vccd1 vccd1 _08861_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07812_ _07812_/A _07811_/X vssd1 vssd1 vccd1 vccd1 _07812_/X sky130_fd_sc_hd__or2b_1
X_08792_ _08791_/A _08791_/B _08181_/B _08790_/Y _08791_/Y vssd1 vssd1 vccd1 vccd1
+ _08792_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07743_ _07485_/A _07765_/A _07686_/A _07868_/A vssd1 vssd1 vccd1 vccd1 _07743_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07674_ _07659_/Y _07662_/X _07659_/Y _07662_/X vssd1 vssd1 vccd1 vccd1 _07674_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06625_ _10377_/Q vssd1 vssd1 vccd1 vccd1 _06625_/Y sky130_fd_sc_hd__inv_2
X_09413_ _09411_/X _09412_/X _09411_/X _09412_/X vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06556_ _08432_/A _06489_/X _06560_/C _06552_/X vssd1 vssd1 vccd1 vccd1 _06556_/Y
+ sky130_fd_sc_hd__o22ai_1
X_09344_ _09344_/A _09343_/X vssd1 vssd1 vccd1 vccd1 _09344_/X sky130_fd_sc_hd__or2b_1
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__inv_2
X_06487_ _06487_/A vssd1 vssd1 vccd1 vccd1 _06496_/A sky130_fd_sc_hd__clkbuf_2
X_05507_ _07152_/D vssd1 vssd1 vccd1 vccd1 _07164_/B sky130_fd_sc_hd__inv_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08226_ _08160_/X _08224_/B _08184_/A _08225_/Y vssd1 vssd1 vccd1 vccd1 _08226_/Y
+ sky130_fd_sc_hd__a211oi_4
X_05438_ _05438_/A vssd1 vssd1 vccd1 vccd1 _10322_/D sky130_fd_sc_hd__inv_2
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08157_ _10352_/Q _08155_/X _10374_/Q _08293_/A vssd1 vssd1 vccd1 vccd1 _08157_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05369_ _05369_/A _10209_/Q vssd1 vssd1 vccd1 vccd1 _05399_/A sky130_fd_sc_hd__or2_1
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07108_ _07108_/A _07108_/B _07197_/A vssd1 vssd1 vccd1 vccd1 _07109_/B sky130_fd_sc_hd__and3_1
X_08088_ _08084_/Y _06253_/A _06635_/Y _10193_/Q _08087_/X vssd1 vssd1 vccd1 vccd1
+ _08098_/B sky130_fd_sc_hd__o221a_1
XFILLER_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07039_ _06927_/X _06938_/X _06881_/X _06939_/X vssd1 vssd1 vccd1 vccd1 _07039_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _10447_/CLK _10050_/D vssd1 vssd1 vccd1 vccd1 _10050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ _10330_/CLK _10317_/D vssd1 vssd1 vccd1 vccd1 _10317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10248_ _10249_/CLK _10248_/D vssd1 vssd1 vccd1 vccd1 _10248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _10447_/CLK _10179_/D vssd1 vssd1 vccd1 vccd1 _10179_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06410_ _06407_/X _06409_/Y _06407_/X _06409_/Y vssd1 vssd1 vccd1 vccd1 _06410_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07390_ _07390_/A vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__inv_2
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06341_ _10241_/Q _08378_/A _06330_/Y _06335_/X vssd1 vssd1 vccd1 vccd1 _06341_/X
+ sky130_fd_sc_hd__o22a_1
X_06272_ _06272_/A _08301_/A vssd1 vssd1 vccd1 vccd1 _06273_/B sky130_fd_sc_hd__or2_2
XFILLER_147_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09060_ _09060_/A _09060_/B vssd1 vssd1 vccd1 vccd1 _09060_/Y sky130_fd_sc_hd__nor2_4
XFILLER_175_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05223_ _05264_/A vssd1 vssd1 vccd1 vccd1 _05223_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08011_ _08011_/A vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__inv_2
XFILLER_162_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05154_ _10401_/Q vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__inv_2
X_09962_ _06614_/B _08309_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09962_/X sky130_fd_sc_hd__mux2_1
X_05085_ _06099_/A vssd1 vssd1 vccd1 vccd1 _05274_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08913_ _08913_/A _08912_/X vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__or2b_1
XFILLER_134_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09893_ _06849_/X _05858_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09893_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08844_ _10294_/Q vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__inv_2
X_08775_ _10352_/Q _08752_/B _08759_/B vssd1 vssd1 vccd1 vccd1 _08775_/Y sky130_fd_sc_hd__a21oi_1
X_05987_ _06183_/A _06082_/B _06184_/A _08329_/D vssd1 vssd1 vccd1 vccd1 _09781_/S
+ sky130_fd_sc_hd__nor4_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07726_ _07719_/Y _07723_/X _07719_/Y _07723_/X vssd1 vssd1 vccd1 vccd1 _07726_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07657_ _07678_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06608_ _06606_/X _06607_/Y _05018_/X _06739_/A vssd1 vssd1 vccd1 vccd1 _06608_/X
+ sky130_fd_sc_hd__a22o_1
X_07588_ _07588_/A _09920_/X vssd1 vssd1 vccd1 vccd1 _07588_/X sky130_fd_sc_hd__or2_1
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06539_ _06539_/A _06539_/B _06539_/C vssd1 vssd1 vccd1 vccd1 _06542_/A sky130_fd_sc_hd__or3_1
X_09327_ _09227_/X _09241_/X _09242_/X _09270_/X vssd1 vssd1 vccd1 vccd1 _09327_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _09258_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__or2_2
XFILLER_181_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08209_ _08121_/X _08208_/B _08211_/B _08240_/A vssd1 vssd1 vccd1 vccd1 _08209_/Y
+ sky130_fd_sc_hd__a211oi_4
X_09189_ _09045_/X _09144_/X _09145_/X _09146_/X vssd1 vssd1 vccd1 vccd1 _09189_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10102_ _10102_/CLK _10102_/D vssd1 vssd1 vccd1 vccd1 _10102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10033_ _10042_/Q _09565_/X _08387_/Y _09566_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10033_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05910_ _05910_/A vssd1 vssd1 vccd1 vccd1 _05910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06890_ _06888_/X _06889_/X _06888_/X _06889_/X vssd1 vssd1 vccd1 vccd1 _06897_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05841_ _10263_/Q _05780_/X _05637_/X _06856_/A _05764_/X vssd1 vssd1 vccd1 vccd1
+ _10263_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08560_ _08130_/X _08558_/B _08559_/X vssd1 vssd1 vccd1 vccd1 _08560_/X sky130_fd_sc_hd__a21o_1
X_05772_ _07594_/C _05467_/X _06176_/A _05771_/X vssd1 vssd1 vccd1 vccd1 _10267_/D
+ sky130_fd_sc_hd__o211a_1
X_08491_ _10073_/Q _08491_/B vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__or2_1
X_07511_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07513_/A sky130_fd_sc_hd__or2_1
XFILLER_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07442_ _07454_/B vssd1 vssd1 vccd1 vccd1 _07442_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ _07340_/X _07360_/X _07340_/X _07360_/X vssd1 vssd1 vccd1 vccd1 _07388_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_210_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09112_/A _09112_/B vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__or2_1
X_06324_ _06324_/A vssd1 vssd1 vccd1 vccd1 _06324_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06255_ _10189_/Q _06255_/B vssd1 vssd1 vccd1 vccd1 _08230_/A sky130_fd_sc_hd__or2_1
X_09043_ _09043_/A vssd1 vssd1 vccd1 vccd1 _09043_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05206_ _05236_/A vssd1 vssd1 vccd1 vccd1 _05206_/X sky130_fd_sc_hd__clkbuf_4
X_06186_ _06224_/A vssd1 vssd1 vccd1 vccd1 _06203_/A sky130_fd_sc_hd__clkbuf_2
X_05137_ _10437_/Q vssd1 vssd1 vccd1 vccd1 _05137_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05068_ _10431_/Q _05064_/X input31/X _05065_/X _05062_/X vssd1 vssd1 vccd1 vccd1
+ _10431_/D sky130_fd_sc_hd__o221a_1
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _09223_/Y _09222_/B _09994_/S vssd1 vssd1 vccd1 vccd1 _09945_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09876_ _09875_/X _08310_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__mux2_1
X_08827_ _06262_/A _08730_/Y _06263_/A _08728_/X _08826_/X vssd1 vssd1 vccd1 vccd1
+ _08827_/X sky130_fd_sc_hd__o221a_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_23 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_12 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08758_ _10352_/Q _08758_/B vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__nor2_2
XFILLER_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08689_ _08169_/X _10069_/Q _08616_/A _10076_/Q _08688_/X vssd1 vssd1 vccd1 vccd1
+ _08695_/C sky130_fd_sc_hd__a221o_1
X_07709_ _07705_/X _07708_/X _07705_/X _07708_/X vssd1 vssd1 vccd1 vccd1 _07709_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10016_ _08005_/A _08036_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10016_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10343_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06040_ _10194_/Q vssd1 vssd1 vccd1 vccd1 _06260_/A sky130_fd_sc_hd__buf_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07991_ _07770_/X _07969_/X _07770_/X _07969_/X vssd1 vssd1 vccd1 vccd1 _08008_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09730_ _06801_/Y _10395_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10061_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06942_ _06942_/A _09894_/X _06942_/C _09895_/X vssd1 vssd1 vccd1 vccd1 _06942_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09661_ _10143_/Q _10159_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06873_ _07056_/A _06868_/Y _05956_/X _06870_/Y _06872_/X vssd1 vssd1 vccd1 vccd1
+ _06880_/A sky130_fd_sc_hd__a41o_1
X_08612_ _08309_/A _08495_/Y _08611_/X vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__a21o_1
X_09592_ _08435_/X _08434_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09592_/X sky130_fd_sc_hd__mux2_1
X_05824_ _05788_/A _10260_/Q _05823_/Y vssd1 vssd1 vccd1 vccd1 _05824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08543_ _10186_/Q _08573_/B _10185_/Q _08542_/Y vssd1 vssd1 vccd1 vccd1 _08592_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05755_ _10275_/Q _05751_/X _09637_/X _05753_/X _05747_/X vssd1 vssd1 vccd1 vccd1
+ _10275_/D sky130_fd_sc_hd__o221a_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ _10056_/Q _08474_/B vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__or2_1
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05686_ _10301_/Q vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__inv_2
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _07425_/A vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__buf_2
XFILLER_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07356_ _06894_/C _07355_/X _06894_/C _07355_/X vssd1 vssd1 vccd1 vccd1 _07356_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06307_ _06304_/A _06302_/X _06304_/A _06302_/X vssd1 vssd1 vccd1 vccd1 _06307_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_07287_ _07285_/X _07286_/Y _07285_/X _07286_/Y vssd1 vssd1 vccd1 vccd1 _07287_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06238_ _10039_/D _06236_/Y _06237_/Y _10039_/Q vssd1 vssd1 vccd1 vccd1 _06238_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ _09038_/A _09128_/A _09074_/C vssd1 vssd1 vccd1 vccd1 _09026_/X sky130_fd_sc_hd__or3_4
XFILLER_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06169_ _06169_/A _09673_/X vssd1 vssd1 vccd1 vccd1 _10122_/D sky130_fd_sc_hd__and2_1
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09928_ _09927_/X _07828_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09928_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09859_ _10373_/Q _09858_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09859_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 io_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05540_ _05538_/Y _05539_/Y _05538_/Y _05539_/Y vssd1 vssd1 vccd1 vccd1 _05540_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05471_ _10015_/X vssd1 vssd1 vccd1 vccd1 _05472_/B sky130_fd_sc_hd__inv_2
X_08190_ _10179_/Q _06245_/B _06246_/B vssd1 vssd1 vccd1 vccd1 _08190_/X sky130_fd_sc_hd__a21o_1
X_07210_ _07210_/A _07210_/B vssd1 vssd1 vccd1 vccd1 _07210_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07141_ _07119_/X _07140_/X _07119_/X _07140_/X vssd1 vssd1 vccd1 vccd1 _07141_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ _07234_/A _07072_/B vssd1 vssd1 vccd1 vccd1 _07073_/A sky130_fd_sc_hd__or2_2
X_06023_ _10199_/Q vssd1 vssd1 vccd1 vccd1 _06265_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07974_ _07948_/X _07952_/X _07953_/X _07973_/X vssd1 vssd1 vccd1 vccd1 _07974_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _10448_/Q _06742_/A _09717_/S vssd1 vssd1 vccd1 vccd1 _09713_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06925_ _06925_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _06925_/Y sky130_fd_sc_hd__nor2_1
X_09644_ _06408_/X _06410_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09644_/X sky130_fd_sc_hd__mux2_1
X_06856_ _06856_/A _06856_/B vssd1 vssd1 vccd1 vccd1 _07023_/B sky130_fd_sc_hd__or2_1
X_05807_ _05804_/A _10255_/Q _05805_/A _05806_/Y vssd1 vssd1 vccd1 vccd1 _05807_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06787_ _06614_/A _06692_/Y _06620_/A _06786_/X vssd1 vssd1 vccd1 vccd1 _09745_/S
+ sky130_fd_sc_hd__o211a_4
X_09575_ _08404_/Y _09574_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09575_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08526_ _08526_/A _08526_/B vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__nor2_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05738_ _10284_/Q _05728_/X _07423_/A _05732_/X _05737_/X vssd1 vssd1 vccd1 vccd1
+ _10284_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08457_/A _10048_/Q vssd1 vssd1 vccd1 vccd1 _08457_/Y sky130_fd_sc_hd__nor2_1
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05669_ _10304_/Q vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__inv_2
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07408_ _07408_/A _07408_/B vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__or2_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08388_ _08388_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08388_/Y sky130_fd_sc_hd__nor2_1
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07339_ _07035_/X _07335_/X _07336_/X _07338_/X vssd1 vssd1 vccd1 vccd1 _07339_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _10447_/CLK _10350_/D vssd1 vssd1 vccd1 vccd1 _10350_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_191_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09009_ _09070_/A _09089_/B vssd1 vssd1 vccd1 vccd1 _09009_/X sky130_fd_sc_hd__or2_2
XFILLER_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _10298_/CLK _10281_/D vssd1 vssd1 vccd1 vccd1 _10281_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06710_ _06710_/A vssd1 vssd1 vccd1 vccd1 _06810_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_34_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10329_/CLK sky130_fd_sc_hd__clkbuf_16
X_07690_ _07685_/X _07689_/X _07685_/X _07689_/X vssd1 vssd1 vccd1 vccd1 _07722_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06641_ _10391_/Q vssd1 vssd1 vccd1 vccd1 _06641_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06572_ _06563_/X _06566_/X _06571_/X vssd1 vssd1 vccd1 vccd1 _06572_/Y sky130_fd_sc_hd__o21ai_2
X_09360_ _09359_/A _09359_/B _09359_/X vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__a21bo_1
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ _06273_/A _06273_/B _09878_/S vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09291_ _09457_/C _09451_/B vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__or2_2
X_05523_ _10003_/X _09995_/X _05486_/Y _05558_/A vssd1 vssd1 vccd1 vccd1 _05523_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08242_ _08245_/B vssd1 vssd1 vccd1 vccd1 _08242_/Y sky130_fd_sc_hd__inv_2
X_05454_ _05449_/B _05439_/X _05452_/Y _05453_/Y _05424_/A vssd1 vssd1 vccd1 vccd1
+ _05455_/A sky130_fd_sc_hd__o32a_1
XFILLER_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08173_ _06664_/A _06072_/X _10363_/Q _08172_/X vssd1 vssd1 vccd1 vccd1 _08173_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05385_ _10318_/Q _05452_/B vssd1 vssd1 vccd1 vccd1 _05448_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07124_ _07111_/X _07112_/X _07111_/X _07112_/X vssd1 vssd1 vccd1 vccd1 _07124_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_173_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07055_ _07055_/A _07054_/X vssd1 vssd1 vccd1 vccd1 _07055_/X sky130_fd_sc_hd__or2b_1
X_06006_ _09881_/X _05998_/X _06273_/A _06002_/X _06005_/X vssd1 vssd1 vccd1 vccd1
+ _10207_/D sky130_fd_sc_hd__o221a_1
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07957_ _07785_/X _07955_/X _07785_/A _07955_/X vssd1 vssd1 vccd1 vccd1 _07957_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06908_ _06897_/A _06897_/B _06897_/X vssd1 vssd1 vccd1 vccd1 _06909_/B sky130_fd_sc_hd__a21bo_1
X_07888_ _07879_/X _07883_/X _07886_/X _07887_/X vssd1 vssd1 vccd1 vccd1 _07888_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09627_ _09626_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09627_/X sky130_fd_sc_hd__mux2_1
X_06839_ _10220_/Q vssd1 vssd1 vccd1 vccd1 _07164_/A sky130_fd_sc_hd__inv_2
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09558_ _10386_/Q _10183_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09558_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08509_ _08509_/A vssd1 vssd1 vccd1 vccd1 _08509_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ vssd1 vssd1 vccd1 vccd1 _09489_/HI _09613_/A1 sky130_fd_sc_hd__conb_1
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ _10436_/CLK _10402_/D vssd1 vssd1 vccd1 vccd1 _10402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ _10334_/CLK _10333_/D vssd1 vssd1 vccd1 vccd1 _10333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10264_ _10298_/CLK _10264_/D vssd1 vssd1 vccd1 vccd1 _10264_/Q sky130_fd_sc_hd__dfxtp_1
X_10195_ _10399_/CLK _10195_/D vssd1 vssd1 vccd1 vccd1 _10195_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 io_wb_dat_i[12] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_4
Xinput11 io_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
XFILLER_190_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05170_ _05153_/X _05168_/Y _05169_/Y _05161_/X vssd1 vssd1 vccd1 vccd1 _05171_/B
+ sky130_fd_sc_hd__o22a_1
Xinput33 io_wb_dat_i[22] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput44 io_wb_dat_i[3] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_4
XFILLER_155_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08860_ _10285_/Q _07421_/Y _08895_/A _08859_/X vssd1 vssd1 vccd1 vccd1 _08860_/X
+ sky130_fd_sc_hd__o22a_1
X_07811_ _07811_/A _07897_/B _07811_/C _09914_/X vssd1 vssd1 vccd1 vccd1 _07811_/X
+ sky130_fd_sc_hd__or4_4
X_08791_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07742_ _07642_/X _07644_/X _07642_/X _07644_/X vssd1 vssd1 vccd1 vccd1 _07742_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07673_ _07663_/X _07664_/X _07671_/X _07672_/X vssd1 vssd1 vccd1 vccd1 _07673_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06624_ _10378_/Q vssd1 vssd1 vccd1 vccd1 _06624_/Y sky130_fd_sc_hd__inv_2
X_09412_ _09341_/X _09351_/X _09352_/X _09356_/X vssd1 vssd1 vccd1 vccd1 _09412_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09343_ _09343_/A _09470_/B _09343_/C vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__or3_1
X_06555_ _10102_/Q _06463_/A _08434_/A _06540_/A vssd1 vssd1 vccd1 vccd1 _06560_/D
+ sky130_fd_sc_hd__a22o_1
X_09274_ _09224_/X _09273_/X _09224_/X _09273_/X vssd1 vssd1 vccd1 vccd1 _09275_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06486_ _10090_/Q vssd1 vssd1 vccd1 vccd1 _08399_/A sky130_fd_sc_hd__inv_2
X_05506_ _05510_/A _05505_/B _05505_/Y vssd1 vssd1 vccd1 vccd1 _07152_/D sky130_fd_sc_hd__a21oi_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08225_ _08228_/B vssd1 vssd1 vccd1 vccd1 _08225_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05437_ _05432_/B _05416_/X _05436_/Y _05389_/A _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05438_/A sky130_fd_sc_hd__o32a_1
X_08156_ _10203_/Q vssd1 vssd1 vccd1 vccd1 _08293_/A sky130_fd_sc_hd__inv_2
X_05368_ _06086_/A _10331_/Q _05296_/B _05312_/B vssd1 vssd1 vccd1 vccd1 _10331_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07107_ _07150_/A _09890_/X vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__or2_2
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08087_ _06638_/Y _08751_/A _08761_/A _08086_/X vssd1 vssd1 vccd1 vccd1 _08087_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05299_ _05299_/A _05355_/A vssd1 vssd1 vccd1 vccd1 _05351_/A sky130_fd_sc_hd__or2_1
XFILLER_161_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07038_ _06949_/X _07037_/X _06949_/X _07037_/X vssd1 vssd1 vccd1 vccd1 _07038_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__nor2_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10316_ _10330_/CLK _10316_/D vssd1 vssd1 vccd1 vccd1 _10316_/Q sky130_fd_sc_hd__dfxtp_1
X_10247_ _10249_/CLK _10247_/D vssd1 vssd1 vccd1 vccd1 _10247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10178_ _10178_/CLK _10178_/D vssd1 vssd1 vccd1 vccd1 _10178_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06340_ _10134_/Q vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__inv_2
X_06271_ _06271_/A _06271_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__or2_1
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05222_ _05240_/A vssd1 vssd1 vccd1 vccd1 _05264_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08010_ _08010_/A vssd1 vssd1 vccd1 vccd1 _08019_/A sky130_fd_sc_hd__inv_2
XFILLER_162_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05153_ _05202_/A vssd1 vssd1 vccd1 vccd1 _05153_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _09960_/X _10370_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09961_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05084_ input20/X _05082_/X _10421_/Q _05083_/X _08623_/A vssd1 vssd1 vccd1 vccd1
+ _10421_/D sky130_fd_sc_hd__a221o_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08912_ _08912_/A _09010_/B _08936_/C vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__or3_4
XFILLER_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09892_ _06848_/X _06413_/Y _10022_/S vssd1 vssd1 vccd1 vccd1 _09892_/X sky130_fd_sc_hd__mux2_2
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08843_ _10295_/Q _07458_/Y _10295_/Q _07458_/Y vssd1 vssd1 vccd1 vccd1 _08843_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08774_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08774_/X sky130_fd_sc_hd__or2_1
XFILLER_111_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05986_ _05038_/X _05970_/X _07854_/D _05971_/X _05985_/X vssd1 vssd1 vccd1 vccd1
+ _10210_/D sky130_fd_sc_hd__a221o_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07725_ _07885_/A _07516_/B _07885_/C _07634_/Y _07724_/X vssd1 vssd1 vccd1 vccd1
+ _07725_/X sky130_fd_sc_hd__a41o_1
XFILLER_65_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07656_ _07768_/A vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__inv_2
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06607_ _10383_/Q vssd1 vssd1 vccd1 vccd1 _06607_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07587_ _07613_/B _07765_/A _07667_/A _07587_/D vssd1 vssd1 vccd1 vccd1 _07587_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06538_ _06538_/A vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__inv_2
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _09308_/X _09325_/X _09308_/X _09325_/X vssd1 vssd1 vccd1 vccd1 _09326_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09257_ _09245_/A _09259_/B _09310_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _09261_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__nor2_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06469_ _10087_/Q vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__inv_2
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09188_ _09186_/X _09187_/X _09186_/X _09187_/X vssd1 vssd1 vccd1 vccd1 _09188_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_181_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08139_ _10353_/Q vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__inv_2
XFILLER_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _10102_/CLK _10101_/D vssd1 vssd1 vccd1 vccd1 _10101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10032_ _10444_/Q _09562_/X _08384_/Y _09563_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10032_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05840_ _05828_/X _05839_/X _05828_/X _05839_/X vssd1 vssd1 vccd1 vccd1 _06856_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05771_ _05771_/A _05771_/B _05771_/C vssd1 vssd1 vccd1 vccd1 _05771_/X sky130_fd_sc_hd__or3_1
X_07510_ _07483_/A _07516_/B _07913_/A vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__a21oi_1
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08490_ _10072_/Q _08490_/B vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__or2_1
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07441_ _10278_/Q _07441_/B vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__or2_1
XFILLER_210_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07372_ _07361_/X _07371_/X _07361_/X _07371_/X vssd1 vssd1 vccd1 vccd1 _07387_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09111_ _09111_/A vssd1 vssd1 vccd1 vccd1 _09112_/B sky130_fd_sc_hd__inv_2
X_06323_ _06311_/A _10132_/Q _06312_/A _06315_/Y vssd1 vssd1 vccd1 vccd1 _06324_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06254_ _06254_/A _08222_/A vssd1 vssd1 vccd1 vccd1 _06255_/B sky130_fd_sc_hd__or2_1
X_09042_ _09258_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__or2_2
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06185_ _06185_/A _09944_/S vssd1 vssd1 vccd1 vccd1 _06224_/A sky130_fd_sc_hd__or2_2
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05205_ _05202_/X _10383_/Q _05203_/X _09898_/X _05198_/X vssd1 vssd1 vccd1 vccd1
+ _10383_/D sky130_fd_sc_hd__o221a_1
X_05136_ _10405_/Q vssd1 vssd1 vccd1 vccd1 _06615_/B sky130_fd_sc_hd__inv_2
XFILLER_143_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05067_ _10432_/Q _05064_/X input32/X _05065_/X _05062_/X vssd1 vssd1 vccd1 vccd1
+ _10432_/D sky130_fd_sc_hd__o221a_1
X_09944_ _09943_/X _10041_/Q _09944_/S vssd1 vssd1 vccd1 vccd1 _09944_/X sky130_fd_sc_hd__mux2_1
X_09875_ _10377_/Q _09874_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09875_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08826_ _08737_/X _08812_/X _08825_/X vssd1 vssd1 vccd1 vccd1 _08826_/X sky130_fd_sc_hd__a21o_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_13 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08757_ _08804_/A _08804_/B _08539_/A _08756_/Y vssd1 vssd1 vccd1 vccd1 _08822_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05969_ _05971_/A vssd1 vssd1 vccd1 vccd1 _05970_/A sky130_fd_sc_hd__inv_2
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08688_ _08307_/A _10075_/Q _08304_/A _10074_/Q vssd1 vssd1 vccd1 vccd1 _08688_/X
+ sky130_fd_sc_hd__a22o_1
X_07708_ _07707_/A _07707_/B _07707_/X vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__a21bo_1
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07639_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07640_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _09246_/X _09249_/X _09250_/X _09264_/X vssd1 vssd1 vccd1 vccd1 _09309_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10015_ _08031_/X _07387_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10015_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07990_ _07971_/A _07971_/B _07971_/X vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__a21bo_1
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06941_ _06942_/A _09894_/X _06961_/A _07021_/B vssd1 vssd1 vccd1 vccd1 _06943_/A
+ sky130_fd_sc_hd__o22a_1
X_09660_ _10126_/Q input25/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08611_ _08309_/A _08495_/Y _08610_/Y vssd1 vssd1 vccd1 vccd1 _08611_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06872_ _07054_/C _06949_/D _07031_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _06872_/X
+ sky130_fd_sc_hd__o22a_1
X_09591_ _08433_/Y _08432_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05823_ _08847_/B _05792_/Y _05793_/X _05822_/X vssd1 vssd1 vccd1 vccd1 _05823_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08542_ _08542_/A vssd1 vssd1 vccd1 vccd1 _08542_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05754_ _05790_/A _05751_/X _09638_/X _05753_/X _05747_/X vssd1 vssd1 vccd1 vccd1
+ _10276_/D sky130_fd_sc_hd__o221a_1
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08473_ _10055_/Q _08473_/B vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__or2_1
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05685_ _05685_/A _05685_/B vssd1 vssd1 vccd1 vccd1 _05685_/Y sky130_fd_sc_hd__nor2_1
X_07424_ _07686_/A vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__buf_2
XFILLER_24_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ _07283_/X _07296_/Y _07297_/X _07299_/A vssd1 vssd1 vccd1 vccd1 _07355_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06306_ _06304_/A _06304_/B _06305_/Y vssd1 vssd1 vccd1 vccd1 _06306_/Y sky130_fd_sc_hd__a21oi_1
X_07286_ _07245_/A _07245_/B _07246_/B vssd1 vssd1 vccd1 vccd1 _07286_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_191_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06237_ _10039_/D vssd1 vssd1 vccd1 vccd1 _06237_/Y sky130_fd_sc_hd__inv_2
X_09025_ _08998_/A _09938_/X _08912_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _09027_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06168_ _06169_/A _09674_/X vssd1 vssd1 vccd1 vccd1 _10123_/D sky130_fd_sc_hd__and2_1
X_05119_ _05116_/X _06614_/B _05118_/Y _05113_/X vssd1 vssd1 vccd1 vccd1 _05120_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06099_ _06099_/A vssd1 vssd1 vccd1 vccd1 _06099_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09927_ _09926_/X _06962_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09858_ _08288_/Y _10373_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09858_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08809_ _08809_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__nor2_1
X_09789_ _09788_/X input49/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05470_ _10011_/X vssd1 vssd1 vccd1 vccd1 _05472_/A sky130_fd_sc_hd__inv_2
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07140_ _07134_/A _07129_/X _07133_/Y _07131_/A _07139_/Y vssd1 vssd1 vccd1 vccd1
+ _07140_/X sky130_fd_sc_hd__o32a_1
XFILLER_173_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07071_ _07055_/X _07057_/Y _07069_/X _07070_/X vssd1 vssd1 vccd1 vccd1 _07071_/X
+ sky130_fd_sc_hd__o22a_1
X_06022_ _09853_/X _06015_/X _10200_/Q _06017_/X _06018_/X vssd1 vssd1 vccd1 vccd1
+ _10200_/D sky130_fd_sc_hd__o221a_1
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _09711_/X _10380_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10046_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07973_ _07954_/X _07958_/X _07959_/X _07972_/X vssd1 vssd1 vccd1 vccd1 _07973_/X
+ sky130_fd_sc_hd__o22a_1
X_06924_ _06924_/A _06924_/B vssd1 vssd1 vccd1 vccd1 _06945_/B sky130_fd_sc_hd__nor2_2
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09643_ _06402_/Y _06403_/Y _10175_/Q vssd1 vssd1 vccd1 vccd1 _09643_/X sky130_fd_sc_hd__mux2_1
X_06855_ _06855_/A _06855_/B vssd1 vssd1 vccd1 vccd1 _06856_/B sky130_fd_sc_hd__or2_1
X_09574_ _08402_/Y _09573_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__mux2_1
X_05806_ _10255_/Q vssd1 vssd1 vccd1 vccd1 _05806_/Y sky130_fd_sc_hd__inv_2
X_08525_ _08524_/Y _08511_/Y _08484_/B vssd1 vssd1 vccd1 vccd1 _08526_/B sky130_fd_sc_hd__o21ai_1
X_06786_ _06614_/B _06694_/Y _06614_/A _06692_/Y _06785_/X vssd1 vssd1 vccd1 vccd1
+ _06786_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05737_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05737_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _10048_/Q vssd1 vssd1 vccd1 vccd1 _08456_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05668_ _05668_/A _05668_/B vssd1 vssd1 vccd1 vccd1 _05668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _09525_/X _08391_/B vssd1 vssd1 vccd1 vccd1 _08387_/Y sky130_fd_sc_hd__nor2_1
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07407_ _07407_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _07408_/B sky130_fd_sc_hd__or2_1
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05599_ _09975_/X _05560_/X _05561_/X _05598_/X vssd1 vssd1 vccd1 vccd1 _05655_/B
+ sky130_fd_sc_hd__o22a_1
X_07338_ _07302_/X _07337_/X _07302_/X _07337_/X vssd1 vssd1 vccd1 vccd1 _07338_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07269_ _07269_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07269_/X sky130_fd_sc_hd__or2_1
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09091_/C sky130_fd_sc_hd__or2_2
X_10280_ _10297_/CLK _10280_/D vssd1 vssd1 vccd1 vccd1 _10280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_0_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10330_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06640_ _10360_/Q vssd1 vssd1 vccd1 vccd1 _06640_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ _08436_/A _06436_/A _08439_/A _06436_/A vssd1 vssd1 vccd1 vccd1 _06571_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08310_ _06272_/A _08305_/Y _08264_/A _08313_/A vssd1 vssd1 vccd1 vccd1 _08310_/X
+ sky130_fd_sc_hd__o211a_1
X_09290_ _09903_/X vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__clkbuf_2
X_05522_ _09989_/X _09991_/X _05489_/Y _05562_/A vssd1 vssd1 vccd1 vccd1 _05558_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08241_ _08241_/A _08241_/B vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__or2_1
X_05453_ _10318_/Q vssd1 vssd1 vccd1 vccd1 _05453_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08172_ _08809_/A vssd1 vssd1 vccd1 vccd1 _08172_/X sky130_fd_sc_hd__buf_2
XFILLER_192_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05384_ _10316_/Q _10315_/Q _10317_/Q vssd1 vssd1 vccd1 vccd1 _05452_/B sky130_fd_sc_hd__and3_1
XFILLER_146_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07123_ _07123_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__or2_1
X_07054_ _07054_/A _07072_/B _07054_/C _07118_/B vssd1 vssd1 vccd1 vccd1 _07054_/X
+ sky130_fd_sc_hd__or4_4
X_06005_ _06032_/A vssd1 vssd1 vccd1 vccd1 _06005_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07956_ _07728_/X _07754_/X _07728_/X _07754_/X vssd1 vssd1 vccd1 vccd1 _07956_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06907_ _06907_/A _06886_/X vssd1 vssd1 vccd1 vccd1 _06909_/A sky130_fd_sc_hd__or2b_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _07879_/X _07883_/X _07879_/X _07883_/X vssd1 vssd1 vccd1 vccd1 _07887_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09626_ _08390_/X _06360_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09626_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06838_ _06837_/A _06837_/B _06855_/B vssd1 vssd1 vccd1 vccd1 _06838_/X sky130_fd_sc_hd__a21bo_1
X_06769_ _10395_/Q _06801_/B _10394_/Q _06800_/B _06768_/X vssd1 vssd1 vccd1 vccd1
+ _06769_/X sky130_fd_sc_hd__a221o_1
X_09557_ _08373_/Y _10117_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__mux2_1
X_08508_ _10066_/Q _08484_/B _08485_/B vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__a21bo_1
XFILLER_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _06606_/X _05012_/A _05013_/X _09487_/X _05468_/X vssd1 vssd1 vccd1 vccd1
+ _10450_/D sky130_fd_sc_hd__o221a_1
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08439_ _08439_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08439_/Y sky130_fd_sc_hd__nor2_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10401_ _10436_/CLK _10401_/D vssd1 vssd1 vccd1 vccd1 _10401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10332_ _10346_/CLK _10332_/D vssd1 vssd1 vccd1 vccd1 _10332_/Q sky130_fd_sc_hd__dfxtp_1
X_10263_ _10300_/CLK _10263_/D vssd1 vssd1 vccd1 vccd1 _10263_/Q sky130_fd_sc_hd__dfxtp_1
X_10194_ _10399_/CLK _10194_/D vssd1 vssd1 vccd1 vccd1 _10194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput12 io_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
XFILLER_190_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 io_wb_dat_i[23] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 io_wb_dat_i[13] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
Xinput45 io_wb_dat_i[4] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_6
XFILLER_182_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08790_ _08790_/A vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07810_ _07811_/A _07897_/B _07811_/C _07864_/A vssd1 vssd1 vccd1 vccd1 _07812_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07741_ _07739_/X _07740_/X _07739_/X _07740_/X vssd1 vssd1 vccd1 vccd1 _07741_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_96_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07672_ _07672_/A _07676_/B _07672_/C vssd1 vssd1 vccd1 vccd1 _07672_/X sky130_fd_sc_hd__or3_1
X_09411_ _09404_/X _09410_/X _09404_/X _09410_/X vssd1 vssd1 vccd1 vccd1 _09411_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06623_ _06623_/A _06795_/A vssd1 vssd1 vccd1 vccd1 _06623_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06554_ _10102_/Q vssd1 vssd1 vccd1 vccd1 _08434_/A sky130_fd_sc_hd__inv_2
X_09342_ _09447_/A _09945_/X _09343_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09344_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05505_ _05505_/A _05505_/B vssd1 vssd1 vccd1 vccd1 _05505_/Y sky130_fd_sc_hd__nor2_4
X_09273_ _09271_/X _09272_/X _09271_/X _09272_/X vssd1 vssd1 vccd1 vccd1 _09273_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06485_ _06495_/A _06484_/X _06495_/A _06484_/X vssd1 vssd1 vccd1 vccd1 _06485_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_08224_ _08765_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__or2_1
XFILLER_119_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05436_ _10322_/Q _05436_/B vssd1 vssd1 vccd1 vccd1 _05436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08155_ _08200_/A vssd1 vssd1 vccd1 vccd1 _08155_/X sky130_fd_sc_hd__buf_2
X_05367_ _05367_/A vssd1 vssd1 vccd1 vccd1 _10332_/D sky130_fd_sc_hd__inv_2
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07106_ _07150_/A _09888_/X vssd1 vssd1 vccd1 vccd1 _07112_/C sky130_fd_sc_hd__nor2_1
X_08086_ _08774_/A vssd1 vssd1 vccd1 vccd1 _08086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05298_ _05298_/A _05362_/A _05298_/C vssd1 vssd1 vccd1 vccd1 _05355_/A sky130_fd_sc_hd__or3_1
X_07037_ _07074_/A _07036_/Y _07074_/A _07036_/Y vssd1 vssd1 vccd1 vccd1 _07037_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08988_ _08988_/A vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__inv_2
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _07935_/X _07936_/X _07937_/X _07938_/X vssd1 vssd1 vccd1 vccd1 _07939_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _10422_/Q _08072_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_33_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10328_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10315_ _10330_/CLK _10315_/D vssd1 vssd1 vccd1 vccd1 _10315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10246_ _10249_/CLK _10246_/D vssd1 vssd1 vccd1 vccd1 _10246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10177_ _10450_/CLK _10177_/D vssd1 vssd1 vccd1 vccd1 _10177_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06270_ _06270_/A _08291_/A vssd1 vssd1 vccd1 vccd1 _06271_/B sky130_fd_sc_hd__or2_1
XFILLER_187_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05221_ _05239_/A vssd1 vssd1 vccd1 vccd1 _05221_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05152_ _05157_/A _05152_/B vssd1 vssd1 vccd1 vccd1 _10402_/D sky130_fd_sc_hd__nor2_1
XFILLER_155_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _10402_/Q _10199_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05083_ _05095_/A vssd1 vssd1 vccd1 vccd1 _05083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _08998_/A _09010_/B _08912_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _08913_/A
+ sky130_fd_sc_hd__o22a_1
X_09891_ _06838_/X _05849_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__mux2_1
X_08842_ _08842_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08842_/Y sky130_fd_sc_hd__nor2_1
X_08773_ _08153_/Y _08770_/Y _08762_/B vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__o21ai_1
X_05985_ _06099_/A vssd1 vssd1 vccd1 vccd1 _05985_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07724_ _07897_/A _07539_/B _07802_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07724_/X
+ sky130_fd_sc_hd__o22a_1
X_07655_ _07676_/A _07677_/A vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__or2_1
XFILLER_198_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06606_ _10450_/Q vssd1 vssd1 vccd1 vccd1 _06606_/X sky130_fd_sc_hd__buf_2
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07586_ _09919_/X vssd1 vssd1 vccd1 vccd1 _07765_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _09323_/X _09324_/X _09323_/X _09324_/X vssd1 vssd1 vccd1 vccd1 _09325_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06537_ _08427_/A _06540_/A _10099_/Q _06463_/A vssd1 vssd1 vccd1 vccd1 _06538_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09256_ _09254_/X _09314_/A _09254_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _09262_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06468_ _06471_/A _06467_/X _06471_/A _06467_/X vssd1 vssd1 vccd1 vccd1 _06468_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ _08545_/A _06249_/B _08206_/Y vssd1 vssd1 vccd1 vccd1 _08207_/X sky130_fd_sc_hd__a21o_1
X_05419_ _05413_/B _05416_/X _05418_/Y _05393_/A _05409_/X vssd1 vssd1 vccd1 vccd1
+ _05420_/A sky130_fd_sc_hd__o32a_1
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09187_ _09187_/A _09187_/B vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__or2_1
X_06399_ _06399_/A vssd1 vssd1 vccd1 vccd1 _06399_/X sky130_fd_sc_hd__buf_1
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08138_ _08782_/A vssd1 vssd1 vccd1 vccd1 _08138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08069_ _08069_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08069_/Y sky130_fd_sc_hd__nor2_1
X_10100_ _10442_/CLK _10100_/D vssd1 vssd1 vccd1 vccd1 _10100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10031_ _10450_/Q _09559_/X _08379_/Y _09560_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10031_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10229_ _10289_/CLK _10229_/D vssd1 vssd1 vccd1 vccd1 _10229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05770_ _05770_/A _10127_/Q vssd1 vssd1 vccd1 vccd1 _05771_/C sky130_fd_sc_hd__nor2_1
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07440_ _10277_/Q _07440_/B vssd1 vssd1 vccd1 vccd1 _07441_/B sky130_fd_sc_hd__or2_1
X_07371_ _07333_/X _07371_/B vssd1 vssd1 vccd1 vccd1 _07371_/X sky130_fd_sc_hd__and2b_1
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09110_ _09043_/A _09109_/X _09043_/A _09109_/X vssd1 vssd1 vccd1 vccd1 _09111_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06322_ _06322_/A vssd1 vssd1 vccd1 vccd1 _06322_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09041_ _09024_/X _09040_/X _09024_/X _09040_/X vssd1 vssd1 vccd1 vccd1 _09057_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_209_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06253_ _06253_/A _06253_/B vssd1 vssd1 vccd1 vccd1 _08222_/A sky130_fd_sc_hd__or2_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06184_ _06184_/A _08325_/A vssd1 vssd1 vccd1 vccd1 _09944_/S sky130_fd_sc_hd__nor2_8
X_05204_ _05202_/X _10384_/Q _05203_/X _09899_/X _05198_/X vssd1 vssd1 vccd1 vccd1
+ _10384_/D sky130_fd_sc_hd__o221a_1
XFILLER_190_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05135_ _05678_/A vssd1 vssd1 vccd1 vccd1 _05157_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05066_ _10433_/Q _05064_/X input33/X _05065_/X _05062_/X vssd1 vssd1 vccd1 vccd1
+ _10433_/D sky130_fd_sc_hd__o221a_1
X_09943_ _10041_/Q input19/X _09943_/S vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__mux2_1
X_09874_ _08308_/Y _10377_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09874_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08825_ _06262_/A _08730_/Y _08824_/X vssd1 vssd1 vccd1 vccd1 _08825_/X sky130_fd_sc_hd__a21bo_1
XINSDIODE2_14 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _08756_/A vssd1 vssd1 vccd1 vccd1 _08756_/Y sky130_fd_sc_hd__inv_2
X_05968_ _05968_/A _08318_/A vssd1 vssd1 vccd1 vccd1 _05971_/A sky130_fd_sc_hd__or2_4
X_08687_ _08294_/A _10072_/Q _08299_/A _10073_/Q vssd1 vssd1 vccd1 vccd1 _08695_/B
+ sky130_fd_sc_hd__a22o_1
X_05899_ _10248_/Q _05896_/X input24/X _05897_/X _05885_/X vssd1 vssd1 vccd1 vccd1
+ _10248_/D sky130_fd_sc_hd__o221a_1
X_07707_ _07707_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _07707_/X sky130_fd_sc_hd__or2_1
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07638_ _07621_/A _07627_/A _07621_/Y vssd1 vssd1 vccd1 vccd1 _07638_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07569_ _07564_/X _07568_/X _07564_/X _07568_/X vssd1 vssd1 vccd1 vccd1 _07569_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09308_ _09286_/X _09307_/X _09286_/X _09307_/X vssd1 vssd1 vccd1 vccd1 _09308_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _09238_/A _09238_/B _09303_/A vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10014_ _08012_/A _08050_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10014_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06940_ _06881_/X _06939_/X _06881_/X _06939_/X vssd1 vssd1 vccd1 vccd1 _06940_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06871_ _06911_/B vssd1 vssd1 vccd1 vccd1 _06949_/D sky130_fd_sc_hd__clkbuf_2
X_08610_ _06271_/A _08496_/Y _08609_/Y vssd1 vssd1 vccd1 vccd1 _08610_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05822_ _07445_/A _05795_/Y _05796_/X _05821_/X vssd1 vssd1 vccd1 vccd1 _05822_/X
+ sky130_fd_sc_hd__o22a_1
X_09590_ _08431_/Y _08430_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__mux2_2
X_08541_ _10054_/Q _08472_/B _08473_/B vssd1 vssd1 vccd1 vccd1 _08542_/A sky130_fd_sc_hd__a21bo_1
X_05753_ _05761_/A vssd1 vssd1 vccd1 vccd1 _05753_/X sky130_fd_sc_hd__clkbuf_2
X_08472_ _10054_/Q _08472_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__or2_1
X_05684_ _05684_/A vssd1 vssd1 vccd1 vccd1 _05684_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07423_ _07423_/A vssd1 vssd1 vccd1 vccd1 _07423_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _07350_/X _07351_/X _07350_/X _07351_/X vssd1 vssd1 vccd1 vccd1 _07358_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06305_ _06305_/A vssd1 vssd1 vccd1 vccd1 _06305_/Y sky130_fd_sc_hd__inv_2
X_07285_ _07188_/X _07199_/X _07188_/X _07199_/X vssd1 vssd1 vccd1 vccd1 _07285_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_191_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06236_ _10039_/Q vssd1 vssd1 vccd1 vccd1 _06236_/Y sky130_fd_sc_hd__inv_2
X_09024_ _08997_/X _09004_/X _09005_/X _09006_/X vssd1 vssd1 vccd1 vccd1 _09024_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06167_ _06169_/A _09675_/X vssd1 vssd1 vccd1 vccd1 _10124_/D sky130_fd_sc_hd__and2_1
X_05118_ _10441_/Q vssd1 vssd1 vccd1 vccd1 _05118_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06098_ _10340_/Q _06093_/X _10168_/Q _06094_/X _05985_/X vssd1 vssd1 vccd1 vccd1
+ _10168_/D sky130_fd_sc_hd__a221o_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05049_ _10442_/Q _05047_/X input43/X _05048_/X _05036_/X vssd1 vssd1 vccd1 vccd1
+ _10442_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09926_ _09925_/X _09447_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09926_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09857_ _09856_/X input36/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09857_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08808_ _08808_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__and2_1
X_09788_ _09787_/X _08212_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09788_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08739_ _06635_/Y _08738_/Y _08734_/X vssd1 vssd1 vccd1 vccd1 _08739_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07070_ _07055_/X _07057_/Y _07055_/X _07057_/Y vssd1 vssd1 vccd1 vccd1 _07070_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06021_ _09857_/X _06015_/X _06020_/X _06017_/X _06018_/X vssd1 vssd1 vccd1 vccd1
+ _10201_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09711_ _10447_/Q _06647_/Y _09717_/S vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07972_ _07960_/X _07965_/X _07966_/X _07971_/X vssd1 vssd1 vccd1 vccd1 _07972_/X
+ sky130_fd_sc_hd__o22a_1
X_06923_ _06923_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _06924_/B sky130_fd_sc_hd__or2_1
X_09642_ _06393_/X _06395_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__mux2_1
X_06854_ _06942_/C vssd1 vssd1 vccd1 vccd1 _06961_/A sky130_fd_sc_hd__clkbuf_2
X_06785_ _06614_/C _06698_/A _06614_/B _06694_/Y _06784_/Y vssd1 vssd1 vccd1 vccd1
+ _06785_/X sky130_fd_sc_hd__o221a_1
X_09573_ _08403_/Y _10123_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__mux2_1
X_05805_ _05805_/A vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__buf_2
X_08524_ _10065_/Q vssd1 vssd1 vccd1 vccd1 _08524_/Y sky130_fd_sc_hd__inv_2
X_05736_ _10268_/Q vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__buf_2
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ _10049_/Q vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__inv_2
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05667_ _05667_/A vssd1 vssd1 vccd1 vccd1 _05667_/Y sky130_fd_sc_hd__inv_2
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05598_ _09946_/X _05564_/X _05662_/A vssd1 vssd1 vccd1 vccd1 _05598_/X sky130_fd_sc_hd__o21a_1
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _07406_/A _07406_/B vssd1 vssd1 vccd1 vccd1 _07407_/B sky130_fd_sc_hd__or2_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08386_ _08386_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__or2_1
XFILLER_211_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07337_ _07263_/X _07337_/B vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__and2b_1
XFILLER_176_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07269_/B sky130_fd_sc_hd__nor2_1
XFILLER_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06219_ _09689_/X _06217_/X _10090_/Q _06218_/X vssd1 vssd1 vccd1 vccd1 _10090_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09007_ _09005_/X _09006_/X _09005_/X _09006_/X vssd1 vssd1 vccd1 vccd1 _09007_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07199_ _07191_/X _07194_/X _07197_/X _07198_/X vssd1 vssd1 vccd1 vccd1 _07199_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09909_ _08355_/X _06299_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06570_ _08442_/A _06435_/A _10105_/Q _06465_/A vssd1 vssd1 vccd1 vccd1 _06570_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05521_ _10012_/X _09990_/X _05490_/X _05520_/X vssd1 vssd1 vccd1 vccd1 _05562_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08240_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08240_/X sky130_fd_sc_hd__clkbuf_4
X_05452_ _10318_/Q _05452_/B vssd1 vssd1 vccd1 vccd1 _05452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08171_ _08245_/A vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05383_ _10319_/Q vssd1 vssd1 vccd1 vccd1 _05386_/A sky130_fd_sc_hd__inv_2
X_07122_ _07111_/A _07111_/B _07111_/X vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__a21bo_1
XFILLER_118_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ _07054_/A _07072_/B _07054_/C _07118_/B vssd1 vssd1 vccd1 vccd1 _07055_/A
+ sky130_fd_sc_hd__o22a_1
X_06004_ _06070_/A vssd1 vssd1 vccd1 vccd1 _06032_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07955_ _07849_/A _07849_/B _07850_/B vssd1 vssd1 vccd1 vccd1 _07955_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06906_ _06911_/A _09893_/X _07100_/A _06911_/B vssd1 vssd1 vccd1 vccd1 _06907_/A
+ sky130_fd_sc_hd__o22a_1
X_09625_ _09624_/X _07806_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09625_/X sky130_fd_sc_hd__mux2_1
X_07886_ _07886_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__or2_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06837_ _06837_/A _06837_/B vssd1 vssd1 vccd1 vccd1 _06855_/B sky130_fd_sc_hd__or2_1
X_06768_ _10393_/Q _06799_/B _10394_/Q _06800_/B _06767_/X vssd1 vssd1 vccd1 vccd1
+ _06768_/X sky130_fd_sc_hd__o221a_1
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09555_/X _10353_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09556_/X sky130_fd_sc_hd__mux2_1
X_08507_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__nand2_1
XFILLER_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06699_ _10374_/Q vssd1 vssd1 vccd1 vccd1 _06699_/Y sky130_fd_sc_hd__inv_2
X_09487_ _05016_/A _05016_/B _09486_/Y input48/X _05016_/Y vssd1 vssd1 vccd1 vccd1
+ _09487_/X sky130_fd_sc_hd__o32a_1
XFILLER_102_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05719_ _05761_/A vssd1 vssd1 vccd1 vccd1 _05719_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08438_ _09982_/X _08449_/B vssd1 vssd1 vccd1 vccd1 _08438_/Y sky130_fd_sc_hd__nor2_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _09310_/A vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__buf_4
XFILLER_137_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10400_ _10433_/CLK _10400_/D vssd1 vssd1 vccd1 vccd1 _10400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _10346_/CLK _10331_/D vssd1 vssd1 vccd1 vccd1 _10331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _10300_/CLK _10262_/D vssd1 vssd1 vccd1 vccd1 _10262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10193_ _10399_/CLK _10193_/D vssd1 vssd1 vccd1 vccd1 _10193_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 io_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput35 io_wb_dat_i[24] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput24 io_wb_dat_i[14] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_6
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput46 io_wb_dat_i[5] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_6
XFILLER_128_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07740_ _07698_/A _07698_/B _07699_/B vssd1 vssd1 vccd1 vccd1 _07740_/X sky130_fd_sc_hd__a21bo_1
XFILLER_203_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07671_/X sky130_fd_sc_hd__or2_1
XFILLER_203_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09410_ _09409_/A _09409_/B _09409_/Y vssd1 vssd1 vccd1 vccd1 _09410_/X sky130_fd_sc_hd__a21o_1
X_06622_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06553_ _06560_/C _06552_/X _06560_/C _06552_/X vssd1 vssd1 vccd1 vccd1 _06553_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_09341_ _09341_/A _09340_/X vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__or2b_1
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05504_ _10250_/Q vssd1 vssd1 vccd1 vccd1 _05505_/B sky130_fd_sc_hd__inv_2
XFILLER_178_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _09171_/X _09177_/X _09178_/X _09212_/X vssd1 vssd1 vccd1 vccd1 _09272_/X
+ sky130_fd_sc_hd__o22a_1
X_06484_ _06495_/C _06484_/B vssd1 vssd1 vccd1 vccd1 _06484_/X sky130_fd_sc_hd__and2_1
X_08223_ _06253_/A _06253_/B _08222_/Y vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__a21o_1
X_05435_ _05435_/A vssd1 vssd1 vccd1 vccd1 _05436_/B sky130_fd_sc_hd__inv_2
X_08154_ _10181_/Q vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__inv_2
X_05366_ _05362_/Y _05333_/A _05365_/Y _05336_/A _05296_/A vssd1 vssd1 vccd1 vccd1
+ _05367_/A sky130_fd_sc_hd__o32a_1
XFILLER_161_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08085_ _08211_/A vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__inv_2
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07105_ _07103_/X _07104_/X _07103_/X _07104_/X vssd1 vssd1 vccd1 vccd1 _07111_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_05297_ _10334_/Q vssd1 vssd1 vccd1 vccd1 _05298_/C sky130_fd_sc_hd__inv_2
X_07036_ _07011_/X _07035_/X _07011_/X _07035_/X vssd1 vssd1 vccd1 vccd1 _07036_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08987_ _08851_/X _08863_/X _08851_/X _08863_/X vssd1 vssd1 vccd1 vccd1 _08988_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07938_ _07935_/X _07936_/X _07935_/X _07936_/X vssd1 vssd1 vccd1 vccd1 _07938_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07869_ _07869_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _10421_/Q _08071_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09608_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _09538_/X _10348_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09539_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ _10422_/CLK _10314_/D vssd1 vssd1 vccd1 vccd1 _10314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10245_ _10249_/CLK _10245_/D vssd1 vssd1 vccd1 vccd1 _10245_/Q sky130_fd_sc_hd__dfxtp_1
X_10176_ _10176_/CLK _10176_/D vssd1 vssd1 vccd1 vccd1 _10176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05220_ _10376_/Q _05215_/X input40/X _05216_/X _05218_/X vssd1 vssd1 vccd1 vccd1
+ _10376_/D sky130_fd_sc_hd__o221a_1
X_05151_ _05129_/X _06616_/A _05150_/Y _05138_/X vssd1 vssd1 vccd1 vccd1 _05152_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05082_ _05094_/A vssd1 vssd1 vccd1 vccd1 _05082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ _08908_/Y _08907_/X _08930_/A vssd1 vssd1 vccd1 vccd1 _08910_/Y sky130_fd_sc_hd__o21ai_1
X_09890_ _06833_/X _05876_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09890_/X sky130_fd_sc_hd__mux2_2
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08841_ _10296_/Q vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__inv_2
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08772_ _08772_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05984_ _10210_/Q vssd1 vssd1 vccd1 vccd1 _07854_/D sky130_fd_sc_hd__clkbuf_2
X_07723_ _07720_/X _07722_/X _07720_/X _07722_/X vssd1 vssd1 vccd1 vccd1 _07723_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07654_ _07581_/X _07652_/X _07537_/X _07653_/X vssd1 vssd1 vccd1 vccd1 _07654_/X
+ sky130_fd_sc_hd__o211a_1
X_06605_ _05018_/X _06739_/A _05024_/X _06600_/Y _06604_/X vssd1 vssd1 vccd1 vccd1
+ _06605_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07585_ _07585_/A _07584_/X vssd1 vssd1 vccd1 vccd1 _07585_/X sky130_fd_sc_hd__or2b_1
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _09244_/A _09267_/X _09269_/B vssd1 vssd1 vccd1 vccd1 _09324_/X sky130_fd_sc_hd__o21a_1
X_06536_ _06536_/A vssd1 vssd1 vccd1 vccd1 _06540_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ _09354_/C _09258_/B _09104_/A _09202_/A _09203_/A vssd1 vssd1 vccd1 vccd1
+ _09314_/A sky130_fd_sc_hd__o32a_1
X_06467_ _10085_/Q _06466_/X _06454_/X _06456_/Y vssd1 vssd1 vccd1 vccd1 _06467_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08206_ _08206_/A vssd1 vssd1 vccd1 vccd1 _08206_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05418_ _10326_/Q _05418_/B vssd1 vssd1 vccd1 vccd1 _05418_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09186_ _09185_/A _09185_/B _09185_/X vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__a21bo_1
X_06398_ _10248_/Q _08409_/A _06397_/Y _10141_/Q vssd1 vssd1 vccd1 vccd1 _06399_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ _08137_/A vssd1 vssd1 vccd1 vccd1 _08782_/A sky130_fd_sc_hd__clkbuf_2
X_05349_ _05344_/B _05333_/X _05348_/Y _05336_/X _05301_/A vssd1 vssd1 vccd1 vccd1
+ _05350_/A sky130_fd_sc_hd__o32a_1
XFILLER_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08068_ _08075_/B _10306_/Q vssd1 vssd1 vccd1 vccd1 _08068_/Y sky130_fd_sc_hd__nor2b_1
X_07019_ _07019_/A vssd1 vssd1 vccd1 vccd1 _07019_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10030_ _10449_/Q _09556_/X _08372_/Y _09557_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10030_/X sky130_fd_sc_hd__mux4_2
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10228_ _10289_/CLK _10228_/D vssd1 vssd1 vccd1 vccd1 _10228_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _10346_/CLK _10159_/D vssd1 vssd1 vccd1 vccd1 _10159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07370_ _07326_/X _07363_/X _07326_/X _07363_/X vssd1 vssd1 vccd1 vccd1 _07386_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_203_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06321_ _10240_/Q _08370_/A _06320_/Y _10133_/Q vssd1 vssd1 vccd1 vccd1 _06322_/A
+ sky130_fd_sc_hd__o22a_2
X_06252_ _10186_/Q _08213_/A vssd1 vssd1 vccd1 vccd1 _06253_/B sky130_fd_sc_hd__or2_1
X_09040_ _09037_/X _09039_/X _09037_/X _09039_/X vssd1 vssd1 vccd1 vccd1 _09040_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05203_ _05203_/A vssd1 vssd1 vccd1 vccd1 _05203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06183_ _06183_/A _08324_/C _08324_/B vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__or3_4
XFILLER_171_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05134_ input52/X vssd1 vssd1 vccd1 vccd1 _05678_/A sky130_fd_sc_hd__clkbuf_4
X_05065_ _05073_/A vssd1 vssd1 vccd1 vccd1 _05065_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09942_ _09941_/X _10040_/Q _09944_/S vssd1 vssd1 vccd1 vccd1 _09942_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09873_ _09872_/X input40/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__mux2_1
X_08824_ _08824_/A _08824_/B _08824_/C vssd1 vssd1 vccd1 vccd1 _08824_/X sky130_fd_sc_hd__or3_2
XINSDIODE2_15 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08755_ _08753_/A _08753_/B _08753_/Y vssd1 vssd1 vccd1 vccd1 _08756_/A sky130_fd_sc_hd__a21oi_2
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05967_ _05967_/A _06137_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__or2_4
X_07706_ _07706_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07707_/B sky130_fd_sc_hd__nor2_1
X_08686_ _10206_/Q _08454_/Y _06000_/A _08613_/Y vssd1 vssd1 vccd1 vccd1 _08695_/A
+ sky130_fd_sc_hd__a22o_1
X_05898_ _10249_/Q _05896_/X input25/X _05897_/X _05885_/X vssd1 vssd1 vccd1 vccd1
+ _10249_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10225_/CLK sky130_fd_sc_hd__clkbuf_16
X_07637_ _10210_/Q _07566_/B _07820_/A _07634_/Y _07636_/X vssd1 vssd1 vccd1 vccd1
+ _07637_/X sky130_fd_sc_hd__a41o_1
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07568_ _07558_/C _07567_/A _07557_/A _07567_/Y vssd1 vssd1 vccd1 vccd1 _07568_/X
+ sky130_fd_sc_hd__a22o_1
X_09307_ _09288_/X _09306_/X _09288_/X _09306_/X vssd1 vssd1 vccd1 vccd1 _09307_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06519_ _06519_/A _06519_/B vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__or2_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07499_ _07485_/X _07488_/X _07496_/X _07498_/X vssd1 vssd1 vccd1 vccd1 _07499_/X
+ sky130_fd_sc_hd__o22a_1
X_09238_ _09238_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__nor2_2
XFILLER_166_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _09168_/A _09168_/C _09168_/B vssd1 vssd1 vccd1 vccd1 _09170_/C sky130_fd_sc_hd__o21ai_1
XFILLER_119_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10013_ _08037_/X _07390_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _10013_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06870_ _07028_/B vssd1 vssd1 vccd1 vccd1 _06870_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05821_ _05797_/Y _05798_/Y _05799_/X _05820_/X vssd1 vssd1 vccd1 vccd1 _05821_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08540_ _10055_/Q _08473_/B _08474_/B vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__a21boi_1
X_05752_ _05788_/A _05751_/X _09639_/X _05743_/X _05747_/X vssd1 vssd1 vccd1 vccd1
+ _10277_/D sky130_fd_sc_hd__o221a_1
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _10053_/Q _08471_/B vssd1 vssd1 vccd1 vccd1 _08472_/B sky130_fd_sc_hd__or2_1
X_05683_ _08618_/A _05683_/B vssd1 vssd1 vccd1 vccd1 _10302_/D sky130_fd_sc_hd__nor2_1
XFILLER_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07422_ _07421_/A _07417_/B _07418_/B vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__a21bo_1
XFILLER_210_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _07347_/X _07352_/X _07347_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07353_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06304_ _06304_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06305_/A sky130_fd_sc_hd__or2_1
X_07284_ _07283_/A _07283_/B _07283_/X vssd1 vssd1 vccd1 vccd1 _07296_/A sky130_fd_sc_hd__a21boi_2
XFILLER_191_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06235_ _06235_/A vssd1 vssd1 vccd1 vccd1 _06235_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09023_ _09022_/A _09022_/B _09067_/A vssd1 vssd1 vccd1 vccd1 _09023_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_191_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06166_ _06169_/A _09676_/X vssd1 vssd1 vccd1 vccd1 _10125_/D sky130_fd_sc_hd__and2_1
X_05117_ _10409_/Q vssd1 vssd1 vccd1 vccd1 _06614_/B sky130_fd_sc_hd__inv_2
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06097_ _10341_/Q _06093_/X _10169_/Q _06094_/X _05985_/X vssd1 vssd1 vccd1 vccd1
+ _10169_/D sky130_fd_sc_hd__a221o_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05048_ _05073_/A vssd1 vssd1 vccd1 vccd1 _05048_/X sky130_fd_sc_hd__clkbuf_4
X_09925_ _08343_/X _06281_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09925_/X sky130_fd_sc_hd__mux2_1
X_09856_ _09855_/X _08287_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09856_/X sky130_fd_sc_hd__mux2_1
X_08807_ _08823_/C _08806_/Y vssd1 vssd1 vccd1 vccd1 _08808_/B sky130_fd_sc_hd__or2b_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09787_ _10355_/Q _09786_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09787_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06999_ _07116_/B vssd1 vssd1 vccd1 vccd1 _06999_/Y sky130_fd_sc_hd__inv_2
X_08738_ _08738_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08738_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08669_ _06265_/A _08505_/Y _06026_/X _08668_/Y vssd1 vssd1 vccd1 vccd1 _08674_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06020_ _10201_/Q vssd1 vssd1 vccd1 vccd1 _06020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _07971_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _07971_/X sky130_fd_sc_hd__or2_1
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09710_ _06623_/Y _10379_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10045_/D sky130_fd_sc_hd__mux2_1
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06922_ _06898_/C _06895_/B _06895_/Y vssd1 vssd1 vccd1 vccd1 _06923_/B sky130_fd_sc_hd__o21ai_1
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09641_ _06385_/Y _06386_/Y _10175_/Q vssd1 vssd1 vccd1 vccd1 _09641_/X sky130_fd_sc_hd__mux2_2
X_06853_ _07112_/A vssd1 vssd1 vccd1 vccd1 _06942_/C sky130_fd_sc_hd__clkbuf_2
X_06784_ _10407_/Q _06815_/B _10408_/Q _06816_/B _06783_/X vssd1 vssd1 vccd1 vccd1
+ _06784_/Y sky130_fd_sc_hd__o221ai_1
X_09572_ _08400_/X _09571_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__mux2_2
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05804_ _05804_/A vssd1 vssd1 vccd1 vccd1 _05805_/A sky130_fd_sc_hd__inv_2
X_08523_ _08514_/Y _08517_/X _08520_/Y _08596_/C vssd1 vssd1 vccd1 vccd1 _08523_/X
+ sky130_fd_sc_hd__o22a_1
X_05735_ _10285_/Q _05728_/X _07421_/A _05732_/X _05724_/X vssd1 vssd1 vccd1 vccd1
+ _10285_/D sky130_fd_sc_hd__o221a_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _10075_/Q vssd1 vssd1 vccd1 vccd1 _08454_/Y sky130_fd_sc_hd__inv_2
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05666_ _05677_/A _05666_/B vssd1 vssd1 vccd1 vccd1 _10305_/D sky130_fd_sc_hd__nor2_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08385_ _08385_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08385_/Y sky130_fd_sc_hd__nor2_1
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05597_ _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05662_/A sky130_fd_sc_hd__nand2_1
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07405_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07406_/B sky130_fd_sc_hd__or2_1
X_07336_ _07035_/X _07335_/X _07035_/X _07335_/X vssd1 vssd1 vccd1 vccd1 _07336_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09006_ _08962_/X _08975_/X _08945_/X _08976_/X vssd1 vssd1 vccd1 vccd1 _09006_/X
+ sky130_fd_sc_hd__o22a_1
X_07267_ _07241_/A _07247_/A _07241_/Y vssd1 vssd1 vccd1 vccd1 _07267_/X sky130_fd_sc_hd__a21o_1
X_06218_ _06225_/A vssd1 vssd1 vccd1 vccd1 _06218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07198_ _07191_/X _07194_/X _07191_/X _07194_/X vssd1 vssd1 vccd1 vccd1 _07198_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06149_ _06157_/A vssd1 vssd1 vccd1 vccd1 _06149_/X sky130_fd_sc_hd__buf_1
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09908_ _05782_/X _07460_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09908_/X sky130_fd_sc_hd__mux2_1
X_09839_ _10368_/Q _09838_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09839_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05520_ _10014_/X _10017_/X _05491_/X _05519_/X vssd1 vssd1 vccd1 vccd1 _05520_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05451_ _05451_/A vssd1 vssd1 vccd1 vccd1 _10319_/D sky130_fd_sc_hd__inv_2
X_08170_ _10192_/Q vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__inv_2
XFILLER_192_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05382_ _10320_/Q vssd1 vssd1 vccd1 vccd1 _05387_/A sky130_fd_sc_hd__inv_2
X_07121_ _07121_/A _07102_/X vssd1 vssd1 vccd1 vccd1 _07123_/A sky130_fd_sc_hd__or2b_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07052_ _07052_/A _07052_/B vssd1 vssd1 vccd1 vccd1 _07052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06003_ _10444_/Q input5/X input52/X vssd1 vssd1 vccd1 vccd1 _06070_/A sky130_fd_sc_hd__a21oi_4
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07954_ _07950_/X _07951_/X _07950_/X _07951_/X vssd1 vssd1 vccd1 vccd1 _07954_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07885_ _07885_/A _07885_/B _07885_/C _07885_/D vssd1 vssd1 vccd1 vccd1 _07886_/B
+ sky130_fd_sc_hd__and4_1
X_06905_ _06901_/X _06904_/X _06901_/X _06904_/X vssd1 vssd1 vccd1 vccd1 _06905_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09624_ _09623_/X _07054_/C _09999_/S vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06836_ _06836_/A _06836_/B vssd1 vssd1 vccd1 vccd1 _06837_/B sky130_fd_sc_hd__or2_1
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06767_ _10393_/Q _06799_/B _10392_/Q _06798_/B _06766_/X vssd1 vssd1 vccd1 vccd1
+ _06767_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09555_ _10385_/Q _10182_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09555_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ _08505_/Y _08502_/Y _08487_/B vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__o21ai_1
X_06698_ _06698_/A vssd1 vssd1 vccd1 vccd1 _06816_/B sky130_fd_sc_hd__inv_2
X_09486_ input48/X vssd1 vssd1 vccd1 vccd1 _09486_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05718_ _05718_/A vssd1 vssd1 vccd1 vccd1 _05761_/A sky130_fd_sc_hd__buf_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _08453_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__clkbuf_2
X_05649_ _05649_/A _05649_/B vssd1 vssd1 vccd1 vccd1 _05649_/Y sky130_fd_sc_hd__nor2_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08368_ _09259_/A vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__buf_1
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08304_/B sky130_fd_sc_hd__or2_2
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07319_ _07317_/X _07318_/X _07317_/X _07318_/X vssd1 vssd1 vccd1 vccd1 _07319_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10330_ _10330_/CLK _10330_/D vssd1 vssd1 vccd1 vccd1 _10330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10261_ _10300_/CLK _10261_/D vssd1 vssd1 vccd1 vccd1 _10261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _10436_/CLK _10192_/D vssd1 vssd1 vccd1 vccd1 _10192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput36 io_wb_dat_i[25] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput25 io_wb_dat_i[15] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_6
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 io_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput47 io_wb_dat_i[6] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_6
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ _07663_/A _07765_/A _07660_/A _07672_/A _07669_/Y vssd1 vssd1 vccd1 vccd1
+ _07671_/B sky130_fd_sc_hd__o41a_1
XFILLER_203_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06621_ _06621_/A vssd1 vssd1 vccd1 vccd1 _06623_/A sky130_fd_sc_hd__inv_2
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06552_ _06560_/A _06560_/B _06543_/Y _06551_/X vssd1 vssd1 vccd1 vccd1 _06552_/X
+ sky130_fd_sc_hd__o31a_1
X_09340_ _09457_/C _09922_/X _09468_/A _09903_/X vssd1 vssd1 vccd1 vccd1 _09340_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_92_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09242_/X _09270_/X _09242_/X _09270_/X vssd1 vssd1 vccd1 vccd1 _09271_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05503_ _05505_/A vssd1 vssd1 vccd1 vccd1 _05510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_166_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08222_ _08222_/A vssd1 vssd1 vccd1 vccd1 _08222_/Y sky130_fd_sc_hd__inv_2
X_06483_ _08385_/A _06432_/A _08388_/A _06432_/A vssd1 vssd1 vccd1 vccd1 _06484_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05434_ _05434_/A vssd1 vssd1 vccd1 vccd1 _10323_/D sky130_fd_sc_hd__inv_2
X_08153_ _08761_/A vssd1 vssd1 vccd1 vccd1 _08153_/Y sky130_fd_sc_hd__inv_2
X_05365_ _10332_/Q _10331_/Q vssd1 vssd1 vccd1 vccd1 _05365_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _10358_/Q vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07104_ _07155_/A _09888_/X vssd1 vssd1 vccd1 vccd1 _07104_/X sky130_fd_sc_hd__or2_1
XFILLER_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05296_ _05296_/A _05296_/B vssd1 vssd1 vccd1 vccd1 _05362_/A sky130_fd_sc_hd__or2_2
X_07035_ _06995_/A _06995_/B _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _07035_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_161_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08985_/A _08985_/B _09018_/A vssd1 vssd1 vccd1 vccd1 _08986_/X sky130_fd_sc_hd__a21bo_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07937_ _07760_/A _07760_/B _07761_/B vssd1 vssd1 vccd1 vccd1 _07937_/X sky130_fd_sc_hd__a21bo_1
XFILLER_180_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07868_ _07868_/A _07868_/B _07867_/X vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__or3b_1
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09607_ _10420_/Q _08070_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09607_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06819_ _07152_/D _06819_/B vssd1 vssd1 vccd1 vccd1 _06820_/B sky130_fd_sc_hd__or2_1
X_07799_ _07867_/B vssd1 vssd1 vccd1 vccd1 _07885_/D sky130_fd_sc_hd__inv_2
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09538_ _10380_/Q _10177_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09538_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _09396_/X _09403_/X _09404_/X _09410_/X vssd1 vssd1 vccd1 vccd1 _09469_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10313_ _10426_/CLK _10313_/D vssd1 vssd1 vccd1 vccd1 _10313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10244_ _10244_/CLK _10244_/D vssd1 vssd1 vccd1 vccd1 _10244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10175_ _10244_/CLK _10175_/D vssd1 vssd1 vccd1 vccd1 _10175_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05150_ _10434_/Q vssd1 vssd1 vccd1 vccd1 _05150_/Y sky130_fd_sc_hd__inv_2
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05081_ _10422_/Q _05094_/A input21/X _05095_/A _05078_/X vssd1 vssd1 vccd1 vccd1
+ _10422_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ _10297_/Q _05782_/X _10297_/Q _07854_/A vssd1 vssd1 vccd1 vccd1 _08840_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08771_ _08760_/A _08760_/B _08770_/Y vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__a21oi_2
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05983_ _07820_/A _05970_/A input30/X _05971_/A _05978_/X vssd1 vssd1 vccd1 vccd1
+ _10211_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07722_ _07722_/A _07722_/B vssd1 vssd1 vccd1 vccd1 _07722_/X sky130_fd_sc_hd__or2_1
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07653_ _07555_/X _07558_/X _07559_/X _07580_/X vssd1 vssd1 vccd1 vccd1 _07653_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06604_ _06603_/X _10380_/Q _05024_/X _06600_/Y vssd1 vssd1 vccd1 vccd1 _06604_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _09309_/X _09322_/Y _09309_/X _09322_/Y vssd1 vssd1 vccd1 vccd1 _09323_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07584_ _07603_/A _09920_/X _07587_/D _09921_/X vssd1 vssd1 vccd1 vccd1 _07584_/X
+ sky130_fd_sc_hd__or4_4
X_06535_ _10099_/Q vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__inv_2
XFILLER_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06466_ _06466_/A vssd1 vssd1 vccd1 vccd1 _06466_/X sky130_fd_sc_hd__buf_2
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09254_ _05933_/X _09251_/X _09252_/X _09253_/Y vssd1 vssd1 vccd1 vccd1 _09254_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08205_ _08797_/A _08201_/Y _08208_/B _08188_/X vssd1 vssd1 vccd1 vccd1 _08205_/X
+ sky130_fd_sc_hd__o211a_1
X_09185_ _09185_/A _09185_/B vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__or2_1
X_05417_ _05417_/A vssd1 vssd1 vccd1 vccd1 _05418_/B sky130_fd_sc_hd__inv_2
XFILLER_193_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08136_ _10373_/Q _08134_/X _06624_/Y _06000_/A _08135_/X vssd1 vssd1 vccd1 vccd1
+ _08143_/C sky130_fd_sc_hd__o221a_1
X_06397_ _10248_/Q vssd1 vssd1 vccd1 vccd1 _06397_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05348_ _10337_/Q _05348_/B vssd1 vssd1 vccd1 vccd1 _05348_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05279_ _09897_/X vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__inv_2
X_08067_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_122_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07018_ _10220_/Q _06929_/Y _05964_/X _06930_/Y _06937_/Y vssd1 vssd1 vccd1 vccd1
+ _07019_/A sky130_fd_sc_hd__a41o_1
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _08967_/X _08968_/Y _08967_/X _08968_/Y vssd1 vssd1 vccd1 vccd1 _08970_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _10289_/CLK _10227_/D vssd1 vssd1 vccd1 vccd1 _10227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10158_ _10328_/CLK _10158_/D vssd1 vssd1 vccd1 vccd1 _10158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10089_ _10346_/CLK _10089_/D vssd1 vssd1 vccd1 vccd1 _10089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06320_ _10240_/Q vssd1 vssd1 vccd1 vccd1 _06320_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06251_ _10185_/Q _06251_/B vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__or2_1
XFILLER_175_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05202_ _05202_/A vssd1 vssd1 vccd1 vccd1 _05202_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06182_ _06182_/A _09661_/X vssd1 vssd1 vccd1 vccd1 _10111_/D sky130_fd_sc_hd__and2_1
XFILLER_209_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05133_ _05133_/A _05133_/B vssd1 vssd1 vccd1 vccd1 _10406_/D sky130_fd_sc_hd__nor2_1
XFILLER_171_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05064_ _05072_/A vssd1 vssd1 vccd1 vccd1 _05064_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _10040_/Q input30/X _09943_/S vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09872_ _09871_/X _08306_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09872_/X sky130_fd_sc_hd__mux2_1
X_08823_ _08823_/A _08823_/B _08823_/C _08808_/A vssd1 vssd1 vccd1 vccd1 _08824_/B
+ sky130_fd_sc_hd__or4b_4
XINSDIODE2_16 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ _06640_/Y _08753_/Y _08748_/Y vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__o21bai_1
X_05966_ _10217_/Q vssd1 vssd1 vccd1 vccd1 _05966_/X sky130_fd_sc_hd__buf_2
X_07705_ _07654_/X _07702_/X _07703_/X _07704_/X vssd1 vssd1 vccd1 vccd1 _07705_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08685_ _06265_/A _08505_/Y _08674_/A _08684_/X vssd1 vssd1 vccd1 vccd1 _08685_/X
+ sky130_fd_sc_hd__o22a_1
X_05897_ _05911_/A vssd1 vssd1 vccd1 vccd1 _05897_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07636_ _07877_/A _07539_/B _07815_/A _07634_/A vssd1 vssd1 vccd1 vccd1 _07636_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07567_ _07567_/A vssd1 vssd1 vccd1 vccd1 _07567_/Y sky130_fd_sc_hd__inv_2
X_09306_ _09291_/X _09305_/X _09291_/X _09305_/X vssd1 vssd1 vccd1 vccd1 _09306_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06518_ _06498_/A _06516_/X _06498_/B _06517_/X vssd1 vssd1 vccd1 vccd1 _06519_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09235_/X _09297_/A _09235_/X _09297_/A vssd1 vssd1 vccd1 vccd1 _09238_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _07802_/A _07558_/B _07498_/C vssd1 vssd1 vccd1 vccd1 _07498_/X sky130_fd_sc_hd__or3_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06449_ _10084_/Q vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__inv_2
XFILLER_181_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09168_ _09168_/A _09168_/B _09168_/C vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__or3_1
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08119_ _08119_/A _08119_/B _08119_/C _08119_/D vssd1 vssd1 vccd1 vccd1 _08176_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ _09093_/X _09098_/X _09093_/X _09098_/X vssd1 vssd1 vccd1 vccd1 _09192_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_119_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ _08011_/A _08048_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10012_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05820_ _05801_/X _05802_/Y _05803_/X _05819_/X vssd1 vssd1 vccd1 vccd1 _05820_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05751_ _05871_/A vssd1 vssd1 vccd1 vccd1 _05751_/X sky130_fd_sc_hd__buf_1
X_08470_ _10052_/Q _08470_/B vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__or2_1
X_05682_ _05653_/X _05679_/Y _05680_/Y _08062_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05683_/B sky130_fd_sc_hd__o32a_1
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _07421_/A vssd1 vssd1 vccd1 vccd1 _07421_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07352_ _06984_/X _07349_/X _07350_/X _07351_/X vssd1 vssd1 vccd1 vccd1 _07352_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06303_ _06285_/X _06294_/A _06302_/X vssd1 vssd1 vccd1 vccd1 _06304_/B sky130_fd_sc_hd__o21ba_1
X_07283_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__or2_1
X_06234_ _10036_/Q _06233_/Y _10036_/Q _06233_/Y vssd1 vssd1 vccd1 vccd1 _06235_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__nand2_1
X_06165_ _06169_/A _09677_/X vssd1 vssd1 vccd1 vccd1 _10126_/D sky130_fd_sc_hd__and2_1
XFILLER_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05116_ _05202_/A vssd1 vssd1 vccd1 vccd1 _05116_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06096_ _10342_/Q _06093_/X _10170_/Q _06094_/X _05985_/X vssd1 vssd1 vccd1 vccd1
+ _10170_/D sky130_fd_sc_hd__a221o_1
XFILLER_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05047_ _05094_/A vssd1 vssd1 vccd1 vccd1 _05047_/X sky130_fd_sc_hd__clkbuf_4
X_09924_ _07453_/Y _07457_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__mux2_2
X_09855_ _10372_/Q _09854_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09855_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08806_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09786_ _08210_/Y _10355_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06998_ _09888_/X vssd1 vssd1 vccd1 vccd1 _07116_/B sky130_fd_sc_hd__clkbuf_2
X_08737_ _08741_/A _08741_/C vssd1 vssd1 vccd1 vccd1 _08737_/X sky130_fd_sc_hd__or2b_1
X_05949_ _06119_/A vssd1 vssd1 vccd1 vccd1 _06111_/A sky130_fd_sc_hd__buf_2
X_08668_ _10067_/Q vssd1 vssd1 vccd1 vccd1 _08668_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07619_ _07619_/A vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__inv_2
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08599_ _08599_/A _08599_/B vssd1 vssd1 vccd1 vccd1 _08599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_198_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10249_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07970_ _07820_/C _07968_/X _07770_/X _07969_/X vssd1 vssd1 vccd1 vccd1 _07971_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06921_ _06909_/A _06909_/B _06945_/A vssd1 vssd1 vccd1 vccd1 _06924_/A sky130_fd_sc_hd__a21o_1
X_09640_ _06374_/X _06376_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__mux2_2
X_06852_ _07155_/A vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__clkbuf_2
X_06783_ _10406_/Q _06814_/B _10407_/Q _06815_/B _06782_/X vssd1 vssd1 vccd1 vccd1
+ _06783_/X sky130_fd_sc_hd__a221o_1
X_09571_ _08398_/Y _09570_/X _09583_/S vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05803_ _05800_/A _10256_/Q _05801_/A _05802_/Y vssd1 vssd1 vccd1 vccd1 _05803_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08522_ _08255_/A _08516_/A _08521_/X _08514_/A _08517_/X vssd1 vssd1 vccd1 vccd1
+ _08596_/C sky130_fd_sc_hd__o2111ai_4
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05734_ _10269_/Q vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__buf_2
X_08453_ _09604_/X _08453_/B vssd1 vssd1 vccd1 vccd1 _08453_/Y sky130_fd_sc_hd__nor2_1
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05665_ _05653_/X _05662_/Y _05663_/Y _08066_/A _05644_/X vssd1 vssd1 vccd1 vccd1
+ _05666_/B sky130_fd_sc_hd__o32a_1
X_07404_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__or2_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ _09509_/X _08391_/B vssd1 vssd1 vccd1 vccd1 _08384_/Y sky130_fd_sc_hd__nor2_1
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05596_ _09987_/X _05566_/X _05667_/A vssd1 vssd1 vccd1 vccd1 _05663_/B sky130_fd_sc_hd__o21ai_1
XFILLER_176_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07335_ _06924_/A _06924_/B _06945_/B vssd1 vssd1 vccd1 vccd1 _07335_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07266_ _07206_/B _07265_/Y _07206_/B _07265_/Y vssd1 vssd1 vccd1 vccd1 _07266_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06217_ _06224_/A vssd1 vssd1 vccd1 vccd1 _06217_/X sky130_fd_sc_hd__clkbuf_2
X_09005_ _08997_/X _09004_/X _08997_/X _09004_/X vssd1 vssd1 vccd1 vccd1 _09005_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07197_ _07197_/A _07197_/B vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__or2_1
XFILLER_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06148_ _06156_/A vssd1 vssd1 vccd1 vccd1 _06148_/X sky130_fd_sc_hd__buf_1
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06079_ _10176_/Q vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__buf_2
XFILLER_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _09443_/X _09441_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09907_/X sky130_fd_sc_hd__mux2_2
XFILLER_116_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09838_ _08268_/X _10368_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09838_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _09768_/X input44/X _09781_/S vssd1 vssd1 vccd1 vccd1 _09769_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05450_ _05445_/B _05439_/X _05449_/Y _05386_/A _05424_/A vssd1 vssd1 vccd1 vccd1
+ _05451_/A sky130_fd_sc_hd__o32a_1
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05381_ _10321_/Q vssd1 vssd1 vccd1 vccd1 _05388_/A sky130_fd_sc_hd__inv_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _07146_/A _07102_/B _07161_/A _07189_/A vssd1 vssd1 vccd1 vccd1 _07121_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_173_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ _07046_/X _07048_/Y _07049_/X _07050_/Y vssd1 vssd1 vccd1 vccd1 _07052_/B
+ sky130_fd_sc_hd__o22a_1
X_06002_ _06031_/A vssd1 vssd1 vccd1 vccd1 _06002_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07953_ _07948_/X _07952_/X _07948_/X _07952_/X vssd1 vssd1 vccd1 vccd1 _07953_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07884_ _07897_/A _07868_/B _07802_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07886_/A
+ sky130_fd_sc_hd__o22a_1
X_06904_ _07118_/A _07031_/B _06904_/C vssd1 vssd1 vccd1 vccd1 _06904_/X sky130_fd_sc_hd__or3_4
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09623_ _09622_/X _09452_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06835_ _06835_/A _06835_/B vssd1 vssd1 vccd1 vccd1 _06836_/B sky130_fd_sc_hd__or2_1
XFILLER_209_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06766_ _10392_/Q _06798_/B _10391_/Q _06795_/B _06765_/X vssd1 vssd1 vccd1 vccd1
+ _06766_/X sky130_fd_sc_hd__o221a_1
X_09554_ _08365_/Y _10116_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09554_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08505_ _10068_/Q vssd1 vssd1 vccd1 vccd1 _08505_/Y sky130_fd_sc_hd__inv_2
X_06697_ _10375_/Q _08711_/A _06695_/Y vssd1 vssd1 vccd1 vccd1 _06815_/B sky130_fd_sc_hd__a21oi_2
X_09485_ _09442_/X _09484_/Y _09442_/X _09484_/Y vssd1 vssd1 vccd1 vccd1 _09485_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05717_ _10292_/Q _05715_/X _05790_/A _05705_/X _05711_/X vssd1 vssd1 vccd1 vccd1
+ _10292_/D sky130_fd_sc_hd__o221a_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08436_ _08436_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_168_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05648_ _05648_/A vssd1 vssd1 vccd1 vccd1 _05648_/Y sky130_fd_sc_hd__inv_2
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08367_ _09008_/A vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05579_ _05579_/A _05516_/X vssd1 vssd1 vccd1 vccd1 _05695_/A sky130_fd_sc_hd__or2b_2
X_07318_ _07052_/A _07052_/B _07052_/Y vssd1 vssd1 vccd1 vccd1 _07318_/X sky130_fd_sc_hd__a21o_1
X_08298_ _08299_/A _08291_/Y _06271_/B vssd1 vssd1 vccd1 vccd1 _08298_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07249_ _07226_/X _07228_/Y _07229_/X _07248_/X _07210_/Y vssd1 vssd1 vccd1 vccd1
+ _07249_/X sky130_fd_sc_hd__o221a_1
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _10300_/CLK _10260_/D vssd1 vssd1 vccd1 vccd1 _10260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10191_ _10436_/CLK _10191_/D vssd1 vssd1 vccd1 vccd1 _10191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 io_wb_dat_i[26] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 io_wb_dat_i[16] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_4
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 io_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 io_wb_dat_i[7] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_6
XFILLER_184_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10421_/CLK _10389_/D vssd1 vssd1 vccd1 vccd1 _10389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06620_ _06620_/A vssd1 vssd1 vccd1 vccd1 _09717_/S sky130_fd_sc_hd__buf_2
XFILLER_203_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06551_ _08427_/A _06540_/X _08430_/A _06540_/X vssd1 vssd1 vccd1 vccd1 _06551_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09270_ _09244_/Y _09269_/X _09244_/Y _09269_/X vssd1 vssd1 vccd1 vccd1 _09270_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06482_ _06482_/A _06482_/B vssd1 vssd1 vccd1 vccd1 _06495_/C sky130_fd_sc_hd__or2_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05502_ _10267_/Q vssd1 vssd1 vccd1 vccd1 _05505_/A sky130_fd_sc_hd__inv_2
XFILLER_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08221_ _08801_/A _08216_/Y _08219_/X _08224_/B vssd1 vssd1 vccd1 vccd1 _08221_/X
+ sky130_fd_sc_hd__o211a_1
X_05433_ _05428_/B _05416_/X _05432_/Y _05390_/A _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05434_/A sky130_fd_sc_hd__o32a_1
XFILLER_193_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08152_ _10353_/Q _08569_/A _08146_/Y _10177_/Q _08151_/X vssd1 vssd1 vccd1 vccd1
+ _08175_/A sky130_fd_sc_hd__o221a_1
X_05364_ _05322_/X _05298_/A _05363_/X vssd1 vssd1 vccd1 vccd1 _10333_/D sky130_fd_sc_hd__o21ai_1
X_08083_ _06634_/Y _06260_/A _10370_/Q _08079_/X _08082_/X vssd1 vssd1 vccd1 vccd1
+ _08083_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05295_ _10331_/Q vssd1 vssd1 vccd1 vccd1 _05296_/B sky130_fd_sc_hd__inv_2
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07103_ _07150_/A _09887_/X vssd1 vssd1 vccd1 vccd1 _07103_/X sky130_fd_sc_hd__or2_1
XFILLER_161_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07034_ _07054_/A _07118_/B vssd1 vssd1 vccd1 vccd1 _07074_/A sky130_fd_sc_hd__or2_1
XFILLER_161_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _08985_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__or2_1
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07936_ _07894_/A _07894_/B _07894_/X vssd1 vssd1 vccd1 vccd1 _07936_/X sky130_fd_sc_hd__a21bo_1
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07867_ _07897_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07867_/X sky130_fd_sc_hd__or2_1
X_06818_ _06818_/A _06818_/B vssd1 vssd1 vccd1 vccd1 _06818_/Y sky130_fd_sc_hd__nor2_1
X_09606_ _10419_/Q _08069_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07798_ _07837_/B vssd1 vssd1 vccd1 vccd1 _07867_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _08760_/A _06666_/B _06667_/B vssd1 vssd1 vccd1 vccd1 _06790_/B sky130_fd_sc_hd__a21bo_1
X_09537_ _09536_/X _10111_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _09468_/A _09906_/X vssd1 vssd1 vccd1 vccd1 _09468_/Y sky130_fd_sc_hd__nor2_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08419_ _09527_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08419_/Y sky130_fd_sc_hd__nor2_1
X_09399_ _09447_/A _09451_/B _09457_/C _09906_/X vssd1 vssd1 vccd1 vccd1 _09399_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10312_ _10312_/CLK _10312_/D vssd1 vssd1 vccd1 vccd1 _10312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10243_ _10249_/CLK _10243_/D vssd1 vssd1 vccd1 vccd1 _10243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _10334_/CLK _10174_/D vssd1 vssd1 vccd1 vccd1 _10174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05080_ _10423_/Q _05094_/A input22/X _05095_/A _05078_/X vssd1 vssd1 vccd1 vccd1
+ _10423_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08770_ _08770_/A vssd1 vssd1 vccd1 vccd1 _08770_/Y sky130_fd_sc_hd__inv_2
X_05982_ _10211_/Q vssd1 vssd1 vccd1 vccd1 _07820_/A sky130_fd_sc_hd__clkbuf_2
X_07721_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07722_/B sky130_fd_sc_hd__nor2_1
X_07652_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _07652_/X sky130_fd_sc_hd__or2_1
X_06603_ _08626_/A vssd1 vssd1 vccd1 vccd1 _06603_/X sky130_fd_sc_hd__buf_2
X_07583_ _07613_/B _09920_/X _07587_/D _09921_/X vssd1 vssd1 vccd1 vccd1 _07585_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09322_ _09321_/A _09321_/B _09321_/Y vssd1 vssd1 vccd1 vccd1 _09322_/Y sky130_fd_sc_hd__o21ai_1
X_06534_ _06539_/B _06533_/Y _06539_/B _06533_/Y vssd1 vssd1 vccd1 vccd1 _06534_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06465_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06466_/A sky130_fd_sc_hd__clkbuf_2
X_09253_ _05933_/X _09251_/X _09252_/X vssd1 vssd1 vccd1 vccd1 _09253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08204_ _08204_/A _08204_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__or2_4
X_09184_ _09083_/A _09085_/Y _09139_/Y _09183_/X vssd1 vssd1 vccd1 vccd1 _09185_/B
+ sky130_fd_sc_hd__a31oi_2
X_06396_ _10141_/Q vssd1 vssd1 vccd1 vccd1 _08409_/A sky130_fd_sc_hd__inv_2
X_05416_ _05439_/A vssd1 vssd1 vccd1 vccd1 _05416_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _06629_/Y _06020_/X _06623_/A _08179_/A vssd1 vssd1 vccd1 vccd1 _08135_/X
+ sky130_fd_sc_hd__o22a_1
X_05347_ _05347_/A vssd1 vssd1 vccd1 vccd1 _05348_/B sky130_fd_sc_hd__inv_2
XFILLER_174_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05278_ _10175_/Q vssd1 vssd1 vccd1 vccd1 _06086_/A sky130_fd_sc_hd__inv_2
X_08066_ _08066_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07017_ _06997_/X _07012_/X _07013_/X _07016_/X vssd1 vssd1 vccd1 vccd1 _07017_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08968_ _08939_/C _08918_/Y _10227_/Q _09142_/A vssd1 vssd1 vccd1 vccd1 _08968_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08899_ _10227_/Q _08978_/A _08899_/C vssd1 vssd1 vccd1 vccd1 _08899_/X sky130_fd_sc_hd__and3_1
X_07919_ _07919_/A vssd1 vssd1 vccd1 vccd1 _07919_/X sky130_fd_sc_hd__buf_1
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10226_ _10289_/CLK _10226_/D vssd1 vssd1 vccd1 vccd1 _10226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10157_ _10330_/CLK _10157_/D vssd1 vssd1 vccd1 vccd1 _10157_/Q sky130_fd_sc_hd__dfxtp_1
X_10088_ _10334_/CLK _10088_/D vssd1 vssd1 vccd1 vccd1 _10088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06250_ _10184_/Q _08206_/A vssd1 vssd1 vccd1 vccd1 _06251_/B sky130_fd_sc_hd__or2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05201_ _05193_/X _10385_/Q _05194_/X _09753_/X _05198_/X vssd1 vssd1 vccd1 vccd1
+ _10385_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06181_ _06181_/A _09662_/X vssd1 vssd1 vccd1 vccd1 _10112_/D sky130_fd_sc_hd__and2_1
XFILLER_209_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05132_ _05129_/X _06615_/A _05131_/Y _05113_/X vssd1 vssd1 vccd1 vccd1 _05133_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05063_ _10434_/Q _05055_/X input34/X _05057_/X _05062_/X vssd1 vssd1 vccd1 vccd1
+ _10434_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _10042_/Q input50/X _09940_/S vssd1 vssd1 vccd1 vccd1 _09940_/X sky130_fd_sc_hd__mux2_1
X_09871_ _10376_/Q _09870_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09871_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08822_ _08822_/A _08822_/B _08806_/A vssd1 vssd1 vccd1 vccd1 _08823_/B sky130_fd_sc_hd__or3b_1
XINSDIODE2_17 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08753_/Y sky130_fd_sc_hd__nor2_1
X_05965_ _05038_/X _05947_/X _05964_/X _05948_/X _05274_/X vssd1 vssd1 vccd1 vccd1
+ _10218_/D sky130_fd_sc_hd__a221o_1
X_07704_ _07654_/X _07702_/X _07654_/X _07702_/X vssd1 vssd1 vccd1 vccd1 _07704_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08684_ _08674_/C _08683_/X _08679_/X vssd1 vssd1 vccd1 vccd1 _08684_/X sky130_fd_sc_hd__o21a_1
X_05896_ _05910_/A vssd1 vssd1 vccd1 vccd1 _05896_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07635_ _07814_/A vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _10213_/Q _07566_/B _07577_/A vssd1 vssd1 vccd1 vccd1 _07567_/A sky130_fd_sc_hd__and3_1
X_06517_ _08411_/A _06536_/A _08415_/A _06496_/X _06507_/X vssd1 vssd1 vccd1 vccd1
+ _06517_/X sky130_fd_sc_hd__o221a_1
X_09305_ _09392_/A _09304_/B _09304_/Y vssd1 vssd1 vccd1 vccd1 _09305_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _09174_/A _09229_/B _09122_/A _09173_/X _09174_/X vssd1 vssd1 vccd1 vccd1
+ _09297_/A sky130_fd_sc_hd__o32a_1
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07497_ _07868_/A vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06448_ _06447_/A _06447_/B _06447_/X vssd1 vssd1 vccd1 vccd1 _06448_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09166_/A _09166_/B _09222_/A vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__a21o_1
X_06379_ _06377_/Y _10139_/Q _10246_/Q _08401_/A vssd1 vssd1 vccd1 vccd1 _06384_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08118_ _08632_/A _10180_/Q _06633_/Y _06262_/A _08117_/X vssd1 vssd1 vccd1 vccd1
+ _08119_/D sky130_fd_sc_hd__o221a_1
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09098_ _09095_/Y _09097_/X _09095_/Y _09097_/X vssd1 vssd1 vccd1 vccd1 _09098_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08049_ _07403_/A _07403_/B _07404_/B vssd1 vssd1 vccd1 vccd1 _08049_/X sky130_fd_sc_hd__a21bo_1
XFILLER_122_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10011_ _08003_/A _08032_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10011_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10209_ _10414_/CLK _10209_/D vssd1 vssd1 vccd1 vccd1 _10209_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05750_ _05750_/A vssd1 vssd1 vccd1 vccd1 _05871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05681_ _10302_/Q vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__inv_2
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ _08855_/B _07418_/B _07419_/Y vssd1 vssd1 vccd1 vccd1 _07420_/X sky130_fd_sc_hd__a21o_1
XFILLER_210_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07351_ _07280_/X _07299_/Y _07280_/X _07299_/Y vssd1 vssd1 vccd1 vccd1 _07351_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06302_ _10237_/Q _08349_/A _06294_/B _06297_/X vssd1 vssd1 vccd1 vccd1 _06302_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ _07185_/X _07200_/X _07185_/X _07200_/X vssd1 vssd1 vccd1 vccd1 _07283_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_06233_ _10036_/D vssd1 vssd1 vccd1 vccd1 _06233_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09021_ _08864_/X _09020_/X _08864_/X _09020_/X vssd1 vssd1 vccd1 vccd1 _09022_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06164_ _06176_/A vssd1 vssd1 vccd1 vccd1 _06169_/A sky130_fd_sc_hd__buf_1
X_05115_ _05133_/A _05115_/B vssd1 vssd1 vccd1 vccd1 _10410_/D sky130_fd_sc_hd__nor2_1
XFILLER_144_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06095_ _10343_/Q _06093_/X _10171_/Q _06094_/X _05985_/X vssd1 vssd1 vccd1 vccd1
+ _10171_/D sky130_fd_sc_hd__a221o_1
XFILLER_131_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09923_ _09219_/X _09217_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09923_/X sky130_fd_sc_hd__mux2_2
X_05046_ _05072_/A vssd1 vssd1 vccd1 vccd1 _05094_/A sky130_fd_sc_hd__clkbuf_2
X_09854_ _08284_/X _10372_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09854_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08805_ _08822_/A _08803_/X _08821_/C vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__o21bai_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _09784_/X input48/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06997_ _06980_/X _06996_/X _06980_/X _06996_/X vssd1 vssd1 vccd1 vccd1 _06997_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08736_ _08733_/A _08733_/B _08255_/A _08735_/X vssd1 vssd1 vccd1 vccd1 _08741_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_05948_ _05948_/A vssd1 vssd1 vccd1 vccd1 _05948_/X sky130_fd_sc_hd__clkbuf_2
X_08667_ _08121_/X _10052_/Q _08655_/X _08663_/Y _08705_/A vssd1 vssd1 vccd1 vccd1
+ _08667_/Y sky130_fd_sc_hd__a221oi_2
X_05879_ _05816_/X _05878_/X _05816_/X _05878_/X vssd1 vssd1 vccd1 vccd1 _06821_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_202_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07618_ _07598_/X _07599_/X _07598_/X _07599_/X vssd1 vssd1 vccd1 vccd1 _07619_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08598_ _08598_/A vssd1 vssd1 vccd1 vccd1 _08598_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07549_ _07819_/A _09934_/X _07815_/A _09936_/X _07548_/Y vssd1 vssd1 vccd1 vccd1
+ _07550_/B sky130_fd_sc_hd__o41a_1
XFILLER_194_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09219_ _09218_/A _09218_/B _09276_/A vssd1 vssd1 vccd1 vccd1 _09219_/X sky130_fd_sc_hd__a21bo_1
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06920_ _06920_/A vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__inv_2
X_06851_ _10219_/Q vssd1 vssd1 vccd1 vccd1 _07155_/A sky130_fd_sc_hd__inv_2
X_06782_ _10405_/Q _06813_/B _10406_/Q _06814_/B _06781_/X vssd1 vssd1 vccd1 vccd1
+ _06782_/X sky130_fd_sc_hd__o221a_1
X_09570_ _08399_/Y _10122_/Q _09582_/S vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__mux2_1
X_05802_ _10256_/Q vssd1 vssd1 vccd1 vccd1 _05802_/Y sky130_fd_sc_hd__inv_2
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08521_/X sky130_fd_sc_hd__or2_2
X_05733_ _10286_/Q _05728_/X _08855_/B _05732_/X _05724_/X vssd1 vssd1 vccd1 vccd1
+ _10286_/D sky130_fd_sc_hd__o221a_1
X_08452_ _08452_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08452_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05664_ _10305_/Q vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__inv_2
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ _07403_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__or2_1
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05595_ _05668_/A _05668_/B vssd1 vssd1 vccd1 vccd1 _05667_/A sky130_fd_sc_hd__nand2_1
X_08383_ _08383_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__or2_1
XFILLER_149_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07334_ _07330_/X _07331_/X _07330_/X _07331_/X vssd1 vssd1 vccd1 vccd1 _07334_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07265_ _07129_/X _07202_/Y _07206_/A vssd1 vssd1 vccd1 vccd1 _07265_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_191_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06216_ _09690_/X _06210_/X _10091_/Q _06211_/X vssd1 vssd1 vccd1 vccd1 _10091_/D
+ sky130_fd_sc_hd__a22o_1
X_09004_ _09074_/C _09003_/B _09036_/A vssd1 vssd1 vccd1 vccd1 _09004_/X sky130_fd_sc_hd__a21bo_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ _07178_/B _07180_/B _07178_/B _07195_/X vssd1 vssd1 vccd1 vccd1 _07197_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06147_ _09656_/X _06140_/X _10138_/Q _06141_/X _06146_/X vssd1 vssd1 vccd1 vccd1
+ _10138_/D sky130_fd_sc_hd__o221a_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06078_ _09761_/X _06028_/A _10177_/Q _06031_/A _06032_/A vssd1 vssd1 vccd1 vccd1
+ _10177_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09906_ _09388_/X _09387_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__mux2_2
X_05029_ _10447_/Q _09940_/S _05028_/X _05013_/X _06182_/A vssd1 vssd1 vccd1 vccd1
+ _10447_/D sky130_fd_sc_hd__o221a_1
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09837_ _09836_/X input31/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09768_ _09767_/X _08194_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08719_ _08719_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09699_ _06548_/X input32/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__mux2_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05380_ _10322_/Q vssd1 vssd1 vccd1 vccd1 _05389_/A sky130_fd_sc_hd__inv_2
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07050_ _07050_/A _07050_/B vssd1 vssd1 vccd1 vccd1 _07050_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06001_ _06069_/A vssd1 vssd1 vccd1 vccd1 _06031_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ _07922_/Y _07949_/X _07950_/X _07951_/X vssd1 vssd1 vccd1 vccd1 _07952_/X
+ sky130_fd_sc_hd__o22a_1
X_07883_ _07880_/X _07882_/X _07880_/X _07882_/X vssd1 vssd1 vccd1 vccd1 _07883_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06903_ _06903_/A vssd1 vssd1 vccd1 vccd1 _06904_/C sky130_fd_sc_hd__inv_2
XFILLER_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09622_ _08370_/X _06320_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09622_/X sky130_fd_sc_hd__mux2_1
X_06834_ _06834_/A _06834_/B vssd1 vssd1 vccd1 vccd1 _06835_/B sky130_fd_sc_hd__or2_1
X_09553_ _09552_/X _10352_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09553_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__or2_1
X_06765_ _10391_/Q _06795_/B _06764_/X vssd1 vssd1 vccd1 vccd1 _06765_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ _06626_/Y _06695_/Y _08707_/A vssd1 vssd1 vccd1 vccd1 _06698_/A sky130_fd_sc_hd__o21ai_2
X_09484_ _09478_/X _09483_/X _09478_/X _09483_/X vssd1 vssd1 vccd1 vccd1 _09484_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_102_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05716_ _10276_/Q vssd1 vssd1 vccd1 vccd1 _05790_/A sky130_fd_sc_hd__buf_2
XFILLER_211_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08435_ _09961_/X _08435_/B vssd1 vssd1 vccd1 vccd1 _08435_/X sky130_fd_sc_hd__and2_1
X_05647_ _05678_/A vssd1 vssd1 vccd1 vccd1 _05677_/A sky130_fd_sc_hd__clkbuf_2
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08366_ _10232_/Q vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__inv_2
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05578_ _06887_/A _07234_/B _07660_/A _07814_/A vssd1 vssd1 vccd1 vccd1 _05579_/A
+ sky130_fd_sc_hd__o22a_1
X_07317_ _06953_/X _06958_/X _06953_/X _06958_/X vssd1 vssd1 vccd1 vccd1 _07317_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08297_ _08297_/A vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07248_ _07242_/A _07269_/A _07241_/Y _07239_/A _07247_/Y vssd1 vssd1 vccd1 vccd1
+ _07248_/X sky130_fd_sc_hd__o32a_1
XFILLER_191_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07179_ _07167_/X _07168_/X _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07180_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _10426_/CLK _10190_/D vssd1 vssd1 vccd1 vccd1 _10190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_30_clock clkbuf_2_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10447_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput27 io_wb_dat_i[17] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_4
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 io_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
Xinput38 io_wb_dat_i[27] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput49 io_wb_dat_i[8] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10388_ _10422_/CLK _10388_/D vssd1 vssd1 vccd1 vccd1 _10388_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06550_ _10101_/Q _06464_/A _08432_/A _06540_/A vssd1 vssd1 vccd1 vccd1 _06560_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06481_ _08392_/A _06432_/A _10089_/Q _06462_/A vssd1 vssd1 vccd1 vccd1 _06495_/A
+ sky130_fd_sc_hd__a22o_1
X_05501_ _07150_/A vssd1 vssd1 vccd1 vccd1 _06887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__or2_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05432_ _10323_/Q _05432_/B vssd1 vssd1 vccd1 vccd1 _05432_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08151_ _10362_/Q _08533_/A _06633_/A _08265_/A vssd1 vssd1 vccd1 vccd1 _08151_/X
+ sky130_fd_sc_hd__o22a_1
X_05363_ _10333_/Q _05362_/Y _05298_/A _05362_/A _05282_/X vssd1 vssd1 vccd1 vccd1
+ _05363_/X sky130_fd_sc_hd__a221o_1
X_08082_ _06714_/Y _08733_/A _08762_/A _08081_/X vssd1 vssd1 vccd1 vccd1 _08082_/X
+ sky130_fd_sc_hd__a22o_1
X_05294_ _10332_/Q vssd1 vssd1 vccd1 vccd1 _05296_/A sky130_fd_sc_hd__inv_2
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07102_ _07125_/A _07102_/B _07161_/A _09890_/X vssd1 vssd1 vccd1 vccd1 _07102_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07033_ _09887_/X vssd1 vssd1 vccd1 vccd1 _07118_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08984_ _08984_/A vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__inv_2
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07935_ _07912_/X _07913_/Y _07912_/X _07913_/Y vssd1 vssd1 vccd1 vccd1 _07935_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09605_ _10418_/Q _08068_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09605_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07866_ _07483_/A _07800_/X _07885_/A _07864_/Y _07865_/X vssd1 vssd1 vccd1 vccd1
+ _07869_/A sky130_fd_sc_hd__a41o_1
X_06817_ _06818_/A _06817_/B vssd1 vssd1 vccd1 vccd1 _06817_/Y sky130_fd_sc_hd__nor2_1
X_07797_ _09916_/X vssd1 vssd1 vccd1 vccd1 _07837_/B sky130_fd_sc_hd__buf_1
X_06748_ _10386_/Q vssd1 vssd1 vccd1 vccd1 _06748_/Y sky130_fd_sc_hd__inv_2
X_09536_ _10079_/Q _10041_/Q _09544_/S vssd1 vssd1 vccd1 vccd1 _09536_/X sky130_fd_sc_hd__mux2_1
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09462_/X _09466_/X _09462_/X _09466_/X vssd1 vssd1 vccd1 vccd1 _09467_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06679_ _10367_/Q _08729_/A vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__or2_2
X_08418_ _08418_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08418_/Y sky130_fd_sc_hd__nor2_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09398_ _09906_/X vssd1 vssd1 vccd1 vccd1 _09398_/Y sky130_fd_sc_hd__inv_2
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ _08349_/A _09748_/S vssd1 vssd1 vccd1 vccd1 _08349_/X sky130_fd_sc_hd__or2_1
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10426_/CLK _10311_/D vssd1 vssd1 vccd1 vccd1 _10311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10242_ _10249_/CLK _10242_/D vssd1 vssd1 vccd1 vccd1 _10242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _10334_/CLK _10173_/D vssd1 vssd1 vccd1 vccd1 _10173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05981_ _10212_/Q _05970_/A input41/X _05971_/A _05978_/X vssd1 vssd1 vccd1 vccd1
+ _10212_/D sky130_fd_sc_hd__o221a_1
X_07720_ _07694_/A _07700_/A _07694_/Y vssd1 vssd1 vccd1 vccd1 _07720_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07651_ _07573_/A _07579_/A _07573_/Y vssd1 vssd1 vccd1 vccd1 _07652_/B sky130_fd_sc_hd__a21o_1
X_06602_ _08461_/A vssd1 vssd1 vccd1 vccd1 _08626_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _07578_/A _07578_/B _07648_/B vssd1 vssd1 vccd1 vccd1 _07582_/X sky130_fd_sc_hd__a21o_1
X_09321_ _09321_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09321_/Y sky130_fd_sc_hd__nand2_1
X_06533_ _08423_/A _06489_/X _06539_/A _06529_/X vssd1 vssd1 vccd1 vccd1 _06533_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06464_ _06464_/A vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__clkbuf_2
X_09252_ _09252_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__or2_1
XFILLER_193_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _08569_/A _08198_/Y _06249_/B vssd1 vssd1 vccd1 vccd1 _08203_/Y sky130_fd_sc_hd__o21ai_1
X_09183_ _09083_/B _09137_/Y _09136_/Y vssd1 vssd1 vccd1 vccd1 _09183_/X sky130_fd_sc_hd__o21a_1
X_06395_ _06391_/X _06394_/X _06391_/X _06394_/X vssd1 vssd1 vccd1 vccd1 _06395_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_05415_ _05415_/A vssd1 vssd1 vccd1 vccd1 _10327_/D sky130_fd_sc_hd__inv_2
X_08134_ _08289_/A vssd1 vssd1 vccd1 vccd1 _08134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05346_ _05346_/A vssd1 vssd1 vccd1 vccd1 _10338_/D sky130_fd_sc_hd__inv_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05277_ _05038_/X _05215_/X _06621_/A _05216_/X _05274_/X vssd1 vssd1 vccd1 vccd1
+ _10347_/D sky130_fd_sc_hd__a221o_1
XFILLER_146_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08065_ _08065_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07016_ _07016_/A vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08967_ _08912_/X _08966_/X _08912_/X _08966_/X vssd1 vssd1 vccd1 vccd1 _08967_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08898_ _08915_/A _09985_/X vssd1 vssd1 vccd1 vccd1 _08939_/C sky130_fd_sc_hd__nor2_4
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07918_ _07915_/X _07917_/X _07915_/X _07917_/X vssd1 vssd1 vccd1 vccd1 _07918_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07849_ _07849_/A _07849_/B vssd1 vssd1 vccd1 vccd1 _07850_/B sky130_fd_sc_hd__or2_2
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _09518_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10225_ _10225_/CLK _10225_/D vssd1 vssd1 vccd1 vccd1 _10225_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _10328_/CLK _10156_/D vssd1 vssd1 vccd1 vccd1 _10156_/Q sky130_fd_sc_hd__dfxtp_1
X_10087_ _10334_/CLK _10087_/D vssd1 vssd1 vccd1 vccd1 _10087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05200_ _05193_/X _10386_/Q _05194_/X _09605_/X _05198_/X vssd1 vssd1 vccd1 vccd1
+ _10386_/D sky130_fd_sc_hd__o221a_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06180_ _06181_/A _09663_/X vssd1 vssd1 vccd1 vccd1 _10113_/D sky130_fd_sc_hd__and2_1
XFILLER_209_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05131_ _10438_/Q vssd1 vssd1 vccd1 vccd1 _05131_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05062_ _05189_/A vssd1 vssd1 vccd1 vccd1 _05062_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _08302_/X _10376_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08821_ _08821_/A _08821_/B _08821_/C _08765_/X vssd1 vssd1 vccd1 vccd1 _08822_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_18 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ _08752_/A _08752_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__or2_2
XFILLER_85_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05964_ _10218_/Q vssd1 vssd1 vccd1 vccd1 _05964_/X sky130_fd_sc_hd__clkbuf_2
X_08683_ _06038_/X _08676_/Y _06035_/X _08524_/Y _08682_/Y vssd1 vssd1 vccd1 vccd1
+ _08683_/X sky130_fd_sc_hd__o221a_1
X_07703_ _07528_/A _07528_/B _07706_/B vssd1 vssd1 vccd1 vccd1 _07703_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05895_ _05911_/A vssd1 vssd1 vccd1 vccd1 _05910_/A sky130_fd_sc_hd__inv_2
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07634_ _07634_/A vssd1 vssd1 vccd1 vccd1 _07634_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07565_ _07837_/A _07634_/A vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__or2_1
XFILLER_139_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06516_ _06516_/A _06516_/B _06516_/C _06516_/D vssd1 vssd1 vccd1 vccd1 _06516_/X
+ sky130_fd_sc_hd__or4_4
X_09304_ _09392_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _09304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07496_ _07496_/A _07496_/B vssd1 vssd1 vccd1 vccd1 _07496_/X sky130_fd_sc_hd__or2_1
X_06447_ _06447_/A _06447_/B vssd1 vssd1 vccd1 vccd1 _06447_/X sky130_fd_sc_hd__or2_2
X_09235_ _05939_/X _09232_/Y _09233_/X _09234_/Y vssd1 vssd1 vccd1 vccd1 _09235_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09166_ _09166_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__nor2_2
X_06378_ _10139_/Q vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__inv_2
X_08117_ _06634_/Y _06260_/A _08624_/B _08116_/X vssd1 vssd1 vccd1 vccd1 _08117_/X
+ sky130_fd_sc_hd__o22a_1
X_09097_ _09097_/A _09245_/B _09009_/X vssd1 vssd1 vccd1 vccd1 _09097_/X sky130_fd_sc_hd__or3b_1
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05329_ _05329_/A vssd1 vssd1 vccd1 vccd1 _05330_/B sky130_fd_sc_hd__inv_2
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ _08018_/A _08018_/B _08019_/B vssd1 vssd1 vccd1 vccd1 _08048_/X sky130_fd_sc_hd__a21bo_1
X_10010_ _08004_/A _08034_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09999_ _09998_/X _07028_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09999_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _10414_/CLK _10208_/D vssd1 vssd1 vccd1 vccd1 _10208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ _10328_/CLK _10139_/D vssd1 vssd1 vccd1 vccd1 _10139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05680_ _05680_/A _05680_/B vssd1 vssd1 vccd1 vccd1 _05680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _06984_/X _07349_/X _06984_/X _07349_/X vssd1 vssd1 vccd1 vccd1 _07350_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06301_ _06299_/Y _10131_/Q _10238_/Q _08355_/A vssd1 vssd1 vccd1 vccd1 _06304_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ _08850_/A _08850_/B _08850_/Y vssd1 vssd1 vccd1 vccd1 _09020_/X sky130_fd_sc_hd__a21o_1
X_07281_ _07246_/A _07246_/B _07268_/B vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__a21o_1
X_06232_ _09678_/X _06203_/A _10079_/Q _06204_/A vssd1 vssd1 vccd1 vccd1 _10079_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06163_ _09645_/X _06156_/A _10127_/Q _06157_/A _05468_/X vssd1 vssd1 vccd1 vccd1
+ _10127_/D sky130_fd_sc_hd__o221a_1
X_05114_ _06614_/A _05193_/A _05109_/Y _05113_/X vssd1 vssd1 vccd1 vccd1 _05115_/B
+ sky130_fd_sc_hd__o22a_1
X_06094_ _06102_/A vssd1 vssd1 vccd1 vccd1 _06094_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05045_ _05073_/A vssd1 vssd1 vccd1 vccd1 _05072_/A sky130_fd_sc_hd__inv_2
X_09922_ _09337_/Y _09336_/B _09994_/S vssd1 vssd1 vccd1 vccd1 _09922_/X sky130_fd_sc_hd__mux2_2
X_09853_ _09852_/X input35/X _09881_/S vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _08821_/C sky130_fd_sc_hd__nor2_1
X_09784_ _09783_/X _08209_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09784_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08735_ _06715_/Y _08636_/Y _10365_/Q _08734_/X vssd1 vssd1 vccd1 vccd1 _08735_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06996_ _06984_/X _06990_/Y _07227_/B _06991_/Y _06995_/X vssd1 vssd1 vccd1 vccd1
+ _06996_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05947_ _05947_/A vssd1 vssd1 vccd1 vccd1 _05947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08666_ _08666_/A _08666_/B _08666_/C _08646_/X vssd1 vssd1 vccd1 vccd1 _08705_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05878_ _07415_/A _10253_/Q _05811_/Y vssd1 vssd1 vccd1 vccd1 _05878_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _08597_/A _08597_/B _08597_/C _08596_/Y vssd1 vssd1 vccd1 vccd1 _08598_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07617_ _07611_/X _07616_/X _07611_/X _07616_/X vssd1 vssd1 vccd1 vccd1 _07640_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07548_ _07552_/C _07548_/B vssd1 vssd1 vccd1 vccd1 _07548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07479_ _07547_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ _09218_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__or2_1
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09149_ _09147_/Y _09193_/B _09147_/Y _09193_/B vssd1 vssd1 vccd1 vccd1 _09150_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06850_ _06834_/A _06834_/B _06835_/B vssd1 vssd1 vccd1 vccd1 _06850_/X sky130_fd_sc_hd__a21bo_1
XFILLER_67_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05801_ _05801_/A vssd1 vssd1 vccd1 vccd1 _05801_/X sky130_fd_sc_hd__clkbuf_2
X_06781_ _10405_/Q _06813_/B _10404_/Q _06812_/B _06780_/X vssd1 vssd1 vccd1 vccd1
+ _06781_/X sky130_fd_sc_hd__a221o_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _08521_/A _08521_/B _08809_/A _08519_/X vssd1 vssd1 vccd1 vccd1 _08520_/Y
+ sky130_fd_sc_hd__a22oi_2
X_05732_ _05761_/A vssd1 vssd1 vccd1 vccd1 _05732_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_208_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ _09963_/X _08453_/B vssd1 vssd1 vccd1 vccd1 _08451_/Y sky130_fd_sc_hd__nor2_1
X_05663_ _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_196_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07402_ _07402_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07403_/B sky130_fd_sc_hd__or2_1
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _08382_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08382_/Y sky130_fd_sc_hd__nor2_1
X_05594_ _09974_/X _05568_/X _05672_/A vssd1 vssd1 vccd1 vccd1 _05668_/B sky130_fd_sc_hd__o21ai_1
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07333_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07333_/X sky130_fd_sc_hd__and2_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07264_ _07260_/X _07261_/X _07260_/X _07261_/X vssd1 vssd1 vccd1 vccd1 _07264_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06215_ _09691_/X _06210_/X _10092_/Q _06211_/X vssd1 vssd1 vccd1 vccd1 _10092_/D
+ sky130_fd_sc_hd__a22o_1
X_09003_ _09074_/C _09003_/B vssd1 vssd1 vccd1 vccd1 _09036_/A sky130_fd_sc_hd__or2_2
X_07195_ _07180_/A _07180_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07195_/X sky130_fd_sc_hd__a21bo_1
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06146_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06146_/X sky130_fd_sc_hd__clkbuf_2
X_06077_ _09765_/X _06067_/X _08657_/A _06069_/X _06070_/X vssd1 vssd1 vccd1 vccd1
+ _10178_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05028_ input45/X vssd1 vssd1 vccd1 vccd1 _05028_/X sky130_fd_sc_hd__clkbuf_4
X_09905_ _07414_/X _07369_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09836_ _09835_/X _08266_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09836_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09767_ _10350_/Q _09766_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__mux2_1
X_06979_ _07235_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _06985_/A sky130_fd_sc_hd__or2_2
XFILLER_39_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08718_ _08715_/A _08717_/B _06629_/Y _08717_/Y vssd1 vssd1 vccd1 vccd1 _08718_/X
+ sky130_fd_sc_hd__o22a_1
X_09698_ _06544_/X input31/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08649_ _08664_/A _08649_/B vssd1 vssd1 vccd1 vccd1 _08649_/X sky130_fd_sc_hd__or2_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06000_ _06000_/A vssd1 vssd1 vccd1 vccd1 _06273_/A sky130_fd_sc_hd__buf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07951_ _07922_/Y _07949_/X _07922_/Y _07949_/X vssd1 vssd1 vccd1 vccd1 _07951_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_141_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06902_ _06962_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__or2_2
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ _07882_/A _07882_/B vssd1 vssd1 vccd1 vccd1 _07882_/X sky130_fd_sc_hd__or2_1
XFILLER_95_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _09620_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__mux2_1
X_06833_ _06826_/A _06826_/B _06827_/B vssd1 vssd1 vccd1 vccd1 _06833_/X sky130_fd_sc_hd__a21bo_1
X_06764_ _10390_/Q _06794_/B _06763_/Y vssd1 vssd1 vccd1 vccd1 _06764_/X sky130_fd_sc_hd__a21bo_1
X_09552_ _10384_/Q _10181_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09552_/X sky130_fd_sc_hd__mux2_1
X_08503_ _10067_/Q _08485_/B _08502_/Y vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05715_ _05741_/A vssd1 vssd1 vccd1 vccd1 _05715_/X sky130_fd_sc_hd__clkbuf_2
X_06695_ _08709_/A vssd1 vssd1 vccd1 vccd1 _06695_/Y sky130_fd_sc_hd__inv_2
X_09483_ _09479_/Y _09482_/Y _09479_/Y _09482_/Y vssd1 vssd1 vccd1 vccd1 _09483_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08434_ _08434_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08434_/Y sky130_fd_sc_hd__nor2_1
X_05646_ _05646_/A _05646_/B vssd1 vssd1 vccd1 vccd1 _10309_/D sky130_fd_sc_hd__nor2_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ _08365_/A _09544_/S vssd1 vssd1 vccd1 vccd1 _08365_/Y sky130_fd_sc_hd__nor2_1
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05577_ _05498_/X _05516_/X _05498_/X _05516_/X vssd1 vssd1 vccd1 vccd1 _05577_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_07316_ _07309_/A _07309_/B _07309_/X vssd1 vssd1 vccd1 vccd1 _07316_/X sky130_fd_sc_hd__a21bo_1
X_08296_ _08294_/A _08294_/B _08193_/X _08295_/Y vssd1 vssd1 vccd1 vccd1 _08296_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_176_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07247_ _07247_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07178_ _07182_/B _07178_/B vssd1 vssd1 vccd1 vccd1 _07178_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06129_ _10148_/Q _06126_/X _10320_/Q _06122_/X _06128_/X vssd1 vssd1 vccd1 vccd1
+ _10148_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09819_ _10363_/Q _09818_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 io_wb_dat_i[18] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 io_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
Xinput39 io_wb_dat_i[28] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10387_ _10422_/CLK _10387_/D vssd1 vssd1 vccd1 vccd1 _10387_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06480_ _10089_/Q vssd1 vssd1 vccd1 vccd1 _08392_/A sky130_fd_sc_hd__inv_2
X_05500_ _07147_/A vssd1 vssd1 vccd1 vccd1 _07150_/A sky130_fd_sc_hd__clkbuf_2
X_05431_ _05431_/A vssd1 vssd1 vccd1 vccd1 _05432_/B sky130_fd_sc_hd__inv_2
X_08150_ _08526_/A vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__buf_2
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05362_ _05362_/A vssd1 vssd1 vccd1 vccd1 _05362_/Y sky130_fd_sc_hd__inv_2
X_07101_ _07165_/A _06999_/Y _07099_/Y _07099_/A _07100_/X vssd1 vssd1 vccd1 vccd1
+ _07101_/X sky130_fd_sc_hd__a32o_1
X_08081_ _08215_/A vssd1 vssd1 vccd1 vccd1 _08081_/X sky130_fd_sc_hd__buf_2
X_05293_ _10333_/Q vssd1 vssd1 vccd1 vccd1 _05298_/A sky130_fd_sc_hd__inv_2
XFILLER_173_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07032_ _07030_/X _07031_/Y _07030_/X _07031_/Y vssd1 vssd1 vccd1 vccd1 _07032_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _08947_/X _08982_/X _08947_/X _08982_/X vssd1 vssd1 vccd1 vccd1 _08984_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07934_ _07930_/X _07933_/X _07930_/X _07933_/X vssd1 vssd1 vccd1 vccd1 _07934_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07865_ _07678_/A _07867_/B _07485_/A _07864_/A vssd1 vssd1 vccd1 vccd1 _07865_/X
+ sky130_fd_sc_hd__o22a_1
X_09604_ _09603_/X _06624_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09604_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06816_ _06818_/A _06816_/B vssd1 vssd1 vccd1 vccd1 _06816_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07796_ _07786_/X _07795_/X _07786_/X _07795_/X vssd1 vssd1 vccd1 vccd1 _07903_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_09535_ _09534_/X _10347_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09535_/X sky130_fd_sc_hd__mux2_1
X_06747_ _06733_/Y _06788_/B _06607_/Y _06736_/X _06746_/X vssd1 vssd1 vccd1 vccd1
+ _06747_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06678_ _10366_/Q _08731_/A vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__or2_2
X_09466_ _09463_/X _09465_/X _09463_/X _09465_/X vssd1 vssd1 vccd1 vccd1 _09466_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_196_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ _08452_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__clkbuf_2
X_05629_ _05619_/X _05626_/Y _05627_/Y _08074_/A _05623_/X vssd1 vssd1 vccd1 vccd1
+ _05630_/B sky130_fd_sc_hd__o32a_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ _09451_/B vssd1 vssd1 vccd1 vccd1 _09397_/Y sky130_fd_sc_hd__inv_2
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _09343_/A vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08279_ _08079_/X _08277_/B _08240_/X _08278_/Y vssd1 vssd1 vccd1 vccd1 _08279_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ _10420_/CLK _10310_/D vssd1 vssd1 vccd1 vccd1 _10310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10241_ _10249_/CLK _10241_/D vssd1 vssd1 vccd1 vccd1 _10241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _10334_/CLK _10172_/D vssd1 vssd1 vccd1 vccd1 _10172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10439_ _10442_/CLK _10439_/D vssd1 vssd1 vccd1 vccd1 _10439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05980_ _10213_/Q _05970_/A input44/X _05971_/A _05978_/X vssd1 vssd1 vccd1 vccd1
+ _10213_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _07650_/A _07650_/B vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__or2_1
X_06601_ _10447_/Q vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__inv_2
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ _07559_/X _07580_/X _07559_/X _07580_/X vssd1 vssd1 vccd1 vccd1 _07581_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09320_ _09320_/A _09430_/A vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__or2_1
X_06532_ _10098_/Q _06464_/A _08425_/A _06434_/A vssd1 vssd1 vccd1 vccd1 _06539_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09251_ _09251_/A vssd1 vssd1 vccd1 vccd1 _09251_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06463_ _06463_/A vssd1 vssd1 vccd1 vccd1 _06464_/A sky130_fd_sc_hd__clkbuf_2
X_08202_ _08155_/X _08200_/B _08201_/Y _08193_/X vssd1 vssd1 vccd1 vccd1 _08202_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09182_ _09181_/A _09181_/B _09181_/X vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__a21bo_1
X_06394_ _10246_/Q _08401_/A _06384_/A _06381_/X vssd1 vssd1 vccd1 vccd1 _06394_/X
+ sky130_fd_sc_hd__o22a_1
X_05414_ _05407_/B _05372_/X _05413_/Y _05394_/A _05409_/X vssd1 vssd1 vccd1 vccd1
+ _05415_/A sky130_fd_sc_hd__o32a_1
X_08133_ _10202_/Q vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__inv_2
X_05345_ _05340_/B _05333_/X _05344_/Y _05336_/X _05302_/A vssd1 vssd1 vccd1 vccd1
+ _05346_/A sky130_fd_sc_hd__o32a_1
XFILLER_146_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08064_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08071_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_161_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05276_ _10347_/Q vssd1 vssd1 vccd1 vccd1 _06621_/A sky130_fd_sc_hd__buf_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07015_ _06970_/A _06993_/B _06991_/Y _07014_/Y vssd1 vssd1 vccd1 vccd1 _07016_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _09294_/A _09142_/A _08993_/C _08965_/X vssd1 vssd1 vccd1 vccd1 _08966_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08897_ _08934_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _08936_/C sky130_fd_sc_hd__or2_2
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07917_ _07921_/B _07916_/C _07767_/X _07778_/X _07916_/X vssd1 vssd1 vccd1 vccd1
+ _07917_/X sky130_fd_sc_hd__o221a_1
XFILLER_84_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07848_ _07824_/C _07821_/B _07821_/Y vssd1 vssd1 vccd1 vccd1 _07849_/B sky130_fd_sc_hd__o21ai_1
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ _08413_/X _06405_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09518_/X sky130_fd_sc_hd__mux2_1
X_07779_ _07767_/X _07778_/X _07767_/X _07778_/X vssd1 vssd1 vccd1 vccd1 _07779_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09447_/Y _09448_/X _09447_/Y _09448_/X vssd1 vssd1 vccd1 vccd1 _09449_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10224_ _10225_/CLK _10224_/D vssd1 vssd1 vccd1 vccd1 _10224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10155_ _10328_/CLK _10155_/D vssd1 vssd1 vccd1 vccd1 _10155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10086_ _10334_/CLK _10086_/D vssd1 vssd1 vccd1 vccd1 _10086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05130_ _10406_/Q vssd1 vssd1 vccd1 vccd1 _06615_/A sky130_fd_sc_hd__inv_2
XFILLER_128_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05061_ _10435_/Q _05055_/X input35/X _05057_/X _05053_/X vssd1 vssd1 vccd1 vccd1
+ _10435_/D sky130_fd_sc_hd__o221a_1
XFILLER_171_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ _08820_/A _08820_/B _08820_/C _08801_/X vssd1 vssd1 vccd1 vccd1 _08821_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_97_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_19 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__or2_1
X_05963_ _07108_/A _05947_/A _05101_/X _05948_/A _05960_/X vssd1 vssd1 vccd1 vccd1
+ _10219_/D sky130_fd_sc_hd__o221a_1
XFILLER_57_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08682_ _08674_/B _08673_/X _08677_/X vssd1 vssd1 vccd1 vccd1 _08682_/Y sky130_fd_sc_hd__o21ai_1
X_05894_ _06083_/A _08315_/A vssd1 vssd1 vccd1 vccd1 _05911_/A sky130_fd_sc_hd__or2_2
X_07702_ _07675_/X _07680_/X _07681_/X _07701_/X _07658_/Y vssd1 vssd1 vccd1 vccd1
+ _07702_/X sky130_fd_sc_hd__o221a_1
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07633_ _07631_/X _07632_/X _07631_/X _07632_/X vssd1 vssd1 vccd1 vccd1 _07633_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07564_ _07550_/X _07552_/X _07550_/X _07552_/X vssd1 vssd1 vccd1 vccd1 _07564_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_179_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06515_ _10095_/Q _06463_/A _08418_/A _06536_/A vssd1 vssd1 vccd1 vccd1 _06519_/A
+ sky130_fd_sc_hd__a22o_1
X_09303_ _09303_/A _09393_/A vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__nor2_2
X_07495_ _07485_/A _07539_/B _07868_/A _07515_/B _07494_/Y vssd1 vssd1 vccd1 vccd1
+ _07496_/B sky130_fd_sc_hd__o41a_1
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06446_ _06421_/Y _06442_/X _08351_/A _06442_/X _06445_/X vssd1 vssd1 vccd1 vccd1
+ _06447_/B sky130_fd_sc_hd__o221a_1
X_09234_ _05939_/X _09232_/Y _09233_/X vssd1 vssd1 vccd1 vccd1 _09234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09165_ _09165_/A vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__inv_2
X_08116_ _08783_/A vssd1 vssd1 vccd1 vccd1 _08116_/X sky130_fd_sc_hd__buf_2
X_06377_ _10246_/Q vssd1 vssd1 vccd1 vccd1 _06377_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ _09096_/A vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__buf_1
XFILLER_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05328_ _05328_/A vssd1 vssd1 vccd1 vccd1 _10342_/D sky130_fd_sc_hd__inv_2
XFILLER_162_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05259_ _10355_/Q vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__clkbuf_4
X_08047_ _07404_/A _07404_/B _07405_/B vssd1 vssd1 vccd1 vccd1 _08047_/X sky130_fd_sc_hd__a21bo_1
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _09997_/X _09408_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08949_ _08949_/A vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__inv_2
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10207_/CLK _10207_/D vssd1 vssd1 vccd1 vccd1 _10207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10138_ _10244_/CLK _10138_/D vssd1 vssd1 vccd1 vccd1 _10138_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_208_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _10202_/CLK _10069_/D vssd1 vssd1 vccd1 vccd1 _10069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06300_ _10131_/Q vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__inv_2
X_07280_ _07275_/X _07279_/X _07275_/X _07279_/X vssd1 vssd1 vccd1 vccd1 _07280_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_188_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06231_ _09679_/X _06203_/A _10080_/Q _06204_/A vssd1 vssd1 vccd1 vccd1 _10080_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06162_ _09646_/X _06156_/X _10128_/Q _06157_/X _05468_/X vssd1 vssd1 vccd1 vccd1
+ _10128_/D sky130_fd_sc_hd__o221a_1
X_05113_ _05161_/A vssd1 vssd1 vccd1 vccd1 _05113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06093_ _06101_/A vssd1 vssd1 vccd1 vccd1 _06093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05044_ _05968_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _05073_/A sky130_fd_sc_hd__or2_4
X_09921_ _07421_/Y _07422_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09921_/X sky130_fd_sc_hd__mux2_2
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09852_ _09851_/X _08282_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08803_ _08539_/A _08756_/Y _08765_/X _08802_/Y vssd1 vssd1 vccd1 vccd1 _08803_/X
+ sky130_fd_sc_hd__o211a_1
X_09783_ _10354_/Q _09782_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__mux2_1
X_08734_ _08734_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _08734_/X sky130_fd_sc_hd__or2_1
X_06995_ _06995_/A _06995_/B _07219_/B vssd1 vssd1 vccd1 vccd1 _06995_/X sky130_fd_sc_hd__or3_2
X_05946_ _05948_/A vssd1 vssd1 vccd1 vccd1 _05947_/A sky130_fd_sc_hd__inv_2
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08665_ _08086_/X _10053_/Q _08533_/A _10060_/Q _08644_/X vssd1 vssd1 vccd1 vccd1
+ _08666_/C sky130_fd_sc_hd__a221o_1
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05877_ _10254_/Q _05871_/X _05863_/X _06826_/A _05866_/X vssd1 vssd1 vccd1 vccd1
+ _10254_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08596_ _08596_/A _08596_/B _08596_/C vssd1 vssd1 vccd1 vccd1 _08596_/Y sky130_fd_sc_hd__nor3_1
XFILLER_198_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07616_ _07605_/C _07615_/A _07604_/A _07615_/Y vssd1 vssd1 vccd1 vccd1 _07616_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07547_ _07820_/A _07547_/B _07644_/A vssd1 vssd1 vccd1 vccd1 _07548_/B sky130_fd_sc_hd__and3_1
XFILLER_194_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07478_ _09934_/X vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__inv_2
XFILLER_194_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09217_ _09217_/A vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__inv_2
X_06429_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09148_ _09245_/C _09092_/Y _09093_/X _09098_/X vssd1 vssd1 vccd1 vccd1 _09193_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _09949_/X vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05800_ _05800_/A vssd1 vssd1 vccd1 vccd1 _05801_/A sky130_fd_sc_hd__inv_2
X_06780_ _10404_/Q _06812_/B _06779_/X vssd1 vssd1 vccd1 vccd1 _06780_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05731_ _07415_/A vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_208_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08450_ _08450_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08450_/Y sky130_fd_sc_hd__nor2_1
X_05662_ _05662_/A vssd1 vssd1 vccd1 vccd1 _05662_/Y sky130_fd_sc_hd__inv_2
X_08381_ _08415_/B vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__buf_1
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07401_ _07401_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07402_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05593_ _05673_/A _05673_/B vssd1 vssd1 vccd1 vccd1 _05672_/A sky130_fd_sc_hd__nand2_1
X_07332_ _07328_/Y _07329_/X _07330_/X _07331_/X vssd1 vssd1 vccd1 vccd1 _07362_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07263_ _07303_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07263_/X sky130_fd_sc_hd__and2_1
XFILLER_191_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06214_ _09692_/X _06210_/X _10093_/Q _06211_/X vssd1 vssd1 vccd1 vccd1 _10093_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09002_ _09000_/X _09001_/X _09000_/X _09001_/X vssd1 vssd1 vccd1 vccd1 _09003_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_07194_ _07192_/X _07193_/X _07192_/X _07193_/X vssd1 vssd1 vccd1 vccd1 _07194_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06145_ _09657_/X _06140_/X _10139_/Q _06141_/X _06135_/X vssd1 vssd1 vccd1 vccd1
+ _10139_/D sky130_fd_sc_hd__o221a_1
XFILLER_172_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06076_ _10178_/Q vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__buf_2
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05027_ _05016_/B _09940_/S _05024_/X _05013_/X _08623_/A vssd1 vssd1 vccd1 vccd1
+ _10448_/D sky130_fd_sc_hd__a221o_1
X_09904_ _07458_/Y _07459_/Y _10282_/Q vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__mux2_1
X_09835_ _10367_/Q _09834_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09766_ _08190_/X _10350_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09766_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06978_ _09884_/X vssd1 vssd1 vccd1 vccd1 _07223_/B sky130_fd_sc_hd__buf_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08717_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08717_/Y sky130_fd_sc_hd__nor2_1
X_09697_ _06534_/X input29/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09697_/X sky130_fd_sc_hd__mux2_1
X_05929_ _05922_/X _05927_/X _05089_/X _05928_/X _05918_/X vssd1 vssd1 vccd1 vccd1
+ _10233_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08648_ _08086_/X _10053_/Q _08081_/X _10054_/Q vssd1 vssd1 vccd1 vccd1 _08649_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _08594_/C _08577_/Y _08587_/B vssd1 vssd1 vccd1 vccd1 _08580_/C sky130_fd_sc_hd__o21ai_1
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07950_ _07716_/X _07755_/X _07716_/X _07755_/X vssd1 vssd1 vccd1 vccd1 _07950_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06901_ _06885_/X _06886_/X _06899_/X _06900_/X vssd1 vssd1 vccd1 vccd1 _06901_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07881_ _07881_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07882_/B sky130_fd_sc_hd__nor2_1
X_09620_ _09619_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09620_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06832_ _06827_/A _06827_/B _06828_/B vssd1 vssd1 vccd1 vccd1 _06832_/X sky130_fd_sc_hd__a21bo_1
X_06763_ _10390_/Q _06794_/B _06762_/Y vssd1 vssd1 vccd1 vccd1 _06763_/Y sky130_fd_sc_hd__o21ai_1
X_09551_ _08357_/Y _10115_/Q _09554_/S vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__mux2_1
X_08502_ _08502_/A vssd1 vssd1 vccd1 vccd1 _08502_/Y sky130_fd_sc_hd__inv_2
X_05714_ _10293_/Q _05701_/X _05788_/A _05705_/X _05711_/X vssd1 vssd1 vccd1 vccd1
+ _10293_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06694_ _06817_/B vssd1 vssd1 vccd1 vccd1 _06694_/Y sky130_fd_sc_hd__inv_2
X_09482_ _09480_/Y _09481_/X _09480_/Y _09481_/X vssd1 vssd1 vccd1 vccd1 _09482_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08433_ _09955_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08433_/Y sky130_fd_sc_hd__nor2_1
X_05645_ _05619_/X _05640_/Y _05641_/Y _08071_/A _05644_/X vssd1 vssd1 vccd1 vccd1
+ _05646_/B sky130_fd_sc_hd__o32a_1
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08364_ _10000_/X _08364_/B vssd1 vssd1 vccd1 vccd1 _08364_/Y sky130_fd_sc_hd__nor2_1
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05576_ _05574_/Y _05575_/Y _05574_/Y _05575_/Y vssd1 vssd1 vccd1 vccd1 _05576_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_07315_ _07027_/X _07314_/Y _07027_/X _07314_/Y vssd1 vssd1 vccd1 vccd1 _07315_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08295_ _08299_/B vssd1 vssd1 vccd1 vccd1 _08295_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07246_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__nor2_2
X_07177_ _07177_/A _07177_/B vssd1 vssd1 vccd1 vccd1 _07178_/B sky130_fd_sc_hd__or2_1
XFILLER_191_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06128_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06128_/X sky130_fd_sc_hd__clkbuf_2
X_06059_ _10186_/Q vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09818_ _08244_/Y _10363_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09818_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09749_ _09748_/X _10234_/Q _09997_/S vssd1 vssd1 vccd1 vccd1 _09749_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 io_wb_cs_i vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
Xinput29 io_wb_dat_i[19] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10422_/CLK _10386_/D vssd1 vssd1 vccd1 vccd1 _10386_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05430_ _05430_/A vssd1 vssd1 vccd1 vccd1 _10324_/D sky130_fd_sc_hd__inv_2
X_05361_ _05361_/A vssd1 vssd1 vccd1 vccd1 _10334_/D sky130_fd_sc_hd__inv_2
XFILLER_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07100_ _07100_/A _07116_/B vssd1 vssd1 vccd1 vccd1 _07100_/X sky130_fd_sc_hd__or2_1
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08080_ _10185_/Q vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__inv_2
X_05292_ _10335_/Q vssd1 vssd1 vccd1 vccd1 _05299_/A sky130_fd_sc_hd__inv_2
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ _08977_/X _08981_/X _08977_/X _08981_/X vssd1 vssd1 vccd1 vccd1 _08982_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07933_ _07931_/X _07932_/X _07931_/X _07932_/X vssd1 vssd1 vccd1 vccd1 _07933_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07864_ _07864_/A vssd1 vssd1 vccd1 vccd1 _07864_/Y sky130_fd_sc_hd__inv_2
X_09603_ _06614_/A _08616_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__mux2_1
X_06815_ _06818_/A _06815_/B vssd1 vssd1 vccd1 vccd1 _06815_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07795_ _10212_/Q _07788_/Y _07854_/D _07789_/Y _07794_/Y vssd1 vssd1 vccd1 vccd1
+ _07795_/X sky130_fd_sc_hd__a41o_1
X_09534_ _10379_/Q _10176_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09534_/X sky130_fd_sc_hd__mux2_1
X_06746_ _06739_/Y _06745_/X _06607_/Y _06736_/X vssd1 vssd1 vccd1 vccd1 _06746_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06677_ _10365_/Q _08734_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__or2_1
X_09465_ _09416_/X _09420_/X _09171_/X _09421_/X _09464_/Y vssd1 vssd1 vccd1 vccd1
+ _09465_/X sky130_fd_sc_hd__o221a_1
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ _09617_/X _08435_/B vssd1 vssd1 vccd1 vccd1 _08416_/X sky130_fd_sc_hd__and2_1
X_05628_ _10312_/Q vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__inv_2
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ _09391_/X _09395_/Y _09391_/X _09395_/Y vssd1 vssd1 vccd1 vccd1 _09396_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08347_ _09038_/A vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05559_ _05486_/A _05486_/B _05486_/Y vssd1 vssd1 vccd1 vccd1 _05559_/Y sky130_fd_sc_hd__a21oi_1
X_08278_ _08281_/B vssd1 vssd1 vccd1 vccd1 _08278_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07229_ _07226_/X _07228_/Y _07226_/X _07228_/Y vssd1 vssd1 vccd1 vccd1 _07229_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _10249_/CLK _10240_/D vssd1 vssd1 vccd1 vccd1 _10240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10171_ _10330_/CLK _10171_/D vssd1 vssd1 vccd1 vccd1 _10171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ _10442_/CLK _10438_/D vssd1 vssd1 vccd1 vccd1 _10438_/Q sky130_fd_sc_hd__dfxtp_1
X_10369_ _10436_/CLK _10369_/D vssd1 vssd1 vccd1 vccd1 _10369_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ _10381_/Q vssd1 vssd1 vccd1 vccd1 _06600_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _07574_/A _07569_/X _07573_/Y _07571_/A _07579_/Y vssd1 vssd1 vccd1 vccd1
+ _07580_/X sky130_fd_sc_hd__o32a_1
XFILLER_206_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06531_ _10098_/Q vssd1 vssd1 vccd1 vccd1 _08425_/A sky130_fd_sc_hd__inv_2
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09250_ _09246_/X _09249_/X _09246_/X _09249_/X vssd1 vssd1 vccd1 vccd1 _09250_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06462_ _06462_/A vssd1 vssd1 vccd1 vccd1 _06463_/A sky130_fd_sc_hd__clkbuf_2
X_08201_ _08204_/B vssd1 vssd1 vccd1 vccd1 _08201_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09181_ _09181_/A _09181_/B vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__or2_1
X_06393_ _06391_/X _06392_/Y _06391_/X _06392_/Y vssd1 vssd1 vccd1 vccd1 _06393_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05413_ _10327_/Q _05413_/B vssd1 vssd1 vccd1 vccd1 _05413_/Y sky130_fd_sc_hd__nor2_1
X_08132_ _06644_/Y _08801_/A _05273_/X _08130_/X _08131_/X vssd1 vssd1 vccd1 vccd1
+ _08143_/B sky130_fd_sc_hd__o221a_1
X_05344_ _10338_/Q _05344_/B vssd1 vssd1 vccd1 vccd1 _05344_/Y sky130_fd_sc_hd__nor2_1
X_05275_ _05101_/X _05215_/X _05273_/X _05216_/X _05274_/X vssd1 vssd1 vccd1 vccd1
+ _10348_/D sky130_fd_sc_hd__a221o_1
XFILLER_146_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _08063_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08063_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07014_ _07227_/B _06991_/Y _06995_/A vssd1 vssd1 vccd1 vccd1 _07014_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_161_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ _08998_/A _09977_/X _08912_/A _09089_/B vssd1 vssd1 vccd1 vccd1 _08965_/X
+ sky130_fd_sc_hd__o22a_1
X_07916_ _07916_/A _07916_/B _07916_/C vssd1 vssd1 vccd1 vccd1 _07916_/X sky130_fd_sc_hd__or3_2
XFILLER_124_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08896_ _08894_/Y _08893_/X _08909_/A vssd1 vssd1 vccd1 vccd1 _08896_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07847_ _07835_/A _07835_/B _07881_/A vssd1 vssd1 vccd1 vccd1 _07850_/A sky130_fd_sc_hd__a21o_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07778_ _07687_/B _07769_/X _07919_/A _07776_/X _07777_/X vssd1 vssd1 vccd1 vccd1
+ _07778_/X sky130_fd_sc_hd__o221a_1
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06729_ _10358_/Q _06670_/B _06727_/Y vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__a21oi_2
X_09517_ _09516_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09517_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _10228_/Q _09397_/Y _05941_/X _09398_/Y _09402_/Y vssd1 vssd1 vccd1 vccd1
+ _09448_/X sky130_fd_sc_hd__a41o_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _09380_/A _09380_/B vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__and2_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10223_ _10225_/CLK _10223_/D vssd1 vssd1 vccd1 vccd1 _10223_/Q sky130_fd_sc_hd__dfxtp_1
X_10154_ _10330_/CLK _10154_/D vssd1 vssd1 vccd1 vccd1 _10154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ _10450_/CLK _10085_/D vssd1 vssd1 vccd1 vccd1 _10085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05060_ _10436_/Q _05055_/X input36/X _05057_/X _05053_/X vssd1 vssd1 vccd1 vccd1
+ _10436_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08750_ _10191_/Q _08747_/B _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08823_/C
+ sky130_fd_sc_hd__a22o_1
X_05962_ _10219_/Q vssd1 vssd1 vccd1 vccd1 _07108_/A sky130_fd_sc_hd__clkbuf_2
X_08681_ _08654_/X _08667_/Y _08705_/B vssd1 vssd1 vccd1 vccd1 _08681_/X sky130_fd_sc_hd__o21ba_1
X_05893_ _06082_/B _05944_/B vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__or2_4
X_07701_ _07695_/A _07722_/A _07694_/Y _07692_/A _07700_/Y vssd1 vssd1 vccd1 vccd1
+ _07701_/X sky130_fd_sc_hd__o32a_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07632_ _07577_/A _07577_/B _07578_/B vssd1 vssd1 vccd1 vccd1 _07632_/X sky130_fd_sc_hd__a21bo_1
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09302_ _09296_/X _09301_/X _09296_/X _09301_/X vssd1 vssd1 vccd1 vccd1 _09392_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__or2_1
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06514_ _10095_/Q vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__inv_2
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _07498_/C _07494_/B vssd1 vssd1 vccd1 vccd1 _07494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06445_ _06445_/A _06445_/B vssd1 vssd1 vccd1 vccd1 _06445_/X sky130_fd_sc_hd__or2_1
X_09233_ _09289_/A _09945_/X vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__or2_1
X_09164_ _08846_/X _08867_/X _08846_/X _08867_/X vssd1 vssd1 vccd1 vccd1 _09165_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _08191_/A vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06376_ _06372_/Y _06375_/X _06372_/Y _06375_/X vssd1 vssd1 vccd1 vccd1 _06376_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09095_ _09095_/A vssd1 vssd1 vccd1 vccd1 _09095_/Y sky130_fd_sc_hd__inv_2
X_05327_ _05320_/B _05282_/X _05326_/Y _05322_/X _05306_/A vssd1 vssd1 vccd1 vccd1
+ _05328_/A sky130_fd_sc_hd__o32a_1
XFILLER_162_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05258_ input50/X _05251_/X _08762_/A _05252_/X _05253_/X vssd1 vssd1 vccd1 vccd1
+ _10356_/D sky130_fd_sc_hd__a221o_1
X_08046_ _08019_/A _08019_/B _08020_/B vssd1 vssd1 vccd1 vccd1 _08046_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05189_ _05189_/A vssd1 vssd1 vccd1 vccd1 _05189_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _08363_/X _06311_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09997_/X sky130_fd_sc_hd__mux2_1
X_08948_ _08979_/A _08947_/B _08947_/X vssd1 vssd1 vccd1 vccd1 _08949_/A sky130_fd_sc_hd__a21bo_1
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08879_ _05581_/X _07425_/A _08858_/Y vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__o21ai_2
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10206_ _10207_/CLK _10206_/D vssd1 vssd1 vccd1 vccd1 _10206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10137_ _10244_/CLK _10137_/D vssd1 vssd1 vccd1 vccd1 _10137_/Q sky130_fd_sc_hd__dfxtp_1
X_10068_ _10202_/CLK _10068_/D vssd1 vssd1 vccd1 vccd1 _10068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06230_ _09680_/X _06224_/X _10081_/Q _06225_/X vssd1 vssd1 vccd1 vccd1 _10081_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06161_ _09647_/X _06156_/X _10129_/Q _06157_/X _06154_/X vssd1 vssd1 vccd1 vccd1
+ _10129_/D sky130_fd_sc_hd__o221a_1
X_05112_ _05203_/A _09899_/S vssd1 vssd1 vccd1 vccd1 _05161_/A sky130_fd_sc_hd__or2_4
X_06092_ _10172_/Q _06101_/A _10344_/Q _06102_/A _05993_/X vssd1 vssd1 vccd1 vccd1
+ _10172_/D sky130_fd_sc_hd__o221a_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05043_ _08329_/D _08324_/A _06082_/B vssd1 vssd1 vccd1 vccd1 _09981_/S sky130_fd_sc_hd__or3_4
X_09920_ _07415_/Y _07420_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09920_/X sky130_fd_sc_hd__mux2_2
X_09851_ _10371_/Q _09850_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08802_ _06253_/A _08766_/Y _08769_/X _08800_/Y _08801_/X vssd1 vssd1 vccd1 vccd1
+ _08802_/Y sky130_fd_sc_hd__o221ai_2
X_09782_ _08207_/X _10354_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09782_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06994_ _06984_/X _06990_/Y _06984_/A _06990_/Y vssd1 vssd1 vccd1 vccd1 _06995_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_08733_ _08733_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__and2_1
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05945_ _05968_/A _08317_/A vssd1 vssd1 vccd1 vccd1 _05948_/A sky130_fd_sc_hd__or2_4
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08664_ _08664_/A _08664_/B _08649_/B _08652_/Y vssd1 vssd1 vccd1 vccd1 _08666_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05876_ _05876_/A vssd1 vssd1 vccd1 vccd1 _06826_/A sky130_fd_sc_hd__inv_2
XFILLER_198_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08595_ _08595_/A _08595_/B _08595_/C _08580_/B vssd1 vssd1 vccd1 vccd1 _08597_/B
+ sky130_fd_sc_hd__or4b_4
X_07615_ _07615_/A vssd1 vssd1 vccd1 vccd1 _07615_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07546_ _07591_/A _09936_/X vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__or2_1
XFILLER_194_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ _09159_/X _09215_/X _09159_/X _09215_/X vssd1 vssd1 vccd1 vccd1 _09217_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07477_ _07477_/A _07476_/X vssd1 vssd1 vccd1 vccd1 _07477_/X sky130_fd_sc_hd__or2b_1
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06428_ _10082_/Q _06443_/A _08351_/A _06442_/A vssd1 vssd1 vccd1 vccd1 _06445_/B
+ sky130_fd_sc_hd__a22o_1
X_09147_ _09145_/X _09146_/X _09145_/X _09146_/X vssd1 vssd1 vccd1 vccd1 _09147_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
X_06359_ _10137_/Q vssd1 vssd1 vccd1 vccd1 _08390_/A sky130_fd_sc_hd__inv_2
XFILLER_175_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09078_ _09078_/A vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08029_ _07413_/A _07413_/B _07413_/Y vssd1 vssd1 vccd1 vccd1 _08029_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05730_ _10270_/Q vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_208_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05661_ _10306_/Q _05467_/X _05637_/X _05659_/Y _05660_/X vssd1 vssd1 vccd1 vccd1
+ _10306_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08380_ _08380_/A vssd1 vssd1 vccd1 vccd1 _08415_/B sky130_fd_sc_hd__buf_1
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07400_ _07400_/A vssd1 vssd1 vccd1 vccd1 _07401_/B sky130_fd_sc_hd__inv_2
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05592_ _09939_/X _05572_/X _05679_/A vssd1 vssd1 vccd1 vccd1 _05673_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07331_ _07256_/X _07304_/X _07256_/X _07304_/X vssd1 vssd1 vccd1 vccd1 _07331_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07262_ _07258_/X _07259_/X _07260_/X _07261_/X vssd1 vssd1 vccd1 vccd1 _07303_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06213_ _09693_/X _06210_/X _10094_/Q _06211_/X vssd1 vssd1 vccd1 vccd1 _10094_/D
+ sky130_fd_sc_hd__a22o_1
X_09001_ _09029_/A _09938_/X _09001_/C vssd1 vssd1 vccd1 vccd1 _09001_/X sky130_fd_sc_hd__or3_1
X_07193_ _07178_/B _07180_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07193_/X sky130_fd_sc_hd__o21a_1
XFILLER_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06144_ _09658_/X _06140_/X _10140_/Q _06141_/X _06135_/X vssd1 vssd1 vccd1 vccd1
+ _10140_/D sky130_fd_sc_hd__o221a_1
XFILLER_172_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06075_ _09769_/X _06067_/X _10179_/Q _06069_/X _06070_/X vssd1 vssd1 vccd1 vccd1
+ _10179_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05026_ _06099_/A vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__clkbuf_2
X_09903_ _09281_/X _09279_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__mux2_1
X_09834_ _08263_/Y _10367_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ _09764_/X input41/X _09781_/S vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__mux2_1
X_06977_ _06977_/A vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__buf_2
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08716_ _08713_/A _08717_/B _06628_/Y _08715_/Y vssd1 vssd1 vccd1 vccd1 _08716_/X
+ sky130_fd_sc_hd__o22a_1
X_09696_ _06530_/Y input28/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09696_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05928_ _05928_/A vssd1 vssd1 vccd1 vccd1 _05928_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_199_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ _08093_/X _10055_/Q _08081_/X _10054_/Q vssd1 vssd1 vccd1 vccd1 _08664_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05859_ _10259_/Q _05851_/X _05842_/X _06835_/A _05845_/X vssd1 vssd1 vccd1 vccd1
+ _10259_/D sky130_fd_sc_hd__o221a_1
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _08578_/A _08578_/B vssd1 vssd1 vccd1 vccd1 _08587_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ _07529_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07529_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06900_ _06885_/X _06886_/X _06885_/X _06886_/X vssd1 vssd1 vccd1 vccd1 _06900_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07880_ _07845_/A _07851_/A _07845_/Y vssd1 vssd1 vccd1 vccd1 _07880_/X sky130_fd_sc_hd__a21o_1
X_06831_ _06828_/A _06828_/B _06829_/B vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__a21bo_1
X_06762_ _06643_/Y _06793_/B _06761_/X vssd1 vssd1 vccd1 vccd1 _06762_/Y sky130_fd_sc_hd__o21ai_1
X_09550_ _09549_/X _10351_/Q _09982_/S vssd1 vssd1 vccd1 vccd1 _09550_/X sky130_fd_sc_hd__mux2_1
X_08501_ _10069_/Q _08487_/B _08488_/B vssd1 vssd1 vccd1 vccd1 _08599_/B sky130_fd_sc_hd__a21bo_1
X_09481_ _09427_/X _09428_/X _09429_/X _09432_/Y _09434_/X vssd1 vssd1 vccd1 vccd1
+ _09481_/X sky130_fd_sc_hd__o221a_1
X_05713_ _10277_/Q vssd1 vssd1 vccd1 vccd1 _05788_/A sky130_fd_sc_hd__buf_2
X_06693_ _10377_/Q _08707_/A _06690_/Y vssd1 vssd1 vccd1 vccd1 _06817_/B sky130_fd_sc_hd__a21oi_2
X_08432_ _08432_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08432_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05644_ _06126_/A vssd1 vssd1 vccd1 vccd1 _05644_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08363_ _08363_/A _08386_/B vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__or2_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05575_ _05497_/A _05497_/B _05497_/Y vssd1 vssd1 vccd1 vccd1 _05575_/Y sky130_fd_sc_hd__a21oi_1
X_08294_ _08294_/A _08294_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__or2_1
XFILLER_149_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07314_ _07044_/X _07313_/Y _07044_/X _07313_/Y vssd1 vssd1 vccd1 vccd1 _07314_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_176_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07245_ _07245_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07246_/B sky130_fd_sc_hd__nand2_2
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07176_ _07176_/A _07176_/B vssd1 vssd1 vccd1 vccd1 _07177_/B sky130_fd_sc_hd__or2_1
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06127_ _10149_/Q _06126_/X _10321_/Q _06122_/X _06120_/X vssd1 vssd1 vccd1 vccd1
+ _10149_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06058_ _09801_/X _06054_/X _06253_/A _06056_/X _06057_/X vssd1 vssd1 vccd1 vccd1
+ _10187_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05009_ _06183_/A _08324_/C _08329_/D vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__or3_4
X_09817_ _09816_/X input25/X _09821_/S vssd1 vssd1 vccd1 vccd1 _09817_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ _10127_/Q _10266_/Q _09748_/S vssd1 vssd1 vccd1 vccd1 _09748_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09679_ _06419_/X input30/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_wb_dat_i[0] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_6
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10385_ _10422_/CLK _10385_/D vssd1 vssd1 vccd1 vccd1 _10385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05360_ _05356_/B _05333_/A _05359_/X _05336_/A _05298_/C vssd1 vssd1 vccd1 vccd1
+ _05361_/A sky130_fd_sc_hd__o32a_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05291_ _10336_/Q vssd1 vssd1 vccd1 vccd1 _05300_/A sky130_fd_sc_hd__inv_2
XFILLER_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07030_ _05943_/X _06868_/Y _07028_/X _07029_/Y vssd1 vssd1 vccd1 vccd1 _07030_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08981_ _05931_/X _09168_/A _09010_/C _08980_/X vssd1 vssd1 vccd1 vccd1 _08981_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07932_ _07915_/A _07915_/B _07915_/X vssd1 vssd1 vccd1 vccd1 _07932_/X sky130_fd_sc_hd__a21bo_1
X_07863_ _07794_/A _07794_/B _07794_/Y vssd1 vssd1 vccd1 vccd1 _07863_/X sky130_fd_sc_hd__a21o_1
X_06814_ _06814_/A _06814_/B vssd1 vssd1 vccd1 vccd1 _06814_/Y sky130_fd_sc_hd__nor2_1
X_09602_ _09601_/X _06628_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09602_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09533_ _09532_/X _06634_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09533_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07794_/Y sky130_fd_sc_hd__nor2_1
X_06745_ _10382_/Q _06740_/Y _10381_/Q _06742_/Y _06744_/X vssd1 vssd1 vccd1 vccd1
+ _06745_/X sky130_fd_sc_hd__o221a_1
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06676_ _10364_/Q _08738_/A vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__or2_2
X_09464_ _09464_/A vssd1 vssd1 vccd1 vccd1 _09464_/Y sky130_fd_sc_hd__inv_2
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05627_ _05627_/A _05627_/B vssd1 vssd1 vccd1 vccd1 _05627_/Y sky130_fd_sc_hd__nor2_1
X_09395_ _09395_/A vssd1 vssd1 vccd1 vccd1 _09395_/Y sky130_fd_sc_hd__inv_2
X_08415_ _08415_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ _08912_/A vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05558_ _05558_/A vssd1 vssd1 vccd1 vccd1 _05558_/Y sky130_fd_sc_hd__inv_2
X_08277_ _08600_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08281_/B sky130_fd_sc_hd__or2_1
XFILLER_192_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05489_ _05489_/A _05489_/B vssd1 vssd1 vccd1 vccd1 _05489_/Y sky130_fd_sc_hd__nor2_1
X_07228_ _07228_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07228_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07159_ _07164_/A _09885_/X vssd1 vssd1 vccd1 vccd1 _07160_/A sky130_fd_sc_hd__or2_2
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10170_ _10330_/CLK _10170_/D vssd1 vssd1 vccd1 vccd1 _10170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10437_ _10437_/CLK _10437_/D vssd1 vssd1 vccd1 vccd1 _10437_/Q sky130_fd_sc_hd__dfxtp_1
X_10368_ _10436_/CLK _10368_/D vssd1 vssd1 vccd1 vccd1 _10368_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10299_ _10422_/CLK _10299_/D vssd1 vssd1 vccd1 vccd1 _10299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06530_ _06539_/A _06529_/X _06539_/A _06529_/X vssd1 vssd1 vccd1 vccd1 _06530_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06461_ _06461_/A vssd1 vssd1 vccd1 vccd1 _06462_/A sky130_fd_sc_hd__clkbuf_2
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08204_/B sky130_fd_sc_hd__or2_1
X_05412_ _05412_/A vssd1 vssd1 vccd1 vccd1 _05413_/B sky130_fd_sc_hd__inv_2
XFILLER_178_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09180_ _09343_/A _09247_/A _09180_/C vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__or3_1
X_06392_ _06377_/Y _10139_/Q _06384_/X vssd1 vssd1 vccd1 vccd1 _06392_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ _10370_/Q _08079_/X _06722_/Y _06047_/X vssd1 vssd1 vccd1 vccd1 _08131_/X
+ sky130_fd_sc_hd__o22a_1
X_05343_ _05343_/A vssd1 vssd1 vccd1 vccd1 _05344_/B sky130_fd_sc_hd__inv_2
X_05274_ _05274_/A vssd1 vssd1 vccd1 vccd1 _05274_/X sky130_fd_sc_hd__clkbuf_4
X_08062_ _08062_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07013_ _06997_/X _07012_/X _06997_/X _07012_/X vssd1 vssd1 vccd1 vccd1 _07013_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08964_ _09985_/X vssd1 vssd1 vccd1 vccd1 _09089_/B sky130_fd_sc_hd__buf_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07915_ _07915_/A _07915_/B vssd1 vssd1 vccd1 vccd1 _07915_/X sky130_fd_sc_hd__or2_1
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__or2_2
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07846_ _07846_/A vssd1 vssd1 vccd1 vccd1 _07881_/A sky130_fd_sc_hd__inv_2
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07777_ _07777_/A _07777_/B _07777_/C _07770_/X vssd1 vssd1 vccd1 vccd1 _07777_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_140_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06728_ _06642_/Y _06727_/Y _06672_/B vssd1 vssd1 vccd1 vccd1 _06795_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09516_ _09515_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ _09447_/A _09922_/X vssd1 vssd1 vccd1 vccd1 _09447_/Y sky130_fd_sc_hd__nor2_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _05024_/A _06657_/Y _06658_/Y _08625_/B vssd1 vssd1 vccd1 vccd1 _06660_/A
+ sky130_fd_sc_hd__o22a_1
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09378_ _09286_/X _09307_/X _09308_/X _09325_/X vssd1 vssd1 vccd1 vccd1 _09380_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08329_ input9/X input6/X _08329_/C _08329_/D vssd1 vssd1 vccd1 vccd1 _09600_/S sky130_fd_sc_hd__or4_4
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10222_ _10225_/CLK _10222_/D vssd1 vssd1 vccd1 vccd1 _10222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10153_ _10329_/CLK _10153_/D vssd1 vssd1 vccd1 vccd1 _10153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10084_ _10244_/CLK _10084_/D vssd1 vssd1 vccd1 vccd1 _10084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05961_ _10220_/Q _05947_/A input41/X _05948_/A _05960_/X vssd1 vssd1 vccd1 vccd1
+ _10220_/D sky130_fd_sc_hd__o221a_1
X_07700_ _07700_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07700_/Y sky130_fd_sc_hd__nor2_1
X_08680_ _08680_/A _08680_/B _08678_/X _08679_/X vssd1 vssd1 vccd1 vccd1 _08705_/B
+ sky130_fd_sc_hd__or4bb_4
X_05892_ _10250_/Q _05891_/X _05699_/X _07152_/D _05885_/X vssd1 vssd1 vccd1 vccd1
+ _10250_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07631_ _07606_/X _07628_/X _07606_/X _07628_/X vssd1 vssd1 vccd1 vccd1 _07631_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07562_ _07550_/A _07550_/B _07550_/X vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__a21bo_1
X_06513_ _06516_/D _06512_/Y _06516_/D _06512_/Y vssd1 vssd1 vccd1 vccd1 _06513_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09301_ _09298_/Y _09300_/X _09298_/Y _09300_/X vssd1 vssd1 vccd1 vccd1 _09301_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07493_ _07885_/C _07566_/B _07493_/C vssd1 vssd1 vccd1 vccd1 _07494_/B sky130_fd_sc_hd__and3_1
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09232_ _09292_/B vssd1 vssd1 vccd1 vccd1 _09232_/Y sky130_fd_sc_hd__inv_2
X_06444_ _08357_/A _06442_/X _10083_/Q _06460_/A vssd1 vssd1 vccd1 vccd1 _06447_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ _09162_/A _09162_/B _09218_/A vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__a21bo_1
X_06375_ _10244_/Q _08390_/A _06362_/Y _06367_/A vssd1 vssd1 vccd1 vccd1 _06375_/X
+ sky130_fd_sc_hd__o22a_1
X_08114_ _10179_/Q vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__inv_2
XFILLER_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05326_ _10342_/Q _05326_/B vssd1 vssd1 vccd1 vccd1 _05326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09094_ _09094_/A _09050_/X vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__or2b_1
XFILLER_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05257_ _10356_/Q vssd1 vssd1 vccd1 vccd1 _08762_/A sky130_fd_sc_hd__buf_2
X_08045_ _07405_/A _07405_/B _07406_/B vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__a21bo_1
XFILLER_150_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05188_ _05185_/X _10393_/Q _05186_/X _09612_/X _05078_/X vssd1 vssd1 vccd1 vccd1
+ _10393_/D sky130_fd_sc_hd__o221a_1
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _08055_/Y _07385_/X _10022_/S vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08947_ _08979_/A _08947_/B vssd1 vssd1 vccd1 vccd1 _08947_/X sky130_fd_sc_hd__or2_1
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08878_ _09008_/B vssd1 vssd1 vccd1 vccd1 _09042_/B sky130_fd_sc_hd__buf_2
XFILLER_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07829_ _07829_/A vssd1 vssd1 vccd1 vccd1 _07830_/C sky130_fd_sc_hd__inv_2
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10205_/CLK _10205_/D vssd1 vssd1 vccd1 vccd1 _10205_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_180_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _10244_/CLK _10136_/D vssd1 vssd1 vccd1 vccd1 _10136_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10067_ _10202_/CLK _10067_/D vssd1 vssd1 vccd1 vccd1 _10067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06160_ _09648_/X _06156_/X _10130_/Q _06157_/X _06154_/X vssd1 vssd1 vccd1 vccd1
+ _10130_/D sky130_fd_sc_hd__o221a_1
XFILLER_156_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06091_ _10173_/Q _06088_/X _10345_/Q _06089_/X _05993_/X vssd1 vssd1 vccd1 vccd1
+ _10173_/D sky130_fd_sc_hd__o221a_1
X_05111_ _05369_/A vssd1 vssd1 vccd1 vccd1 _05203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05042_ input12/X _05775_/A input11/X vssd1 vssd1 vccd1 vccd1 _06082_/B sky130_fd_sc_hd__or3b_4
XFILLER_171_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09850_ _08280_/Y _10371_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09850_/X sky130_fd_sc_hd__mux2_1
X_08801_ _08801_/A _08801_/B vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__or2_1
X_09781_ _09780_/X input47/X _09781_/S vssd1 vssd1 vccd1 vccd1 _09781_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06993_ _07227_/B _06993_/B vssd1 vssd1 vccd1 vccd1 _06995_/A sky130_fd_sc_hd__or2_1
X_08732_ _10366_/Q _08731_/X _08729_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08733_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_05944_ _08324_/C _05944_/B vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__or2_4
X_08663_ _08656_/X _08661_/Y _08704_/A vssd1 vssd1 vccd1 vccd1 _08663_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05875_ _05810_/X _05817_/X _05810_/X _05817_/X vssd1 vssd1 vccd1 vccd1 _05876_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_198_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08594_ _08594_/A _08594_/B _08594_/C _08593_/X vssd1 vssd1 vccd1 vccd1 _08595_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _10213_/Q _07687_/B _07625_/A vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__and3_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07545_ _07591_/A _09935_/X vssd1 vssd1 vccd1 vccd1 _07552_/C sky130_fd_sc_hd__nor2_1
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07476_ _07766_/A _07504_/B _07806_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _07476_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_179_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _09213_/X _09214_/X _09213_/X _09214_/X vssd1 vssd1 vccd1 vccd1 _09215_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06427_ _10082_/Q vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__inv_2
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09146_ _09009_/X _09095_/A _09252_/A _09245_/B vssd1 vssd1 vccd1 vccd1 _09146_/X
+ sky130_fd_sc_hd__a211o_2
X_06358_ _06353_/A _06357_/X _06353_/A _06357_/X vssd1 vssd1 vccd1 vccd1 _06358_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05309_ _05309_/A _05309_/B vssd1 vssd1 vccd1 vccd1 _05312_/A sky130_fd_sc_hd__or2_1
X_09077_ _09077_/A _09031_/X vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__or2b_1
X_06289_ _06285_/A _06288_/A _06283_/A _06288_/Y vssd1 vssd1 vccd1 vccd1 _06289_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08028_ _08027_/A _08027_/B _07984_/Y _07984_/A _08027_/Y vssd1 vssd1 vccd1 vccd1
+ _08028_/X sky130_fd_sc_hd__o32a_1
XFILLER_190_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09979_ _06614_/C _08304_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09979_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10119_ _10334_/CLK _10119_/D vssd1 vssd1 vccd1 vccd1 _10119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05660_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05660_/X sky130_fd_sc_hd__buf_2
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05591_ _05680_/A _05680_/B vssd1 vssd1 vccd1 vccd1 _05679_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _07328_/Y _07329_/X _07328_/Y _07329_/X vssd1 vssd1 vccd1 vccd1 _07330_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_204_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09000_ _09069_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09000_/X sky130_fd_sc_hd__or2_2
X_07261_ _07258_/X _07259_/X _07258_/X _07259_/X vssd1 vssd1 vccd1 vccd1 _07261_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06212_ _09694_/X _06210_/X _10095_/Q _06211_/X vssd1 vssd1 vccd1 vccd1 _10095_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07192_ _07182_/A _07182_/B _07182_/Y vssd1 vssd1 vccd1 vccd1 _07192_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06143_ _09659_/X _06140_/X _10141_/Q _06141_/X _06135_/X vssd1 vssd1 vccd1 vccd1
+ _10141_/D sky130_fd_sc_hd__o221a_1
XFILLER_172_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06074_ _09773_/X _06067_/X _10180_/Q _06069_/X _06070_/X vssd1 vssd1 vccd1 vccd1
+ _10180_/D sky130_fd_sc_hd__o221a_1
X_09902_ _09333_/X _09331_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09902_/X sky130_fd_sc_hd__mux2_2
XFILLER_132_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05025_ input52/X vssd1 vssd1 vccd1 vccd1 _06099_/A sky130_fd_sc_hd__buf_2
X_09833_ _09832_/X input29/X _09849_/S vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09764_ _09763_/X _08189_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09764_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06976_ _06976_/A vssd1 vssd1 vccd1 vccd1 _07311_/B sky130_fd_sc_hd__inv_2
X_08715_ _08715_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08715_/Y sky130_fd_sc_hd__nor2_1
X_09695_ _06524_/X input27/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09695_/X sky130_fd_sc_hd__mux2_1
X_05927_ _05927_/A vssd1 vssd1 vccd1 vccd1 _05927_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ _08160_/X _10056_/Q _08093_/X _10055_/Q vssd1 vssd1 vccd1 vccd1 _08646_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05858_ _05858_/A vssd1 vssd1 vccd1 vccd1 _06835_/A sky130_fd_sc_hd__inv_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _08537_/X _08593_/C _08575_/Y _08595_/A vssd1 vssd1 vccd1 vccd1 _08577_/Y
+ sky130_fd_sc_hd__a31oi_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05789_ _10260_/Q vssd1 vssd1 vccd1 vccd1 _05853_/B sky130_fd_sc_hd__inv_2
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _07528_/A _07528_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__nor2_2
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07459_ _07458_/Y _07442_/Y _07455_/B vssd1 vssd1 vccd1 vccd1 _07459_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _09129_/A vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06830_ _06829_/A _06829_/B _06834_/B vssd1 vssd1 vccd1 vccd1 _06830_/X sky130_fd_sc_hd__a21bo_1
X_06761_ _06643_/Y _06793_/B _06759_/Y _06760_/Y vssd1 vssd1 vccd1 vccd1 _06761_/X
+ sky130_fd_sc_hd__a22o_1
X_08500_ _10070_/Q _08488_/B _08489_/B vssd1 vssd1 vccd1 vccd1 _08500_/X sky130_fd_sc_hd__a21bo_1
X_06692_ _06818_/B vssd1 vssd1 vccd1 vccd1 _06692_/Y sky130_fd_sc_hd__inv_2
X_09480_ _09414_/X _09425_/X _09426_/X _09435_/X vssd1 vssd1 vccd1 vccd1 _09480_/Y
+ sky130_fd_sc_hd__o22ai_2
X_05712_ _10294_/Q _05701_/X _08845_/B _05705_/X _05711_/X vssd1 vssd1 vccd1 vccd1
+ _10294_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ _09953_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__nor2_1
X_05643_ _05750_/A vssd1 vssd1 vccd1 vccd1 _06126_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08362_ _08413_/B vssd1 vssd1 vccd1 vccd1 _08386_/B sky130_fd_sc_hd__buf_1
X_05574_ _05574_/A vssd1 vssd1 vccd1 vccd1 _05574_/Y sky130_fd_sc_hd__inv_2
X_08293_ _08293_/A vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07313_ _07310_/X _07312_/X _07310_/X _07312_/X vssd1 vssd1 vccd1 vccd1 _07313_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07244_ _07223_/C _07220_/B _07220_/Y vssd1 vssd1 vccd1 vccd1 _07245_/B sky130_fd_sc_hd__o21a_1
XFILLER_191_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _07155_/C _07151_/X _07155_/C _07151_/X vssd1 vssd1 vccd1 vccd1 _07176_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_191_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06126_ _06126_/A vssd1 vssd1 vccd1 vccd1 _06126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06057_ _06070_/A vssd1 vssd1 vccd1 vccd1 _06057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05008_ input16/X _06081_/B _06081_/A vssd1 vssd1 vccd1 vccd1 _08329_/D sky130_fd_sc_hd__or3_4
XFILLER_113_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ _09815_/X _08243_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09747_ _10412_/Q _08060_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06959_ _06940_/X _06952_/X _06953_/X _06958_/X vssd1 vssd1 vccd1 vccd1 _06959_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09678_ _06416_/Y input19/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _05024_/X _08146_/Y _08626_/Y _08628_/Y vssd1 vssd1 vccd1 vccd1 _08629_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ _10422_/CLK _10384_/D vssd1 vssd1 vccd1 vccd1 _10384_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05290_ _10337_/Q vssd1 vssd1 vccd1 vccd1 _05301_/A sky130_fd_sc_hd__inv_2
XFILLER_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _09354_/A _09045_/B _09252_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _08980_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07931_ _07889_/X _07894_/X _07889_/X _07894_/X vssd1 vssd1 vccd1 vccd1 _07931_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_95_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07862_ _07831_/X _07852_/X _07831_/X _07852_/X vssd1 vssd1 vccd1 vccd1 _07862_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06813_ _06814_/A _06813_/B vssd1 vssd1 vccd1 vccd1 _06813_/Y sky130_fd_sc_hd__nor2_1
X_09601_ _06615_/B _08134_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09601_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09532_ _05172_/Y _08253_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__mux2_1
X_07793_ _07855_/A _09924_/X _07792_/X vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__or3b_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06744_ _10380_/Q _06647_/A _10381_/Q _06742_/Y _06743_/X vssd1 vssd1 vccd1 vccd1
+ _06744_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06675_ _10363_/Q _08742_/A vssd1 vssd1 vccd1 vccd1 _08738_/A sky130_fd_sc_hd__or2_1
X_09463_ _10232_/Q _09405_/Y _05933_/X _09232_/Y _09409_/Y vssd1 vssd1 vccd1 vccd1
+ _09463_/X sky130_fd_sc_hd__a41o_1
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05626_ _05626_/A vssd1 vssd1 vccd1 vccd1 _05626_/Y sky130_fd_sc_hd__inv_2
X_09394_ _09303_/A _09392_/Y _09350_/Y _09347_/Y _09393_/X vssd1 vssd1 vccd1 vccd1
+ _09395_/A sky130_fd_sc_hd__a32o_1
X_08414_ _09521_/X _08414_/B vssd1 vssd1 vccd1 vccd1 _08414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05557_ _09947_/X _05556_/X _09947_/X _05556_/X vssd1 vssd1 vccd1 vccd1 _05655_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08345_ _10229_/Q vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__inv_2
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08276_ _06265_/A _06265_/B _08275_/Y vssd1 vssd1 vccd1 vccd1 _08276_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05488_ _09991_/X vssd1 vssd1 vccd1 vccd1 _05489_/B sky130_fd_sc_hd__inv_2
XFILLER_138_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07227_ _07234_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07228_/B sky130_fd_sc_hd__or2_2
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07158_ _07145_/X _07146_/X _07156_/X _07157_/X vssd1 vssd1 vccd1 vccd1 _07158_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06109_ _10332_/Q _06088_/X _10160_/Q _06089_/X _05105_/A vssd1 vssd1 vccd1 vccd1
+ _10160_/D sky130_fd_sc_hd__a221o_1
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07089_ _07089_/A _07095_/A vssd1 vssd1 vccd1 vccd1 _07089_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10436_ _10436_/CLK _10436_/D vssd1 vssd1 vccd1 vccd1 _10436_/Q sky130_fd_sc_hd__dfxtp_1
X_10367_ _10399_/CLK _10367_/D vssd1 vssd1 vccd1 vccd1 _10367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10298_ _10298_/CLK _10298_/D vssd1 vssd1 vccd1 vccd1 _10298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06460_ _06460_/A vssd1 vssd1 vccd1 vccd1 _06461_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05411_ _05411_/A vssd1 vssd1 vccd1 vccd1 _10328_/D sky130_fd_sc_hd__inv_2
X_08130_ _08791_/A vssd1 vssd1 vccd1 vccd1 _08130_/X sky130_fd_sc_hd__clkbuf_2
X_06391_ _06391_/A _06391_/B vssd1 vssd1 vccd1 vccd1 _06391_/X sky130_fd_sc_hd__or2_1
XFILLER_186_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05342_ _05342_/A vssd1 vssd1 vccd1 vccd1 _10339_/D sky130_fd_sc_hd__inv_2
X_05273_ _10348_/Q vssd1 vssd1 vccd1 vccd1 _05273_/X sky130_fd_sc_hd__buf_2
X_08061_ _08061_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07012_ _05943_/X _06999_/Y _07008_/Y _07011_/X vssd1 vssd1 vccd1 vccd1 _07012_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ _09977_/X vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__inv_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07914_ _07909_/X _07911_/Y _07912_/X _07913_/Y vssd1 vssd1 vccd1 vccd1 _07915_/B
+ sky130_fd_sc_hd__o22a_1
X_08894_ _08895_/B vssd1 vssd1 vccd1 vccd1 _08894_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07845_ _07845_/A _07851_/A vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07776_ _07774_/X _07775_/X _07774_/X _07775_/X vssd1 vssd1 vccd1 vccd1 _07776_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06727_ _08752_/A vssd1 vssd1 vccd1 vccd1 _06727_/Y sky130_fd_sc_hd__inv_2
X_09515_ _09514_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09515_/X sky130_fd_sc_hd__mux2_1
X_09446_ _09424_/X _09445_/X _09424_/X _09445_/X vssd1 vssd1 vccd1 vccd1 _09446_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _10448_/Q vssd1 vssd1 vccd1 vccd1 _06658_/Y sky130_fd_sc_hd__inv_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06589_ _10109_/Q vssd1 vssd1 vccd1 vccd1 _08450_/A sky130_fd_sc_hd__inv_2
X_09377_ _09362_/X _09376_/X _09362_/X _09376_/X vssd1 vssd1 vccd1 vccd1 _09380_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_05609_ _05627_/A _05627_/B vssd1 vssd1 vccd1 vccd1 _05626_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08328_ _08328_/A vssd1 vssd1 vccd1 vccd1 _09982_/S sky130_fd_sc_hd__inv_16
X_08259_ _10195_/Q vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__inv_2
XFILLER_137_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10221_ _10300_/CLK _10221_/D vssd1 vssd1 vccd1 vccd1 _10221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10152_ _10329_/CLK _10152_/D vssd1 vssd1 vccd1 vccd1 _10152_/Q sky130_fd_sc_hd__dfxtp_1
X_10083_ _10176_/CLK _10083_/D vssd1 vssd1 vccd1 vccd1 _10083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10419_ _10422_/CLK _10419_/D vssd1 vssd1 vccd1 vccd1 _10419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05960_ _06111_/A vssd1 vssd1 vccd1 vccd1 _05960_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05891_ _06126_/A vssd1 vssd1 vccd1 vccd1 _05891_/X sky130_fd_sc_hd__clkbuf_4
X_07630_ _07582_/X _07629_/X _07582_/X _07629_/X vssd1 vssd1 vccd1 vccd1 _07630_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _07561_/A _07539_/X vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__or2b_1
X_06512_ _08411_/A _06489_/X _06516_/C _06508_/X vssd1 vssd1 vccd1 vccd1 _06512_/Y
+ sky130_fd_sc_hd__o22ai_1
X_09300_ _09300_/A _09470_/B _09173_/X vssd1 vssd1 vccd1 vccd1 _09300_/X sky130_fd_sc_hd__or3b_1
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07492_ _07663_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07493_/C sky130_fd_sc_hd__or2_1
XFILLER_194_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06443_ _06443_/A vssd1 vssd1 vccd1 vccd1 _06460_/A sky130_fd_sc_hd__clkbuf_2
X_09231_ _09983_/X vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__buf_2
XFILLER_194_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ _09162_/A _09162_/B vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__or2_1
X_06374_ _06372_/Y _06373_/X _06372_/Y _06373_/X vssd1 vssd1 vccd1 vccd1 _06374_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08113_ _10378_/Q _08312_/A _06714_/Y _06038_/X _08112_/X vssd1 vssd1 vccd1 vccd1
+ _08119_/C sky130_fd_sc_hd__o221a_1
XFILLER_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05325_ _05325_/A vssd1 vssd1 vccd1 vccd1 _05326_/B sky130_fd_sc_hd__inv_2
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _09190_/C _09092_/A _09245_/C _09092_/Y vssd1 vssd1 vccd1 vccd1 _09093_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05256_ input20/X _05251_/X _08763_/A _05252_/X _05253_/X vssd1 vssd1 vccd1 vccd1
+ _10357_/D sky130_fd_sc_hd__a221o_1
X_08044_ _08020_/A _08020_/B _08021_/B vssd1 vssd1 vccd1 vccd1 _08044_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05187_ _05185_/X _10394_/Q _05186_/X _09613_/X _05078_/X vssd1 vssd1 vccd1 vccd1
+ _10394_/D sky130_fd_sc_hd__o221a_1
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09995_ _08043_/X _07394_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__mux2_2
X_08946_ _08959_/A _08945_/B _08945_/X vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__a21bo_1
XFILLER_69_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08877_ _08882_/A vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07828_ _07828_/A _07864_/A vssd1 vssd1 vccd1 vccd1 _07829_/A sky130_fd_sc_hd__or2_2
X_07759_ _07707_/X _07758_/X _07707_/X _07758_/X vssd1 vssd1 vccd1 vccd1 _07760_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_197_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _09427_/X _09428_/X _09427_/X _09428_/X vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _10437_/CLK _10204_/D vssd1 vssd1 vccd1 vccd1 _10204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10135_ _10244_/CLK _10135_/D vssd1 vssd1 vccd1 vccd1 _10135_/Q sky130_fd_sc_hd__dfxtp_2
X_10066_ _10066_/CLK _10066_/D vssd1 vssd1 vccd1 vccd1 _10066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05110_ _10208_/Q vssd1 vssd1 vccd1 vccd1 _05369_/A sky130_fd_sc_hd__inv_2
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06090_ _10174_/Q _06088_/X _10346_/Q _06089_/X _05993_/X vssd1 vssd1 vccd1 vccd1
+ _10174_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05041_ input9/X input6/X input10/X vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__or3b_4
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08800_ _08772_/Y _08774_/X _08798_/Y _08820_/A vssd1 vssd1 vccd1 vccd1 _08800_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_112_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09780_ _09779_/X _08205_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__mux2_1
X_06992_ _06992_/A vssd1 vssd1 vccd1 vccd1 _06993_/B sky130_fd_sc_hd__buf_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08731_ _08731_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08731_/X sky130_fd_sc_hd__or2_1
XFILLER_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05943_ _10225_/Q vssd1 vssd1 vccd1 vccd1 _05943_/X sky130_fd_sc_hd__clkbuf_2
X_08662_ _08155_/X _10050_/Q _08569_/A _10051_/Q vssd1 vssd1 vccd1 vccd1 _08704_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _07667_/A _07613_/B vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__or2_1
X_05874_ _10255_/Q _05871_/X _05863_/X _06827_/A _05866_/X vssd1 vssd1 vccd1 vccd1
+ _10255_/D sky130_fd_sc_hd__o221a_1
X_08593_ _08593_/A _08593_/B _08593_/C vssd1 vssd1 vccd1 vccd1 _08593_/X sky130_fd_sc_hd__and3_1
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07544_ _07597_/A vssd1 vssd1 vccd1 vccd1 _07815_/A sky130_fd_sc_hd__buf_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07475_ _07676_/A vssd1 vssd1 vccd1 vccd1 _07766_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06426_ _06425_/A _06425_/B _06445_/A vssd1 vssd1 vccd1 vccd1 _06426_/X sky130_fd_sc_hd__o21a_1
X_09214_ _09119_/X _09126_/X _09127_/X _09156_/X vssd1 vssd1 vccd1 vccd1 _09214_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ _09045_/X _09144_/X _09045_/X _09144_/X vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06357_ _10242_/Q _08383_/A _06344_/A _06341_/X vssd1 vssd1 vccd1 vccd1 _06357_/X
+ sky130_fd_sc_hd__o22a_1
X_05308_ _10344_/Q _05317_/B vssd1 vssd1 vccd1 vccd1 _05309_/B sky130_fd_sc_hd__nand2_1
X_09076_ _09180_/C _09075_/A _09073_/A _09075_/Y vssd1 vssd1 vccd1 vccd1 _09076_/X
+ sky130_fd_sc_hd__a22o_1
X_06288_ _06288_/A vssd1 vssd1 vccd1 vccd1 _06288_/Y sky130_fd_sc_hd__inv_2
X_05239_ _05239_/A vssd1 vssd1 vccd1 vccd1 _05239_/X sky130_fd_sc_hd__clkbuf_2
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08027_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ _08905_/Y _08904_/B _09986_/S vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__mux2_2
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _08929_/A vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__inv_2
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10118_ _10244_/CLK _10118_/D vssd1 vssd1 vccd1 vccd1 _10118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10049_ _10447_/CLK _10049_/D vssd1 vssd1 vccd1 vccd1 _10049_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05590_ _09978_/X _05576_/X _05684_/A vssd1 vssd1 vccd1 vccd1 _05680_/B sky130_fd_sc_hd__o21ai_1
XFILLER_35_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07260_ _07093_/A _07093_/B _07094_/B vssd1 vssd1 vccd1 vccd1 _07260_/X sky130_fd_sc_hd__a21bo_1
XFILLER_191_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06211_ _06225_/A vssd1 vssd1 vccd1 vccd1 _06211_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _05964_/X _07126_/B _07108_/A _07189_/Y _07190_/X vssd1 vssd1 vccd1 vccd1
+ _07191_/X sky130_fd_sc_hd__a41o_1
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06142_ _09660_/X _06140_/X _10142_/Q _06141_/X _06135_/X vssd1 vssd1 vccd1 vccd1
+ _10142_/D sky130_fd_sc_hd__o221a_1
X_06073_ _09777_/X _06067_/X _06072_/X _06069_/X _06070_/X vssd1 vssd1 vccd1 vccd1
+ _10181_/D sky130_fd_sc_hd__o221a_1
X_05024_ _05024_/A vssd1 vssd1 vccd1 vccd1 _05024_/X sky130_fd_sc_hd__clkbuf_2
X_09901_ _09277_/X _09275_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09901_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09832_ _09831_/X _08262_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09763_ _10349_/Q _09762_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08714_ _08711_/A _08713_/B _06699_/Y _08713_/Y vssd1 vssd1 vccd1 vccd1 _08714_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06975_ _07235_/B _06992_/A vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__or2_2
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _06520_/Y input26/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09694_/X sky130_fd_sc_hd__mux2_1
X_05926_ _05928_/A vssd1 vssd1 vccd1 vccd1 _05927_/A sky130_fd_sc_hd__inv_2
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08645_ _08107_/X _10058_/Q _08104_/X _10057_/Q vssd1 vssd1 vccd1 vccd1 _08666_/A
+ sky130_fd_sc_hd__o22ai_2
X_05857_ _05793_/X _05822_/X _05793_/X _05822_/X vssd1 vssd1 vccd1 vccd1 _05858_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08576_ _08804_/A _08535_/B _08539_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _08595_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07527_ _07527_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__or2_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05788_ _05788_/A vssd1 vssd1 vccd1 vccd1 _05853_/A sky130_fd_sc_hd__inv_2
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07458_ _10279_/Q vssd1 vssd1 vccd1 vccd1 _07458_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06409_ _10248_/Q _08409_/A _06399_/X _06400_/X vssd1 vssd1 vccd1 vccd1 _06409_/Y
+ sky130_fd_sc_hd__o22ai_1
X_07389_ _07389_/A vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__inv_2
XFILLER_182_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09128_ _09128_/A vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_108_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09059_ _09007_/X _09013_/X _09014_/X _09015_/X vssd1 vssd1 vccd1 vccd1 _09060_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06760_ _10388_/Q _06792_/B vssd1 vssd1 vccd1 vccd1 _06760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06691_ _10378_/Q _06690_/A _06624_/Y _06690_/Y vssd1 vssd1 vccd1 vccd1 _06818_/B
+ sky130_fd_sc_hd__o22a_1
X_05711_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05711_/X sky130_fd_sc_hd__buf_1
X_08430_ _08430_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08430_/Y sky130_fd_sc_hd__nor2_1
X_05642_ _10309_/Q vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__inv_2
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _09354_/C vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__clkbuf_4
X_05573_ _09939_/X _05572_/X _09939_/X _05572_/X vssd1 vssd1 vccd1 vccd1 _05680_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_08292_ _06269_/A _06269_/B _08291_/Y vssd1 vssd1 vccd1 vccd1 _08292_/X sky130_fd_sc_hd__a21o_1
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ _06980_/X _06996_/X _06985_/A _07311_/Y vssd1 vssd1 vccd1 vccd1 _07312_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07243_ _07232_/A _07232_/B _07268_/A vssd1 vssd1 vccd1 vccd1 _07246_/A sky130_fd_sc_hd__a21o_1
XFILLER_176_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ _07173_/A _07173_/B _07180_/A vssd1 vssd1 vccd1 vccd1 _07177_/A sky130_fd_sc_hd__a21bo_1
XFILLER_191_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06125_ _10150_/Q _06117_/X _10322_/Q _06122_/X _06120_/X vssd1 vssd1 vccd1 vccd1
+ _10150_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06056_ _06069_/A vssd1 vssd1 vccd1 vccd1 _06056_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05007_ input17/X _05773_/C vssd1 vssd1 vccd1 vccd1 _06081_/A sky130_fd_sc_hd__or2_1
X_09815_ _10362_/Q _09814_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09815_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09746_ _10411_/Q _08059_/Y _09899_/S vssd1 vssd1 vccd1 vccd1 _09746_/X sky130_fd_sc_hd__mux2_1
X_06958_ _06958_/A _06958_/B vssd1 vssd1 vccd1 vccd1 _06958_/X sky130_fd_sc_hd__or2_1
X_09677_ _10158_/Q _10174_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__mux2_1
X_05909_ _10242_/Q _05902_/X input49/X _05903_/X _05908_/X vssd1 vssd1 vccd1 vccd1
+ _10242_/D sky130_fd_sc_hd__o221a_1
X_08628_ _08628_/A vssd1 vssd1 vccd1 vccd1 _08628_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06889_ _07112_/A _09892_/X vssd1 vssd1 vccd1 vccd1 _06889_/X sky130_fd_sc_hd__or2_1
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08077_/X _08557_/Y _08791_/A _08558_/B _08558_/Y vssd1 vssd1 vccd1 vccd1
+ _08559_/X sky130_fd_sc_hd__o221a_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10383_ _10422_/CLK _10383_/D vssd1 vssd1 vccd1 vccd1 _10383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07930_ _07761_/A _07761_/B _07906_/A vssd1 vssd1 vccd1 vccd1 _07930_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07861_ _07806_/X _07860_/X _07806_/X _07860_/X vssd1 vssd1 vccd1 vccd1 _07861_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_06812_ _06814_/A _06812_/B vssd1 vssd1 vccd1 vccd1 _06812_/Y sky130_fd_sc_hd__nor2_1
X_09600_ _08453_/Y _08452_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09600_/X sky130_fd_sc_hd__mux2_2
X_07792_ _07877_/A _07878_/D vssd1 vssd1 vccd1 vccd1 _07792_/X sky130_fd_sc_hd__or2_2
XFILLER_209_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _09530_/X _06635_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__mux2_2
X_06743_ _10380_/Q _06647_/A _10379_/Q _06623_/A vssd1 vssd1 vccd1 vccd1 _06743_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06674_ _10362_/Q _08745_/A vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__or2_4
X_09462_ _09474_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09462_/X sky130_fd_sc_hd__or3_1
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05625_ _05646_/A _05625_/B vssd1 vssd1 vccd1 vccd1 _10313_/D sky130_fd_sc_hd__nor2_1
X_09393_ _09393_/A _09393_/B vssd1 vssd1 vccd1 vccd1 _09393_/X sky130_fd_sc_hd__or2_1
X_08413_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__or2_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08344_ _09928_/X _08364_/B vssd1 vssd1 vccd1 vccd1 _08344_/Y sky130_fd_sc_hd__nor2_1
X_05556_ _05483_/X _05523_/X _05483_/X _05523_/X vssd1 vssd1 vccd1 vccd1 _05556_/X
+ sky130_fd_sc_hd__a2bb2o_2
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ _08275_/A vssd1 vssd1 vccd1 vccd1 _08275_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05487_ _09989_/X vssd1 vssd1 vccd1 vccd1 _05489_/A sky130_fd_sc_hd__inv_2
XFILLER_192_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07226_ _07211_/Y _07213_/Y _07224_/X _07225_/X vssd1 vssd1 vccd1 vccd1 _07226_/X
+ sky130_fd_sc_hd__o22a_1
X_07157_ _07145_/X _07146_/X _07145_/X _07146_/X vssd1 vssd1 vccd1 vccd1 _07157_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06108_ _10333_/Q _06088_/X _10161_/Q _06089_/X _05105_/A vssd1 vssd1 vccd1 vccd1
+ _10161_/D sky130_fd_sc_hd__a221o_1
XFILLER_105_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07088_ _07073_/A _07083_/Y _07080_/X _07084_/X vssd1 vssd1 vccd1 vccd1 _07095_/A
+ sky130_fd_sc_hd__o22ai_4
X_06039_ _09833_/X _06028_/X _06038_/X _06031_/X _06032_/X vssd1 vssd1 vccd1 vccd1
+ _10195_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _06800_/Y _10394_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10060_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ _10436_/CLK _10435_/D vssd1 vssd1 vccd1 vccd1 _10435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10436_/CLK _10366_/D vssd1 vssd1 vccd1 vccd1 _10366_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ _10297_/CLK _10297_/D vssd1 vssd1 vccd1 vccd1 _10297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05410_ _05404_/Y _05372_/X _05407_/Y _05395_/A _05409_/X vssd1 vssd1 vccd1 vccd1
+ _05411_/A sky130_fd_sc_hd__o32a_1
X_06390_ _06390_/A _10140_/Q vssd1 vssd1 vccd1 vccd1 _06391_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05341_ _05335_/B _05333_/X _05340_/Y _05336_/X _05303_/A vssd1 vssd1 vccd1 vccd1
+ _05342_/A sky130_fd_sc_hd__o32a_1
XFILLER_174_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05272_ _05032_/X _05263_/X _08625_/B _05264_/X _05265_/X vssd1 vssd1 vccd1 vccd1
+ _10349_/D sky130_fd_sc_hd__a221o_1
X_08060_ _08060_/A _08063_/B vssd1 vssd1 vccd1 vccd1 _08060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07011_ _07054_/A _07072_/B _07008_/A vssd1 vssd1 vccd1 vccd1 _07011_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _05939_/X _09418_/B _09001_/C _08961_/X vssd1 vssd1 vccd1 vccd1 _08962_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08893_ _08895_/A _08859_/X _08895_/A _08859_/X vssd1 vssd1 vccd1 vccd1 _08893_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07913_ _07913_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _07913_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07844_ _07829_/A _07839_/Y _07836_/X _07840_/X vssd1 vssd1 vccd1 vccd1 _07851_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07775_ _07425_/A _07777_/C _07766_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07775_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06726_ _10360_/Q _06672_/B _08748_/A vssd1 vssd1 vccd1 vccd1 _06798_/B sky130_fd_sc_hd__a21boi_4
X_09514_ _08401_/X _06377_/Y _09997_/S vssd1 vssd1 vccd1 vccd1 _09514_/X sky130_fd_sc_hd__mux2_1
X_09445_ _09142_/X _09225_/X _09251_/X _05922_/X _09444_/Y vssd1 vssd1 vccd1 vccd1
+ _09445_/X sky130_fd_sc_hd__o311a_1
X_06657_ _10349_/Q vssd1 vssd1 vccd1 vccd1 _06657_/Y sky130_fd_sc_hd__inv_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05608_ _09902_/X _05544_/X _05631_/A vssd1 vssd1 vccd1 vccd1 _05627_/B sky130_fd_sc_hd__o21ai_1
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06588_ _06591_/B _06587_/Y _06591_/B _06587_/Y vssd1 vssd1 vccd1 vccd1 _06588_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09376_ _09375_/A _09375_/B _09434_/A vssd1 vssd1 vccd1 vccd1 _09376_/X sky130_fd_sc_hd__a21bo_1
X_08327_ _08327_/A vssd1 vssd1 vccd1 vccd1 _09583_/S sky130_fd_sc_hd__clkbuf_4
X_05539_ _05472_/A _05472_/B _05472_/Y vssd1 vssd1 vccd1 vccd1 _05539_/Y sky130_fd_sc_hd__a21oi_2
X_08258_ _06038_/X _06261_/B _08257_/Y vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07209_ _07212_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07210_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08189_ _08657_/A _08186_/B _08191_/B _08188_/X vssd1 vssd1 vccd1 vccd1 _08189_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _10300_/CLK _10220_/D vssd1 vssd1 vccd1 vccd1 _10220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10329_/CLK _10151_/D vssd1 vssd1 vccd1 vccd1 _10151_/Q sky130_fd_sc_hd__dfxtp_1
X_10082_ _10450_/CLK _10082_/D vssd1 vssd1 vccd1 vccd1 _10082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10418_ _10422_/CLK _10418_/D vssd1 vssd1 vccd1 vccd1 _10418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _10414_/CLK _10349_/D vssd1 vssd1 vccd1 vccd1 _10349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05890_ _10251_/Q _05871_/X _05699_/X _06819_/B _05885_/X vssd1 vssd1 vccd1 vccd1
+ _10251_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07560_ _07603_/A _07539_/B _07813_/C _07634_/A vssd1 vssd1 vccd1 vccd1 _07561_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06511_ _08415_/A _06496_/A _10094_/Q _06461_/A vssd1 vssd1 vccd1 vccd1 _06516_/D
+ sky130_fd_sc_hd__a22o_1
X_09230_ _09230_/A _09229_/X vssd1 vssd1 vccd1 vccd1 _09238_/A sky130_fd_sc_hd__or2b_1
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07491_ _07663_/A _07537_/D vssd1 vssd1 vccd1 vccd1 _07498_/C sky130_fd_sc_hd__nor2_1
X_06442_ _06442_/A vssd1 vssd1 vccd1 vccd1 _06442_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ _09161_/A vssd1 vssd1 vccd1 vccd1 _09162_/B sky130_fd_sc_hd__inv_2
XFILLER_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06373_ _10244_/Q _08390_/A _06362_/A _06364_/Y vssd1 vssd1 vccd1 vccd1 _06373_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ _10375_/Q _08297_/A _06627_/Y _10204_/Q vssd1 vssd1 vccd1 vccd1 _08112_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09092_ _09092_/A vssd1 vssd1 vccd1 vccd1 _09092_/Y sky130_fd_sc_hd__inv_2
X_05324_ _05324_/A vssd1 vssd1 vccd1 vccd1 _10343_/D sky130_fd_sc_hd__inv_2
XFILLER_147_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ _07406_/A _07406_/B _07407_/B vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__a21bo_1
XFILLER_162_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05255_ _10357_/Q vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05186_ _05203_/A vssd1 vssd1 vccd1 vccd1 _05186_/X sky130_fd_sc_hd__clkbuf_2
X_09994_ _09385_/X _09383_/Y _09994_/S vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08945_ _08959_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08945_/X sky130_fd_sc_hd__or2_1
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08876_ _05581_/X _07921_/A _08857_/X _08858_/Y vssd1 vssd1 vccd1 vccd1 _08876_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07827_ _07812_/X _07813_/X _07825_/X _07826_/X vssd1 vssd1 vccd1 vccd1 _07827_/X
+ sky130_fd_sc_hd__o22a_1
X_07758_ _07523_/A _07529_/A _07523_/Y vssd1 vssd1 vccd1 vccd1 _07758_/X sky130_fd_sc_hd__a21o_1
X_06709_ _10369_/Q _08724_/A _06707_/Y vssd1 vssd1 vccd1 vccd1 _06808_/B sky130_fd_sc_hd__a21oi_2
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07689_ _07680_/B _07688_/A _07679_/A _07688_/Y vssd1 vssd1 vccd1 vccd1 _07689_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09474_/A _09462_/B _09428_/C vssd1 vssd1 vccd1 vccd1 _09428_/X sky130_fd_sc_hd__or3_4
X_09359_ _09359_/A _09359_/B vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__or2_1
XFILLER_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _10437_/CLK _10203_/D vssd1 vssd1 vccd1 vccd1 _10203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10134_ _10244_/CLK _10134_/D vssd1 vssd1 vccd1 vccd1 _10134_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _10066_/CLK _10065_/D vssd1 vssd1 vccd1 vccd1 _10065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05040_ _06184_/A vssd1 vssd1 vccd1 vccd1 _05968_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06991_ _07234_/B _07047_/D vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__nand2_4
X_08730_ _06633_/A _08729_/X _08727_/Y vssd1 vssd1 vccd1 vccd1 _08730_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05942_ _05941_/X _05927_/A input19/X _05928_/A _05934_/X vssd1 vssd1 vccd1 vccd1
+ _10226_/D sky130_fd_sc_hd__o221a_1
XFILLER_85_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08661_ _08138_/X _10049_/Q _08116_/X _08456_/X _08660_/X vssd1 vssd1 vccd1 vccd1
+ _08661_/Y sky130_fd_sc_hd__a221oi_2
X_05873_ _05873_/A vssd1 vssd1 vccd1 vccd1 _06827_/A sky130_fd_sc_hd__inv_2
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07612_ _07612_/A vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__buf_2
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08592_ _08592_/A _08592_/B _08592_/C _08537_/X vssd1 vssd1 vccd1 vccd1 _08594_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07543_ _07540_/X _07542_/X _07540_/X _07542_/X vssd1 vssd1 vccd1 vccd1 _07550_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07474_ _07676_/A _07504_/B _07806_/A _07558_/B vssd1 vssd1 vccd1 vccd1 _07477_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ _09178_/X _09212_/X _09178_/X _09212_/X vssd1 vssd1 vccd1 vccd1 _09213_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06425_ _06425_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06445_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ _09170_/A _09142_/X _09190_/C _09143_/X vssd1 vssd1 vccd1 vccd1 _09144_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_135_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06356_ _06353_/Y _06355_/A _06353_/A _06355_/Y vssd1 vssd1 vccd1 vccd1 _06356_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _09075_/A vssd1 vssd1 vccd1 vccd1 _09075_/Y sky130_fd_sc_hd__inv_2
X_05307_ _05307_/A _05319_/A vssd1 vssd1 vccd1 vccd1 _05317_/B sky130_fd_sc_hd__nor2_4
X_06287_ _10235_/Q _08335_/A _05771_/C _06277_/Y vssd1 vssd1 vccd1 vccd1 _06288_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05238_ _10366_/Q _05230_/X input29/X _05231_/X _05236_/X vssd1 vssd1 vccd1 vccd1
+ _10366_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08026_ _08026_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__or2_2
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05169_ _10430_/Q vssd1 vssd1 vccd1 vccd1 _05169_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09977_ _08910_/Y _08907_/X _09986_/S vssd1 vssd1 vccd1 vccd1 _09977_/X sky130_fd_sc_hd__mux2_2
XFILLER_162_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08928_ _08853_/X _08861_/X _08853_/X _08861_/X vssd1 vssd1 vccd1 vccd1 _08929_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ _10284_/Q _07423_/Y _08858_/Y vssd1 vssd1 vccd1 vccd1 _08859_/X sky130_fd_sc_hd__o21ba_1
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10117_ _10334_/CLK _10117_/D vssd1 vssd1 vccd1 vccd1 _10117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10048_ _10450_/CLK _10048_/D vssd1 vssd1 vccd1 vccd1 _10048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06210_ _06224_/A vssd1 vssd1 vccd1 vccd1 _06210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07190_ _06887_/A _07102_/B _07112_/A _07189_/A vssd1 vssd1 vccd1 vccd1 _07190_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_129_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06141_ _06157_/A vssd1 vssd1 vccd1 vccd1 _06141_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06072_ _10181_/Q vssd1 vssd1 vccd1 vccd1 _06072_/X sky130_fd_sc_hd__buf_2
X_05023_ _10448_/Q vssd1 vssd1 vccd1 vccd1 _05024_/A sky130_fd_sc_hd__buf_1
X_09900_ _09163_/X _09161_/A _09994_/S vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__mux2_2
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09831_ _10366_/Q _09830_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ _08185_/Y _10349_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06974_ _06977_/A _07218_/B vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__or2_2
X_08713_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08713_/Y sky130_fd_sc_hd__nor2_1
X_05925_ _05968_/A _08316_/A vssd1 vssd1 vccd1 vccd1 _05928_/A sky130_fd_sc_hd__or2_4
X_09693_ _06513_/X input25/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _08166_/X _10059_/Q _06047_/X _08643_/Y vssd1 vssd1 vccd1 vccd1 _08644_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05856_ _10260_/Q _05851_/X _05842_/X _06836_/A _05845_/X vssd1 vssd1 vccd1 vccd1
+ _10260_/D sky130_fd_sc_hd__o221a_1
X_08575_ _08592_/C _08572_/Y _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08575_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05787_ _07437_/A _10261_/Q vssd1 vssd1 vccd1 vccd1 _05787_/Y sky130_fd_sc_hd__nor2_1
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07498_/C _07494_/B _07494_/Y vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__o21ai_1
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _05704_/X _07455_/B _07854_/B vssd1 vssd1 vccd1 vccd1 _07457_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06408_ _06404_/X _06407_/X _06404_/X _06407_/X vssd1 vssd1 vccd1 vccd1 _06408_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_07388_ _07388_/A vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__inv_2
XFILLER_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _09119_/X _09126_/X _09119_/X _09126_/X vssd1 vssd1 vccd1 vccd1 _09127_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06339_ _06337_/Y _10135_/Q _10242_/Q _08383_/A vssd1 vssd1 vccd1 vccd1 _06344_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09058_ _09057_/A _09057_/B _09057_/Y vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__a21o_1
XFILLER_135_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08009_ _08009_/A vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__inv_2
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 _10026_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_209_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06690_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06690_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05710_ _07437_/A vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__clkbuf_2
X_05641_ _05641_/A _05641_/B vssd1 vssd1 vccd1 vccd1 _05641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08360_ _09252_/A vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07311_ _07311_/A _07311_/B vssd1 vssd1 vccd1 vccd1 _07311_/Y sky130_fd_sc_hd__nor2_1
X_05572_ _05570_/Y _05571_/Y _05570_/Y _05571_/Y vssd1 vssd1 vccd1 vccd1 _05572_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_08291_ _08291_/A vssd1 vssd1 vccd1 vccd1 _08291_/Y sky130_fd_sc_hd__inv_2
X_07242_ _07242_/A vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__inv_2
X_07173_ _07173_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _07180_/A sky130_fd_sc_hd__or2_1
XFILLER_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06124_ _10151_/Q _06117_/X _10323_/Q _06122_/X _06120_/X vssd1 vssd1 vccd1 vccd1
+ _10151_/D sky130_fd_sc_hd__o221a_1
XFILLER_172_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06055_ _10187_/Q vssd1 vssd1 vccd1 vccd1 _06253_/A sky130_fd_sc_hd__buf_2
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05006_ input8/X input7/X vssd1 vssd1 vccd1 vccd1 _05773_/C sky130_fd_sc_hd__or2_2
X_09814_ _08239_/X _10362_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09814_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09745_ _06818_/Y _10410_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10076_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06957_ _06935_/X _06955_/X _06878_/X _06956_/X vssd1 vssd1 vccd1 vccd1 _06958_/B
+ sky130_fd_sc_hd__o22a_1
X_09676_ _10157_/Q _10173_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09676_/X sky130_fd_sc_hd__mux2_1
X_05908_ _05934_/A vssd1 vssd1 vccd1 vccd1 _05908_/X sky130_fd_sc_hd__buf_1
X_06888_ _06931_/A _09891_/X vssd1 vssd1 vccd1 vccd1 _06888_/X sky130_fd_sc_hd__or2_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ _05024_/X _08146_/Y _06658_/Y _05273_/X vssd1 vssd1 vccd1 vccd1 _08628_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05839_ _08842_/B _10263_/Q _05785_/Y vssd1 vssd1 vccd1 vccd1 _05839_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08791_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08489_ _10071_/Q _08489_/B vssd1 vssd1 vccd1 vccd1 _08490_/B sky130_fd_sc_hd__or2_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07509_ _07509_/A vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_210_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _10414_/CLK _10382_/D vssd1 vssd1 vccd1 vccd1 _10382_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _07807_/X _07859_/X _07807_/X _07859_/X vssd1 vssd1 vccd1 vccd1 _07860_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06811_ _06814_/A _06811_/B vssd1 vssd1 vccd1 vccd1 _06811_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07791_ _10212_/Q _07788_/Y _07854_/D _07789_/Y _07790_/X vssd1 vssd1 vccd1 vccd1
+ _07794_/A sky130_fd_sc_hd__a41o_1
XFILLER_209_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09530_ _05176_/Y _08125_/X _09981_/S vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__mux2_1
X_06742_ _06742_/A vssd1 vssd1 vccd1 vccd1 _06742_/Y sky130_fd_sc_hd__inv_2
X_09461_ _09450_/X _09460_/X _09450_/X _09460_/X vssd1 vssd1 vccd1 vccd1 _09461_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06673_ _10361_/Q _08748_/A vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__or2_2
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08412_ _09501_/X _08419_/B vssd1 vssd1 vccd1 vccd1 _08412_/Y sky130_fd_sc_hd__nor2_2
X_05624_ _05619_/X _05620_/Y _05621_/Y _08075_/A _05623_/X vssd1 vssd1 vccd1 vccd1
+ _05625_/B sky130_fd_sc_hd__o32a_1
X_09392_ _09392_/A vssd1 vssd1 vccd1 vccd1 _09392_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05555_ _09900_/X _05554_/X _09900_/X _05554_/X vssd1 vssd1 vccd1 vccd1 _05649_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_08343_ _08343_/A _09748_/S vssd1 vssd1 vccd1 vccd1 _08343_/X sky130_fd_sc_hd__or2_1
XFILLER_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08274_ _06026_/X _08270_/Y _08264_/X _08277_/B vssd1 vssd1 vccd1 vccd1 _08274_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07225_ _07211_/Y _07213_/Y _07211_/Y _07213_/Y vssd1 vssd1 vccd1 vccd1 _07225_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05486_ _05486_/A _05486_/B vssd1 vssd1 vccd1 vccd1 _05486_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07156_ _07147_/X _07148_/X _07154_/X _07155_/X vssd1 vssd1 vccd1 vccd1 _07156_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06107_ _10334_/Q _06101_/X _10162_/Q _06102_/X _05105_/A vssd1 vssd1 vccd1 vccd1
+ _10162_/D sky130_fd_sc_hd__a221o_1
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07087_ _07087_/A vssd1 vssd1 vccd1 vccd1 _07089_/A sky130_fd_sc_hd__inv_2
X_06038_ _08733_/A vssd1 vssd1 vccd1 vccd1 _06038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09728_ _06799_/Y _10393_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10059_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07989_ _07966_/X _07971_/X _07966_/X _07971_/X vssd1 vssd1 vccd1 vccd1 _08006_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _10125_/Q input24/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10434_ _10436_/CLK _10434_/D vssd1 vssd1 vccd1 vccd1 _10434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10365_ _10436_/CLK _10365_/D vssd1 vssd1 vccd1 vccd1 _10365_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10296_ _10297_/CLK _10296_/D vssd1 vssd1 vccd1 vccd1 _10296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05340_ _10339_/Q _05340_/B vssd1 vssd1 vccd1 vccd1 _05340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05271_ _10349_/Q vssd1 vssd1 vccd1 vccd1 _08625_/B sky130_fd_sc_hd__buf_2
XFILLER_162_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ _07116_/B vssd1 vssd1 vccd1 vccd1 _07072_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _09069_/A _09128_/A _09029_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _08961_/X
+ sky130_fd_sc_hd__o22a_1
X_08892_ _08899_/C _08890_/X _08903_/A vssd1 vssd1 vccd1 vccd1 _08892_/Y sky130_fd_sc_hd__o21ai_1
X_07912_ _07909_/X _07911_/Y _07909_/X _07911_/Y vssd1 vssd1 vccd1 vccd1 _07912_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07843_ _07843_/A vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__inv_2
XFILLER_204_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07774_ _07921_/B _07916_/C _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07774_/X
+ sky130_fd_sc_hd__o22a_1
X_06725_ _10361_/Q _08748_/A _06723_/Y vssd1 vssd1 vccd1 vccd1 _06799_/B sky130_fd_sc_hd__a21oi_4
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _09512_/X _07777_/A _10000_/S vssd1 vssd1 vccd1 vccd1 _09513_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09142_/X _09225_/X _09251_/X vssd1 vssd1 vccd1 vccd1 _09444_/Y sky130_fd_sc_hd__o21ai_1
X_06656_ _08625_/A _10350_/Q vssd1 vssd1 vccd1 vccd1 _06656_/Y sky130_fd_sc_hd__nor2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05607_ _05632_/A _05632_/B vssd1 vssd1 vccd1 vccd1 _05631_/A sky130_fd_sc_hd__or2_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06587_ _08446_/A _06489_/X _06591_/A vssd1 vssd1 vccd1 vccd1 _06587_/Y sky130_fd_sc_hd__o21ai_1
X_09375_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__or2_1
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08326_ _08380_/A _09582_/S _08452_/B vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__or3b_2
X_05538_ _05538_/A vssd1 vssd1 vccd1 vccd1 _05538_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08257_/Y sky130_fd_sc_hd__inv_2
X_05469_ _10018_/X _10006_/X _10018_/X _10006_/X vssd1 vssd1 vccd1 vccd1 _05469_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_192_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08188_ _08264_/A vssd1 vssd1 vccd1 vccd1 _08188_/X sky130_fd_sc_hd__buf_2
XFILLER_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07208_ _07119_/X _07140_/X _07141_/X _07206_/X _07207_/X vssd1 vssd1 vccd1 vccd1
+ _07208_/X sky130_fd_sc_hd__o221a_1
XFILLER_192_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07139_ _07139_/A _07202_/B vssd1 vssd1 vccd1 vccd1 _07139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_160_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _10329_/CLK _10150_/D vssd1 vssd1 vccd1 vccd1 _10150_/Q sky130_fd_sc_hd__dfxtp_1
X_10081_ _10450_/CLK _10081_/D vssd1 vssd1 vccd1 vccd1 _10081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ _10422_/CLK _10417_/D vssd1 vssd1 vccd1 vccd1 _10417_/Q sky130_fd_sc_hd__dfxtp_1
X_10348_ _10442_/CLK _10348_/D vssd1 vssd1 vccd1 vccd1 _10348_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10279_ _10298_/CLK _10279_/D vssd1 vssd1 vccd1 vccd1 _10279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06510_ _10094_/Q vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__inv_2
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07490_ _09934_/X vssd1 vssd1 vccd1 vccd1 _07539_/B sky130_fd_sc_hd__clkbuf_2
X_06441_ _10083_/Q vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__inv_2
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ _09159_/A _09159_/B _09159_/X vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__a21bo_1
X_06372_ _06372_/A vssd1 vssd1 vccd1 vccd1 _06372_/Y sky130_fd_sc_hd__inv_2
X_08111_ _10204_/Q vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__inv_2
XFILLER_159_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09091_ _10233_/Q _09168_/A _09091_/C vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__and3_1
XFILLER_119_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05323_ _05317_/B _05282_/X _05320_/Y _05322_/X _05307_/A vssd1 vssd1 vccd1 vccd1
+ _05324_/A sky130_fd_sc_hd__o32a_1
X_05254_ input21/X _05251_/X _10358_/Q _05252_/X _05253_/X vssd1 vssd1 vccd1 vccd1
+ _10358_/D sky130_fd_sc_hd__a221o_1
X_08042_ _08021_/A _08021_/B _08022_/B vssd1 vssd1 vccd1 vccd1 _08042_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05185_ _05193_/A vssd1 vssd1 vccd1 vccd1 _05185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09993_ _07997_/Y _08052_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08944_ _08943_/A _08943_/B _08943_/Y vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__a21o_1
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08875_ _08872_/X _08874_/X _08872_/X _08874_/X vssd1 vssd1 vccd1 vccd1 _09986_/S
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07826_ _07812_/X _07813_/X _07812_/X _07813_/X vssd1 vssd1 vccd1 vccd1 _07826_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07757_ _07705_/X _07708_/X _07709_/X _07756_/X vssd1 vssd1 vccd1 vccd1 _07760_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06708_ _06706_/Y _06707_/Y _08719_/A vssd1 vssd1 vccd1 vccd1 _06710_/A sky130_fd_sc_hd__o21ai_2
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07688_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07688_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09427_ _09260_/A _09367_/A _09368_/X _09369_/X vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o22a_1
X_06639_ _10392_/Q vssd1 vssd1 vccd1 vccd1 _06639_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09358_ _09291_/X _09305_/X _09288_/X _09306_/X vssd1 vssd1 vccd1 vccd1 _09359_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ _08309_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08313_/A sky130_fd_sc_hd__or2_2
XFILLER_100_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09289_ _09289_/A vssd1 vssd1 vccd1 vccd1 _09457_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ _10202_/CLK _10202_/D vssd1 vssd1 vccd1 vccd1 _10202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10133_ _10244_/CLK _10133_/D vssd1 vssd1 vccd1 vccd1 _10133_/Q sky130_fd_sc_hd__dfxtp_1
X_10064_ _10399_/CLK _10064_/D vssd1 vssd1 vccd1 vccd1 _10064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06990_ _06986_/X _06989_/X _06986_/X _06989_/X vssd1 vssd1 vccd1 vccd1 _06990_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05941_ _10226_/Q vssd1 vssd1 vccd1 vccd1 _05941_/X sky130_fd_sc_hd__buf_2
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08660_ _08130_/X _10046_/Q _08657_/Y _08658_/X _08704_/C vssd1 vssd1 vccd1 vccd1
+ _08660_/X sky130_fd_sc_hd__o311a_1
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05872_ _05807_/X _05818_/X _05807_/X _05818_/X vssd1 vssd1 vccd1 vccd1 _05873_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07611_ _07596_/X _07597_/X _07596_/X _07597_/X vssd1 vssd1 vccd1 vccd1 _07611_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_08591_ _08591_/A _08591_/B _08591_/C _08547_/X vssd1 vssd1 vccd1 vccd1 _08592_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_19_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ _07597_/A _09935_/X vssd1 vssd1 vccd1 vccd1 _07542_/X sky130_fd_sc_hd__or2_1
XFILLER_61_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07473_ _07552_/B vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_179_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ _09210_/X _09211_/X _09210_/X _09211_/X vssd1 vssd1 vccd1 vccd1 _09212_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06424_ _10080_/Q _06443_/A _10079_/Q _06418_/X vssd1 vssd1 vccd1 vccd1 _06425_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09143_ _09258_/A _09089_/B _09259_/A _09096_/A vssd1 vssd1 vccd1 vccd1 _09143_/X
+ sky130_fd_sc_hd__o22a_1
X_06355_ _06355_/A vssd1 vssd1 vccd1 vccd1 _06355_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05306_ _05306_/A _05325_/A vssd1 vssd1 vccd1 vccd1 _05319_/A sky130_fd_sc_hd__or2_2
X_09074_ _09294_/A _09418_/B _09074_/C vssd1 vssd1 vccd1 vccd1 _09075_/A sky130_fd_sc_hd__and3_1
X_06286_ _06285_/A _06285_/B _06285_/X vssd1 vssd1 vccd1 vccd1 _06286_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05237_ _06633_/A _05230_/X input31/X _05231_/X _05236_/X vssd1 vssd1 vccd1 vccd1
+ _10367_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08025_ _08025_/A _08025_/B vssd1 vssd1 vccd1 vccd1 _08026_/B sky130_fd_sc_hd__or2_1
X_05168_ _10398_/Q vssd1 vssd1 vccd1 vccd1 _05168_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09976_ _09068_/X _09066_/A _09986_/S vssd1 vssd1 vccd1 vccd1 _09976_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05099_ _05030_/X _05094_/X _10414_/Q _05095_/X _05097_/X vssd1 vssd1 vccd1 vccd1
+ _10414_/D sky130_fd_sc_hd__a221o_1
X_08927_ _08926_/A _08926_/B _08950_/A vssd1 vssd1 vccd1 vccd1 _08927_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08858_ _05581_/X _07686_/A _08857_/X vssd1 vssd1 vccd1 vccd1 _08858_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07809_ _09917_/X vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__clkbuf_2
X_08789_ _06603_/X _06621_/A _08626_/Y vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__a21oi_2
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ _10334_/CLK _10116_/D vssd1 vssd1 vccd1 vccd1 _10116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10047_ _10450_/CLK _10047_/D vssd1 vssd1 vccd1 vccd1 _10047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06140_ _06156_/A vssd1 vssd1 vccd1 vccd1 _06140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06071_ _09781_/X _06067_/X _08797_/A _06069_/X _06070_/X vssd1 vssd1 vccd1 vccd1
+ _10182_/D sky130_fd_sc_hd__o221a_1
X_05022_ _05013_/X _05017_/Y _05018_/X _09940_/S _06182_/A vssd1 vssd1 vccd1 vccd1
+ _10449_/D sky130_fd_sc_hd__o221a_1
XFILLER_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09830_ _08258_/X _10366_/Q _09874_/S vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _09760_/X input30/X _09801_/S vssd1 vssd1 vccd1 vccd1 _09761_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06973_ _07212_/B vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__buf_2
X_08712_ _08709_/A _08713_/B _06627_/Y _08711_/Y vssd1 vssd1 vccd1 vccd1 _08712_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05924_ _06082_/B _06137_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__or2_4
X_09692_ _06509_/Y input24/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08643_ _10060_/Q vssd1 vssd1 vccd1 vccd1 _08643_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05855_ _05823_/Y _05854_/Y _05853_/Y _05824_/Y vssd1 vssd1 vccd1 vccd1 _06836_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08574_ _08765_/A _08574_/B vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__nand2_1
X_05786_ _05786_/A _10262_/Q vssd1 vssd1 vccd1 vccd1 _05786_/Y sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ _07513_/A _07513_/B _07706_/A vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__a21o_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07456_ _07456_/A vssd1 vssd1 vccd1 vccd1 _07854_/B sky130_fd_sc_hd__inv_2
X_06407_ _10249_/Q _10142_/Q _06405_/Y _08413_/A vssd1 vssd1 vccd1 vccd1 _06407_/X
+ sky130_fd_sc_hd__o22a_1
X_07387_ _07387_/A vssd1 vssd1 vccd1 vccd1 _07412_/A sky130_fd_sc_hd__inv_2
XFILLER_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _05939_/X _09294_/B _09174_/C _09125_/X vssd1 vssd1 vccd1 vccd1 _09126_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06338_ _10135_/Q vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__inv_2
X_06269_ _06269_/A _06269_/B vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__or2_1
XFILLER_163_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _09057_/Y sky130_fd_sc_hd__nor2_4
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _08008_/A vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__inv_2
XFILLER_190_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _09958_/X _06627_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput70 _09589_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput81 _09599_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05640_ _05640_/A vssd1 vssd1 vccd1 vccd1 _05640_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05571_ _05494_/A _05494_/B _05494_/Y vssd1 vssd1 vccd1 vccd1 _05571_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07310_ _07052_/Y _07309_/X _07052_/Y _07309_/X vssd1 vssd1 vccd1 vccd1 _07310_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08290_ _06268_/A _08286_/Y _08264_/X _08294_/B vssd1 vssd1 vccd1 vccd1 _08290_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07241_ _07241_/A _07247_/A vssd1 vssd1 vccd1 vccd1 _07241_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07172_ _07154_/A _07154_/B _07154_/X vssd1 vssd1 vccd1 vccd1 _07173_/B sky130_fd_sc_hd__a21bo_1
XFILLER_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06123_ _10152_/Q _06117_/X _10324_/Q _06122_/X _06120_/X vssd1 vssd1 vccd1 vccd1
+ _10152_/D sky130_fd_sc_hd__o221a_1
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06054_ _06067_/A vssd1 vssd1 vccd1 vccd1 _06054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05005_ input18/X vssd1 vssd1 vccd1 vccd1 _06081_/B sky130_fd_sc_hd__inv_2
X_09813_ _09812_/X input24/X _09821_/S vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ _06817_/Y _10409_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10075_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06956_ _06935_/X _06955_/X _06935_/X _06955_/X vssd1 vssd1 vccd1 vccd1 _06956_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09675_ _10156_/Q _10172_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__mux2_1
X_05907_ _10243_/Q _05902_/X input50/X _05903_/X _05900_/X vssd1 vssd1 vccd1 vccd1
+ _10243_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06887_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06931_/A sky130_fd_sc_hd__clkbuf_2
X_08626_ _08626_/A _10347_/Q vssd1 vssd1 vccd1 vccd1 _08626_/Y sky130_fd_sc_hd__nor2_2
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05838_ _10264_/Q _05780_/X _05637_/X _07023_/A _05764_/X vssd1 vssd1 vccd1 vccd1
+ _10264_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08557_/A vssd1 vssd1 vccd1 vccd1 _08557_/Y sky130_fd_sc_hd__inv_2
X_05769_ _10234_/Q vssd1 vssd1 vccd1 vccd1 _05770_/A sky130_fd_sc_hd__inv_2
X_08488_ _10070_/Q _08488_/B vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__or2_1
XFILLER_195_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07508_ _07566_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_210_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ _10276_/Q _07439_/B vssd1 vssd1 vccd1 vccd1 _07440_/B sky130_fd_sc_hd__or2_1
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ _10450_/CLK _10450_/D vssd1 vssd1 vccd1 vccd1 _10450_/Q sky130_fd_sc_hd__dfxtp_1
X_09109_ _09122_/A _09108_/Y _09122_/A _09108_/Y vssd1 vssd1 vccd1 vccd1 _09109_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10381_ _10422_/CLK _10381_/D vssd1 vssd1 vccd1 vccd1 _10381_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_190_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06810_ _06814_/A _06810_/B vssd1 vssd1 vccd1 vccd1 _06810_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _07828_/A _09904_/X _07877_/A _09908_/X vssd1 vssd1 vccd1 vccd1 _07790_/X
+ sky130_fd_sc_hd__o22a_1
X_06741_ _08626_/A _05273_/X _06660_/A _06645_/Y _06660_/Y vssd1 vssd1 vccd1 vccd1
+ _06742_/A sky130_fd_sc_hd__o32a_1
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09460_ _09340_/X _09459_/Y _09340_/X _09459_/Y vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06672_ _10360_/Q _06672_/B vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__or2_4
X_08411_ _08411_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08411_/Y sky130_fd_sc_hd__nor2_1
X_09391_ _09389_/X _09390_/X _09389_/X _09390_/X vssd1 vssd1 vccd1 vccd1 _09391_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05623_ _05750_/A vssd1 vssd1 vccd1 vccd1 _05623_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08342_ _09292_/A vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__clkbuf_4
X_05554_ _05482_/X _05524_/X _05482_/X _05524_/X vssd1 vssd1 vccd1 vccd1 _05554_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_08273_ _08273_/A _08273_/B vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__or2_1
XFILLER_149_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05485_ _09995_/X vssd1 vssd1 vccd1 vccd1 _05486_/B sky130_fd_sc_hd__inv_2
XFILLER_177_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07224_ _07214_/X _07215_/X _07222_/X _07223_/X vssd1 vssd1 vccd1 vccd1 _07224_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ _07155_/A _09884_/X _07155_/C vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__or3_1
X_06106_ _10335_/Q _06101_/X _10163_/Q _06102_/X _06099_/X vssd1 vssd1 vccd1 vccd1
+ _10163_/D sky130_fd_sc_hd__a221o_1
X_07086_ _07069_/X _07070_/X _07069_/X _07070_/X vssd1 vssd1 vccd1 vccd1 _07087_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06037_ _10195_/Q vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07988_ _07959_/X _07972_/X _07959_/X _07972_/X vssd1 vssd1 vccd1 vccd1 _08005_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ _06798_/Y _10392_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10058_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06939_ _06927_/X _06938_/X _06927_/X _06938_/X vssd1 vssd1 vccd1 vccd1 _06939_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _10124_/Q input23/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08609_ _10205_/Q _08496_/Y _08608_/X vssd1 vssd1 vccd1 vccd1 _08609_/Y sky130_fd_sc_hd__a21boi_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _08428_/Y _08427_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09589_/X sky130_fd_sc_hd__mux2_2
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10433_ _10433_/CLK _10433_/D vssd1 vssd1 vccd1 vccd1 _10433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10364_ _10436_/CLK _10364_/D vssd1 vssd1 vccd1 vccd1 _10364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10295_ _10297_/CLK _10295_/D vssd1 vssd1 vccd1 vccd1 _10295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05270_ _05030_/X _05263_/X _08624_/B _05264_/X _05265_/X vssd1 vssd1 vccd1 vccd1
+ _10350_/D sky130_fd_sc_hd__a221o_1
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08960_ _09986_/X vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08891_ _08899_/C _08891_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _07913_/B vssd1 vssd1 vccd1 vccd1 _07911_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07842_ _07825_/X _07826_/X _07825_/X _07826_/X vssd1 vssd1 vccd1 vccd1 _07843_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09512_ _09511_/X _07054_/A _09999_/S vssd1 vssd1 vccd1 vccd1 _09512_/X sky130_fd_sc_hd__mux2_1
X_07773_ _07773_/A vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__inv_2
X_06724_ _06722_/Y _06723_/Y _08742_/A vssd1 vssd1 vccd1 vccd1 _06800_/B sky130_fd_sc_hd__o21a_1
X_09443_ _09442_/A _09442_/B _09442_/X vssd1 vssd1 vccd1 vccd1 _09443_/X sky130_fd_sc_hd__a21bo_1
X_06655_ _08459_/A vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__clkbuf_2
X_09374_ _09321_/A _09321_/B _09373_/Y _09321_/Y _09373_/A vssd1 vssd1 vccd1 vccd1
+ _09375_/B sky130_fd_sc_hd__a32o_1
X_05606_ _09901_/X _05548_/X _05549_/X _05605_/X vssd1 vssd1 vccd1 vccd1 _05632_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06586_ _10108_/Q _06466_/A _08448_/A _06437_/A vssd1 vssd1 vccd1 vccd1 _06591_/B
+ sky130_fd_sc_hd__a22o_1
X_08325_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08452_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05537_ _09907_/X _05536_/X _09907_/X _05536_/X vssd1 vssd1 vccd1 vccd1 _05621_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_08256_ _06260_/A _08250_/Y _08219_/X _08260_/B vssd1 vssd1 vccd1 vccd1 _08256_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_177_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05468_ _05468_/A vssd1 vssd1 vccd1 vccd1 _05468_/X sky130_fd_sc_hd__buf_2
X_08187_ _08240_/A vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__inv_2
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07207_ _07099_/A _07100_/X _07115_/X _07118_/X vssd1 vssd1 vccd1 vccd1 _07207_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05399_ _05399_/A vssd1 vssd1 vccd1 vccd1 _05718_/A sky130_fd_sc_hd__buf_2
X_07138_ _07138_/A _07138_/B vssd1 vssd1 vccd1 vccd1 _07202_/B sky130_fd_sc_hd__nor2_2
XFILLER_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07069_ _07058_/X _07059_/X _07067_/X _07068_/X vssd1 vssd1 vccd1 vccd1 _07069_/X
+ sky130_fd_sc_hd__o22a_1
X_10080_ _10176_/CLK _10080_/D vssd1 vssd1 vccd1 vccd1 _10080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_0 _07806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10416_ _10422_/CLK _10416_/D vssd1 vssd1 vccd1 vccd1 _10416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10347_ _10442_/CLK _10347_/D vssd1 vssd1 vccd1 vccd1 _10347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10278_ _10298_/CLK _10278_/D vssd1 vssd1 vccd1 vccd1 _10278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06440_ _06445_/B _06439_/Y _06445_/B _06439_/Y vssd1 vssd1 vccd1 vccd1 _06440_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06371_ _06370_/A _10138_/Q _06370_/Y vssd1 vssd1 vccd1 vccd1 _06372_/A sky130_fd_sc_hd__a21oi_2
X_08110_ _10207_/Q vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__inv_2
X_09090_ _09245_/C vssd1 vssd1 vccd1 vccd1 _09190_/C sky130_fd_sc_hd__inv_2
X_05322_ _05336_/A vssd1 vssd1 vccd1 vccd1 _05322_/X sky130_fd_sc_hd__buf_2
XFILLER_119_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05253_ _05274_/A vssd1 vssd1 vccd1 vccd1 _05253_/X sky130_fd_sc_hd__buf_1
X_08041_ _07407_/A _07407_/B _07408_/B vssd1 vssd1 vccd1 vccd1 _08041_/X sky130_fd_sc_hd__a21bo_1
X_05184_ _05646_/A _05184_/B vssd1 vssd1 vccd1 vccd1 _10395_/D sky130_fd_sc_hd__nor2_1
XFILLER_127_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _08008_/A _08042_/X _10282_/Q vssd1 vssd1 vccd1 vccd1 _09992_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _08943_/A _08943_/B vssd1 vssd1 vccd1 vccd1 _08943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08874_ _10298_/Q _10282_/Q _08873_/Y _05831_/Y vssd1 vssd1 vccd1 vccd1 _08874_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07825_ _07814_/X _07815_/X _07823_/X _07824_/X vssd1 vssd1 vccd1 vccd1 _07825_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ _07710_/X _07715_/X _07716_/X _07755_/X vssd1 vssd1 vccd1 vccd1 _07756_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06707_ _08722_/A vssd1 vssd1 vccd1 vccd1 _06707_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _09414_/X _09425_/X _09414_/X _09425_/X vssd1 vssd1 vccd1 vccd1 _09426_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07687_ _10217_/Q _07687_/B _07698_/A vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__and3_1
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06638_ _10361_/Q vssd1 vssd1 vccd1 vccd1 _06638_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06569_ _10105_/Q vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__inv_2
X_09357_ _09352_/X _09356_/X _09352_/X _09356_/X vssd1 vssd1 vccd1 vccd1 _09359_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08308_ _08309_/A _08301_/Y _06273_/B vssd1 vssd1 vccd1 vccd1 _08308_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _09470_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09288_/X sky130_fd_sc_hd__or2_1
X_08239_ _06047_/X _06257_/B _08238_/Y vssd1 vssd1 vccd1 vccd1 _08239_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _10202_/CLK _10201_/D vssd1 vssd1 vccd1 vccd1 _10201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _10249_/CLK _10132_/D vssd1 vssd1 vccd1 vccd1 _10132_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _10399_/CLK _10063_/D vssd1 vssd1 vccd1 vccd1 _10063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05940_ _05939_/X _05927_/A _05101_/X _05928_/A _05934_/X vssd1 vssd1 vccd1 vccd1
+ _10227_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05871_ _05871_/A vssd1 vssd1 vccd1 vccd1 _05871_/X sky130_fd_sc_hd__clkbuf_2
X_08590_ _08179_/A _08557_/A _08559_/X _08554_/X vssd1 vssd1 vccd1 vccd1 _08591_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07610_ _07610_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__or2_1
X_07541_ _10211_/Q vssd1 vssd1 vccd1 vccd1 _07597_/A sky130_fd_sc_hd__inv_2
XFILLER_179_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07472_ _09933_/X vssd1 vssd1 vccd1 vccd1 _07552_/B sky130_fd_sc_hd__clkbuf_2
X_06423_ _10081_/Q _06443_/A _06421_/Y _06442_/A vssd1 vssd1 vccd1 vccd1 _06425_/A
+ sky130_fd_sc_hd__o22a_1
X_09211_ _09153_/X _09154_/X _09107_/Y _09155_/X vssd1 vssd1 vccd1 vccd1 _09211_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _09142_/A vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__buf_2
X_06354_ _06337_/Y _10135_/Q _06345_/A vssd1 vssd1 vccd1 vccd1 _06355_/A sky130_fd_sc_hd__o21ai_2
XFILLER_187_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05305_ _05305_/A _05329_/A vssd1 vssd1 vccd1 vccd1 _05325_/A sky130_fd_sc_hd__or2_1
XFILLER_135_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09073_ _09073_/A vssd1 vssd1 vccd1 vccd1 _09180_/C sky130_fd_sc_hd__inv_2
X_06285_ _06285_/A _06285_/B vssd1 vssd1 vccd1 vccd1 _06285_/X sky130_fd_sc_hd__or2_1
X_05236_ _05236_/A vssd1 vssd1 vccd1 vccd1 _05236_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_146_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08024_ _08024_/A _08024_/B vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__or2_1
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05167_ _05179_/A _05167_/B vssd1 vssd1 vccd1 vccd1 _10399_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _09064_/X _09062_/Y _09994_/S vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__mux2_1
X_05098_ _05028_/X _05094_/X _10415_/Q _05095_/X _05097_/X vssd1 vssd1 vccd1 vccd1
+ _10415_/D sky130_fd_sc_hd__a221o_1
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08926_ _08926_/A _08926_/B vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__or2_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _10284_/Q _07423_/Y _10284_/Q _07423_/Y vssd1 vssd1 vccd1 vccd1 _08857_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07808_ _07828_/A _09924_/X vssd1 vssd1 vccd1 vccd1 _07808_/X sky130_fd_sc_hd__or2_1
X_08788_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _08788_/X sky130_fd_sc_hd__or2_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07739_ _07633_/X _07645_/X _07633_/X _07645_/X vssd1 vssd1 vccd1 vccd1 _07739_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_111_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09409_ _09409_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09409_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _10334_/CLK _10115_/D vssd1 vssd1 vccd1 vccd1 _10115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10046_ _10450_/CLK _10046_/D vssd1 vssd1 vccd1 vccd1 _10046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06070_ _06070_/A vssd1 vssd1 vccd1 vccd1 _06070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05021_ _05468_/A vssd1 vssd1 vccd1 vccd1 _06182_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ _09759_/X _08184_/Y _10044_/Q vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__mux2_1
X_06972_ _09886_/X vssd1 vssd1 vccd1 vccd1 _07212_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08711_ _08711_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08711_/Y sky130_fd_sc_hd__nor2_1
X_09691_ _06504_/X input23/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05923_ _06183_/A _05923_/B vssd1 vssd1 vccd1 vccd1 _06137_/B sky130_fd_sc_hd__or2_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08642_ _06624_/Y _08636_/Y _06818_/B _08709_/B vssd1 vssd1 vccd1 vccd1 _08642_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05854_ _05852_/X _05853_/B _05853_/Y vssd1 vssd1 vccd1 vccd1 _05854_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08573_ _08801_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__or2_1
X_05785_ _08842_/B _10263_/Q vssd1 vssd1 vccd1 vccd1 _05785_/Y sky130_fd_sc_hd__nor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07524_ _07524_/A vssd1 vssd1 vccd1 vccd1 _07706_/A sky130_fd_sc_hd__inv_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07455_ _10280_/Q _07455_/B vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__or2_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06406_ _10142_/Q vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__inv_2
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07386_ _07386_/A vssd1 vssd1 vccd1 vccd1 _07413_/A sky130_fd_sc_hd__inv_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _09289_/A _09452_/B _09300_/A _09354_/D vssd1 vssd1 vccd1 vccd1 _09125_/X
+ sky130_fd_sc_hd__o22a_1
X_06337_ _10242_/Q vssd1 vssd1 vccd1 vccd1 _06337_/Y sky130_fd_sc_hd__inv_2
X_06268_ _06268_/A _08283_/A vssd1 vssd1 vccd1 vccd1 _06269_/B sky130_fd_sc_hd__or2_1
XFILLER_135_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _09055_/A _09055_/B _09193_/A vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__a21o_1
XFILLER_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05219_ _10377_/Q _05215_/X input42/X _05216_/X _05218_/X vssd1 vssd1 vccd1 vccd1
+ _10377_/D sky130_fd_sc_hd__o221a_1
X_08007_ _08007_/A vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__inv_2
X_06199_ _09703_/X _06196_/X _10104_/Q _06197_/X vssd1 vssd1 vccd1 vccd1 _10104_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _06614_/D _08299_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08909_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__or2_1
XFILLER_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09889_ _06832_/X _05873_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09889_/X sky130_fd_sc_hd__mux2_2
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput60 _09572_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput82 _09600_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput71 _09590_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_68_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10029_ _10448_/Q _09553_/X _08364_/Y _09554_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10029_/X sky130_fd_sc_hd__mux4_2
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05570_ _05570_/A vssd1 vssd1 vccd1 vccd1 _05570_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07240_ _06991_/Y _07228_/B _07233_/X _07236_/X vssd1 vssd1 vccd1 vccd1 _07247_/A
+ sky130_fd_sc_hd__o22ai_4
X_07171_ _07171_/A _07146_/X vssd1 vssd1 vccd1 vccd1 _07173_/A sky130_fd_sc_hd__or2b_1
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06122_ _06130_/A vssd1 vssd1 vccd1 vccd1 _06122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06053_ _09805_/X _06043_/X _06254_/A _06044_/X _06045_/X vssd1 vssd1 vccd1 vccd1
+ _10188_/D sky130_fd_sc_hd__o221a_1
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05004_ _05967_/A vssd1 vssd1 vccd1 vccd1 _08324_/C sky130_fd_sc_hd__clkbuf_2
X_09812_ _09811_/X _08237_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09812_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09743_ _06816_/Y _10408_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10074_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06955_ _06946_/A _06946_/B _06946_/X vssd1 vssd1 vccd1 vccd1 _06955_/X sky130_fd_sc_hd__a21bo_1
X_09674_ _10155_/Q _10171_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09674_/X sky130_fd_sc_hd__mux2_1
X_05906_ _10244_/Q _05902_/X input20/X _05903_/X _05900_/X vssd1 vssd1 vccd1 vccd1
+ _10244_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06886_ _06911_/A _09893_/X _07100_/A _06911_/B vssd1 vssd1 vccd1 vccd1 _06886_/X
+ sky130_fd_sc_hd__or4_4
X_08625_ _08625_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05837_ _05837_/A vssd1 vssd1 vccd1 vccd1 _07023_/A sky130_fd_sc_hd__inv_2
X_08556_ _06603_/X _10045_/Q _08461_/Y vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__a21oi_4
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ _10234_/Q _05768_/B vssd1 vssd1 vccd1 vccd1 _05771_/B sky130_fd_sc_hd__nor2_1
X_07507_ _07501_/X _07506_/X _07501_/X _07506_/X vssd1 vssd1 vccd1 vccd1 _07507_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ _10069_/Q _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__or2_1
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05699_ _05863_/A vssd1 vssd1 vccd1 vccd1 _05699_/X sky130_fd_sc_hd__buf_2
XFILLER_167_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07438_ _10275_/Q _07438_/B vssd1 vssd1 vccd1 vccd1 _07439_/B sky130_fd_sc_hd__or2_1
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07369_ _07315_/X _07368_/X _07315_/X _07368_/X vssd1 vssd1 vccd1 vccd1 _07369_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09108_ _09057_/Y _09060_/Y _09106_/X _09107_/Y vssd1 vssd1 vccd1 vccd1 _09108_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ _10414_/CLK _10380_/D vssd1 vssd1 vccd1 vccd1 _10380_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09039_ _08991_/X _08993_/X _08994_/X _08996_/X _09038_/X vssd1 vssd1 vccd1 vccd1
+ _09039_/X sky130_fd_sc_hd__o221a_1
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06740_ _06740_/A vssd1 vssd1 vccd1 vccd1 _06740_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06671_ _10359_/Q _08752_/A vssd1 vssd1 vccd1 vccd1 _06672_/B sky130_fd_sc_hd__or2_2
X_05622_ _10313_/Q vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__inv_2
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08410_ _09505_/X _08414_/B vssd1 vssd1 vccd1 vccd1 _08410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_196_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09390_ _09451_/A _09470_/B _09390_/C vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__or3_4
XFILLER_189_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05553_ _09923_/X _05552_/X _09923_/X _05552_/X vssd1 vssd1 vccd1 vccd1 _05641_/A
+ sky130_fd_sc_hd__a2bb2oi_1
X_08341_ _08998_/A vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ _08273_/A _08267_/Y _06265_/B vssd1 vssd1 vccd1 vccd1 _08272_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_149_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05484_ _10003_/X vssd1 vssd1 vccd1 vccd1 _05486_/A sky130_fd_sc_hd__inv_2
XFILLER_177_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater90 _09874_/S vssd1 vssd1 vccd1 vccd1 _09814_/S sky130_fd_sc_hd__buf_8
XFILLER_149_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07223_ _07223_/A _07223_/B _07223_/C vssd1 vssd1 vccd1 vccd1 _07223_/X sky130_fd_sc_hd__or3_1
XFILLER_164_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07154_ _07154_/A _07154_/B vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__or2_1
X_06105_ _10336_/Q _06101_/X _10164_/Q _06102_/X _06099_/X vssd1 vssd1 vccd1 vccd1
+ _10164_/D sky130_fd_sc_hd__a221o_1
X_07085_ _07080_/X _07084_/X _07080_/X _07084_/X vssd1 vssd1 vccd1 vccd1 _07254_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_06036_ _09837_/X _06028_/X _06035_/X _06031_/X _06032_/X vssd1 vssd1 vccd1 vccd1
+ _10196_/D sky130_fd_sc_hd__o221a_1
XFILLER_154_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _07953_/X _07973_/X _07953_/X _07973_/X vssd1 vssd1 vccd1 vccd1 _08004_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09726_ _06795_/Y _10391_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10057_/D sky130_fd_sc_hd__mux2_1
X_06938_ _06937_/A _06937_/B _06937_/Y vssd1 vssd1 vccd1 vccd1 _06938_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _10123_/Q input22/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__mux2_1
X_06869_ _09892_/X vssd1 vssd1 vccd1 vccd1 _07028_/B sky130_fd_sc_hd__clkbuf_2
X_08608_ _08299_/A _08497_/X _08607_/X vssd1 vssd1 vccd1 vccd1 _08608_/X sky130_fd_sc_hd__a21o_1
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _08426_/X _08425_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__mux2_2
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08539_ _08539_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _08593_/C sky130_fd_sc_hd__or2_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _10433_/CLK _10432_/D vssd1 vssd1 vccd1 vccd1 _10432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10363_ _10436_/CLK _10363_/D vssd1 vssd1 vccd1 vccd1 _10363_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10294_ _10297_/CLK _10294_/D vssd1 vssd1 vccd1 vccd1 _10294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08890_ _08890_/A vssd1 vssd1 vccd1 vccd1 _08890_/X sky130_fd_sc_hd__clkbuf_1
X_07910_ _07910_/A _07910_/B _07910_/C vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__or3_4
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _07836_/X _07840_/X _07836_/X _07840_/X vssd1 vssd1 vccd1 vccd1 _07882_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_07772_ _07916_/B _07910_/C vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06723_ _08745_/A vssd1 vssd1 vccd1 vccd1 _06723_/Y sky130_fd_sc_hd__inv_2
X_09511_ _09510_/X _09474_/A _09998_/S vssd1 vssd1 vccd1 vccd1 _09511_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09442_/X sky130_fd_sc_hd__or2_1
X_06654_ _10449_/Q vssd1 vssd1 vccd1 vccd1 _08459_/A sky130_fd_sc_hd__inv_2
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06585_ _10108_/Q vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__inv_2
X_09373_ _09373_/A vssd1 vssd1 vccd1 vccd1 _09373_/Y sky130_fd_sc_hd__inv_2
X_05605_ _09923_/X _05552_/X _05640_/A vssd1 vssd1 vccd1 vccd1 _05605_/X sky130_fd_sc_hd__o21a_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08324_ _08324_/A _08324_/B _08324_/C vssd1 vssd1 vccd1 vccd1 _09554_/S sky130_fd_sc_hd__nor3_4
X_05536_ _05469_/X _05529_/X _05469_/X _05529_/X vssd1 vssd1 vccd1 vccd1 _05536_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__or2_2
X_05467_ _05741_/A vssd1 vssd1 vccd1 vccd1 _05467_/X sky130_fd_sc_hd__buf_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ _10178_/Q _08186_/B vssd1 vssd1 vccd1 vccd1 _08191_/B sky130_fd_sc_hd__nand2_2
X_05398_ _05399_/A vssd1 vssd1 vccd1 vccd1 _06130_/A sky130_fd_sc_hd__clkbuf_4
X_07206_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07206_/X sky130_fd_sc_hd__or2_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07137_ _07137_/A _07137_/B vssd1 vssd1 vccd1 vccd1 _07138_/B sky130_fd_sc_hd__or2_1
XFILLER_145_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07068_ _07068_/A _07118_/B _07068_/C vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__or3_1
X_06019_ _09861_/X _06015_/X _06268_/A _06017_/X _06018_/X vssd1 vssd1 vccd1 vccd1
+ _10202_/D sky130_fd_sc_hd__o221a_1
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE2_1 _09451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _06597_/X input43/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09709_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _10422_/CLK _10415_/D vssd1 vssd1 vccd1 vccd1 _10415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10346_ _10346_/CLK _10346_/D vssd1 vssd1 vccd1 vccd1 _10346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10277_ _10298_/CLK _10277_/D vssd1 vssd1 vccd1 vccd1 _10277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06370_ _06370_/A _10138_/Q vssd1 vssd1 vccd1 vccd1 _06370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05321_ _10175_/Q vssd1 vssd1 vccd1 vccd1 _05336_/A sky130_fd_sc_hd__buf_1
X_05252_ _05264_/A vssd1 vssd1 vccd1 vccd1 _05252_/X sky130_fd_sc_hd__buf_1
X_08040_ _08022_/A _08022_/B _08023_/B vssd1 vssd1 vccd1 vccd1 _08040_/X sky130_fd_sc_hd__a21bo_1
X_05183_ _05193_/A _05181_/Y _05182_/Y _05161_/A vssd1 vssd1 vccd1 vccd1 _05184_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09991_ _08045_/X _07395_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09991_/X sky130_fd_sc_hd__mux2_2
X_08942_ _08942_/A _08995_/A vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08873_ _10298_/Q vssd1 vssd1 vccd1 vccd1 _08873_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07824_ _07855_/A _07897_/B _07824_/C vssd1 vssd1 vccd1 vccd1 _07824_/X sky130_fd_sc_hd__or3_1
XFILLER_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07755_ _07717_/X _07727_/X _07728_/X _07754_/X vssd1 vssd1 vccd1 vccd1 _07755_/X
+ sky130_fd_sc_hd__o22a_1
X_06706_ _10370_/Q vssd1 vssd1 vccd1 vccd1 _06706_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07686_ _07686_/A _07686_/B vssd1 vssd1 vccd1 vccd1 _07698_/A sky130_fd_sc_hd__or2_1
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _09424_/A _09424_/B _09424_/X vssd1 vssd1 vccd1 vccd1 _09425_/X sky130_fd_sc_hd__a21bo_1
X_06637_ _10393_/Q vssd1 vssd1 vccd1 vccd1 _06637_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06568_ _06566_/X _06567_/Y _06566_/X _06567_/Y vssd1 vssd1 vccd1 vccd1 _06568_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09356_ _09356_/A _09356_/B vssd1 vssd1 vccd1 vccd1 _09356_/X sky130_fd_sc_hd__or2_1
X_08307_ _08307_/A vssd1 vssd1 vccd1 vccd1 _08309_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09287_ _09354_/D vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__clkbuf_2
X_06499_ _06499_/A vssd1 vssd1 vccd1 vccd1 _06499_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05519_ _09993_/X _10005_/X _05494_/Y _05570_/A vssd1 vssd1 vccd1 vccd1 _05519_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08238_ _08238_/A vssd1 vssd1 vccd1 vccd1 _08238_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _10202_/CLK _10200_/D vssd1 vssd1 vccd1 vccd1 _10200_/Q sky130_fd_sc_hd__dfxtp_2
X_08169_ _08281_/A vssd1 vssd1 vccd1 vccd1 _08169_/X sky130_fd_sc_hd__buf_2
XFILLER_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _10249_/CLK _10131_/D vssd1 vssd1 vccd1 vccd1 _10131_/Q sky130_fd_sc_hd__dfxtp_2
X_10062_ _10399_/CLK _10062_/D vssd1 vssd1 vccd1 vccd1 _10062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10329_ _10329_/CLK _10329_/D vssd1 vssd1 vccd1 vccd1 _10329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05870_ _10256_/Q _05851_/X _05863_/X _06828_/A _05866_/X vssd1 vssd1 vccd1 vccd1
+ _10256_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07540_ _07819_/A _09933_/X vssd1 vssd1 vccd1 vccd1 _07540_/X sky130_fd_sc_hd__or2_1
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07471_ _07537_/D vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_201_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09210_ _09208_/X _09209_/X _09208_/X _09209_/X vssd1 vssd1 vccd1 vccd1 _09210_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06422_ _06443_/A vssd1 vssd1 vccd1 vccd1 _06442_/A sky130_fd_sc_hd__inv_2
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09141_ _09139_/Y _09140_/Y _09139_/Y _09140_/Y vssd1 vssd1 vccd1 vccd1 _09141_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06353_ _06353_/A vssd1 vssd1 vccd1 vccd1 _06353_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09292_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__or2_2
X_05304_ _05304_/A _05334_/A vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__or2_1
X_06284_ _06275_/Y _10128_/Q _05771_/B _06277_/Y vssd1 vssd1 vccd1 vccd1 _06285_/B
+ sky130_fd_sc_hd__o22a_1
X_08023_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__or2_1
X_05235_ _10367_/Q vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__buf_2
X_05166_ _05153_/X _06616_/D _05165_/Y _05161_/X vssd1 vssd1 vccd1 vccd1 _05167_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _08951_/X _08949_/A _09986_/S vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__mux2_2
X_05097_ _05274_/A vssd1 vssd1 vccd1 vccd1 _05097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08925_ _08926_/B vssd1 vssd1 vccd1 vccd1 _08925_/Y sky130_fd_sc_hd__inv_2
X_08856_ _10285_/Q _07421_/Y _10285_/Q _07421_/Y vssd1 vssd1 vccd1 vccd1 _08895_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07807_ _07830_/A _07878_/D vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__or2_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05999_ _10207_/Q vssd1 vssd1 vccd1 vccd1 _06000_/A sky130_fd_sc_hd__clkbuf_2
X_08787_ _06603_/X _06621_/A _08628_/A _08626_/Y _08628_/Y vssd1 vssd1 vccd1 vccd1
+ _08791_/B sky130_fd_sc_hd__o32a_1
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07738_ _07737_/A _07737_/B _07737_/X vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__a21boi_4
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07669_ _07672_/C _07669_/B vssd1 vssd1 vccd1 vccd1 _07669_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _09408_/A _09452_/B _09288_/X vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__or3b_1
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09339_ _09457_/C _09922_/X _09468_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09341_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10334_/CLK _10114_/D vssd1 vssd1 vccd1 vccd1 _10114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ _10450_/CLK _10045_/D vssd1 vssd1 vccd1 vccd1 _10045_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05020_ _05034_/A vssd1 vssd1 vccd1 vccd1 _05468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06971_ _07210_/A vssd1 vssd1 vccd1 vccd1 _07311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08710_ _08707_/A _08709_/B _06626_/Y _08709_/Y vssd1 vssd1 vccd1 vccd1 _08710_/X
+ sky130_fd_sc_hd__o22a_1
X_05922_ _09170_/A vssd1 vssd1 vccd1 vccd1 _05922_/X sky130_fd_sc_hd__clkbuf_2
X_09690_ _06500_/X input22/X _09944_/S vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__mux2_1
X_08641_ _08713_/B vssd1 vssd1 vccd1 vccd1 _08709_/B sky130_fd_sc_hd__buf_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05853_ _05853_/A _05853_/B vssd1 vssd1 vccd1 vccd1 _05853_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ _08545_/Y _08547_/X _08570_/Y _08591_/C vssd1 vssd1 vccd1 vccd1 _08572_/Y
+ sky130_fd_sc_hd__a31oi_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05784_ _10281_/Q _10264_/Q _07854_/A _05783_/Y vssd1 vssd1 vccd1 vccd1 _05784_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07523_ _07523_/A _07529_/A vssd1 vssd1 vccd1 vccd1 _07523_/Y sky130_fd_sc_hd__nor2_1
XFILLER_179_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07454_ _10279_/Q _07454_/B vssd1 vssd1 vccd1 vccd1 _07455_/B sky130_fd_sc_hd__or2_1
XFILLER_210_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06405_ _10249_/Q vssd1 vssd1 vccd1 vccd1 _06405_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07385_ _07385_/A vssd1 vssd1 vccd1 vccd1 _07385_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ _09976_/X vssd1 vssd1 vccd1 vccd1 _09354_/D sky130_fd_sc_hd__clkbuf_2
X_06336_ _06332_/Y _06335_/X _06332_/Y _06335_/X vssd1 vssd1 vccd1 vccd1 _06336_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06267_ _10201_/Q _06267_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__or2_1
XFILLER_175_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _09055_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05218_ _05236_/A vssd1 vssd1 vccd1 vccd1 _05218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08006_ _08006_/A vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__inv_2
XFILLER_190_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06198_ _09704_/X _06196_/X _10105_/Q _06197_/X vssd1 vssd1 vccd1 vccd1 _10105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05149_ _10402_/Q vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__inv_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _09956_/X _06633_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08908_ _08909_/A vssd1 vssd1 vccd1 vccd1 _08908_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _06831_/X _05869_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__mux2_1
X_08839_ _08839_/A _09583_/S _09600_/S vssd1 vssd1 vccd1 vccd1 _08839_/X sky130_fd_sc_hd__or3b_4
XFILLER_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput61 _09575_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput72 _09591_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput83 _10027_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[3] sky130_fd_sc_hd__clkbuf_2
X_10028_ _10447_/Q _09550_/X _08356_/Y _09551_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10028_/X sky130_fd_sc_hd__mux4_2
XFILLER_209_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07170_ _07164_/A _07212_/B _07146_/C _07218_/B vssd1 vssd1 vccd1 vccd1 _07171_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06121_ _10153_/Q _06117_/X _10325_/Q _06113_/X _06120_/X vssd1 vssd1 vccd1 vccd1
+ _10153_/D sky130_fd_sc_hd__o221a_1
X_06052_ _10188_/Q vssd1 vssd1 vccd1 vccd1 _06254_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05003_ input11/X _08329_/C vssd1 vssd1 vccd1 vccd1 _05967_/A sky130_fd_sc_hd__or2_1
XFILLER_207_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09811_ _10361_/Q _09810_/X _10043_/Q vssd1 vssd1 vccd1 vccd1 _09811_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09742_ _06815_/Y _10407_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10073_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06954_ _06950_/X _06951_/X _06950_/X _06951_/X vssd1 vssd1 vccd1 vccd1 _06958_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09673_ _10154_/Q _10170_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__mux2_1
X_05905_ _10245_/Q _05902_/X input21/X _05903_/X _05900_/X vssd1 vssd1 vccd1 vccd1
+ _10245_/D sky130_fd_sc_hd__o221a_1
X_06885_ _06885_/A _06884_/X vssd1 vssd1 vccd1 vccd1 _06885_/X sky130_fd_sc_hd__or2b_1
X_08624_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05836_ _05784_/X _05829_/X _05784_/X _05829_/X vssd1 vssd1 vccd1 vccd1 _05837_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08555_ _06603_/X _10045_/Q _08463_/A _08461_/Y _08463_/Y vssd1 vssd1 vccd1 vccd1
+ _08558_/B sky130_fd_sc_hd__o32a_1
X_05767_ _10127_/Q vssd1 vssd1 vccd1 vccd1 _05768_/B sky130_fd_sc_hd__inv_2
XFILLER_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07506_/X sky130_fd_sc_hd__or2_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08486_ _10068_/Q _08502_/A vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__or2_1
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05698_ _08618_/A _05698_/B vssd1 vssd1 vccd1 vccd1 _10299_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07437_ _07437_/A vssd1 vssd1 vccd1 vccd1 _07437_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07368_ _07364_/Y _07367_/Y _07364_/Y _07367_/Y vssd1 vssd1 vccd1 vccd1 _07368_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09107_ _09057_/Y _09060_/Y _09106_/X vssd1 vssd1 vccd1 vccd1 _09107_/Y sky130_fd_sc_hd__o21ai_2
X_06319_ _10133_/Q vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__inv_2
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07299_ _07299_/A vssd1 vssd1 vccd1 vccd1 _07299_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ _09038_/A _09096_/A _09038_/C vssd1 vssd1 vccd1 vccd1 _09038_/X sky130_fd_sc_hd__or3_2
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06670_ _10358_/Q _06670_/B vssd1 vssd1 vccd1 vccd1 _08752_/A sky130_fd_sc_hd__or2_2
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05621_ _05621_/A _05621_/B vssd1 vssd1 vccd1 vccd1 _05621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08340_ _08934_/A vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__buf_1
X_05552_ _05550_/Y _05551_/Y _05550_/Y _05551_/Y vssd1 vssd1 vccd1 vccd1 _05552_/X
+ sky130_fd_sc_hd__a2bb2o_4
X_08271_ _08269_/A _08269_/B _08240_/X _08270_/Y vssd1 vssd1 vccd1 vccd1 _08271_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_189_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05483_ _09992_/X _10021_/X _09992_/X _10021_/X vssd1 vssd1 vccd1 vccd1 _05483_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07222_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07222_/X sky130_fd_sc_hd__or2_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater91 _09878_/S vssd1 vssd1 vccd1 vccd1 _09874_/S sky130_fd_sc_hd__buf_8
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07155_/C _07151_/X _07384_/A vssd1 vssd1 vccd1 vccd1 _07154_/B sky130_fd_sc_hd__a21oi_2
XFILLER_157_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06104_ _10337_/Q _06101_/X _10165_/Q _06102_/X _06099_/X vssd1 vssd1 vccd1 vccd1
+ _10165_/D sky130_fd_sc_hd__a221o_1
XFILLER_172_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07084_ _07074_/B _07083_/A _07073_/A _07083_/Y vssd1 vssd1 vccd1 vccd1 _07084_/X
+ sky130_fd_sc_hd__a22o_1
X_06035_ _06262_/A vssd1 vssd1 vccd1 vccd1 _06035_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07986_ _07947_/X _07974_/X _07947_/X _07974_/X vssd1 vssd1 vccd1 vccd1 _08003_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09725_ _06794_/Y _10390_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10056_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06937_ _06937_/A _06937_/B vssd1 vssd1 vccd1 vccd1 _06937_/Y sky130_fd_sc_hd__nor2_1
X_09656_ _10122_/Q input21/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09656_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08607_ _08297_/A _08497_/X _08294_/A _08498_/X _08606_/X vssd1 vssd1 vccd1 vccd1
+ _08607_/X sky130_fd_sc_hd__o221a_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06868_ _06911_/B vssd1 vssd1 vccd1 vccd1 _06868_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09587_ _08424_/Y _08423_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09587_/X sky130_fd_sc_hd__mux2_2
X_06799_ _06802_/A _06799_/B vssd1 vssd1 vccd1 vccd1 _06799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05819_ _08852_/B _05806_/Y _05807_/X _05818_/X vssd1 vssd1 vccd1 vccd1 _05819_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _10057_/Q _08475_/B _08476_/B vssd1 vssd1 vccd1 vccd1 _08539_/B sky130_fd_sc_hd__a21bo_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _10051_/Q _08469_/B vssd1 vssd1 vccd1 vccd1 _08470_/B sky130_fd_sc_hd__or2_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10431_ _10433_/CLK _10431_/D vssd1 vssd1 vccd1 vccd1 _10431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10362_ _10436_/CLK _10362_/D vssd1 vssd1 vccd1 vccd1 _10362_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_151_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10293_ _10297_/CLK _10293_/D vssd1 vssd1 vccd1 vccd1 _10293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07840_ _07830_/C _07839_/A _07829_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _07840_/X
+ sky130_fd_sc_hd__a22o_1
X_07771_ _07766_/A _07777_/B _07770_/X vssd1 vssd1 vccd1 vccd1 _07910_/C sky130_fd_sc_hd__o21ai_2
X_06722_ _10362_/Q vssd1 vssd1 vccd1 vccd1 _06722_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _08405_/X _06390_/A _09997_/S vssd1 vssd1 vccd1 vccd1 _09510_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09441_ _09441_/A vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__inv_2
X_06653_ _10350_/Q vssd1 vssd1 vccd1 vccd1 _06653_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06584_ _06583_/A _06583_/B _06591_/A vssd1 vssd1 vccd1 vccd1 _06584_/Y sky130_fd_sc_hd__a21boi_1
X_09372_ _09370_/Y _09430_/B _09370_/Y _09430_/B vssd1 vssd1 vccd1 vccd1 _09373_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_05604_ _05641_/A _05641_/B vssd1 vssd1 vccd1 vccd1 _05640_/A sky130_fd_sc_hd__nand2_1
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08323_ _09752_/X _08839_/A vssd1 vssd1 vccd1 vccd1 _08323_/X sky130_fd_sc_hd__and2_1
X_05535_ _05530_/Y _05534_/Y _05530_/Y _05534_/Y vssd1 vssd1 vccd1 vccd1 _05615_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08254_ _08253_/X _08247_/Y _06261_/B vssd1 vssd1 vccd1 vccd1 _08254_/Y sky130_fd_sc_hd__o21ai_1
X_05466_ _05750_/A vssd1 vssd1 vccd1 vccd1 _05741_/A sky130_fd_sc_hd__buf_1
X_08185_ _08554_/A _08182_/A _06245_/B vssd1 vssd1 vccd1 vccd1 _08185_/Y sky130_fd_sc_hd__o21ai_1
X_05397_ _10330_/Q vssd1 vssd1 vccd1 vccd1 _05397_/Y sky130_fd_sc_hd__inv_2
X_07205_ _07133_/A _07139_/A _07133_/Y vssd1 vssd1 vccd1 vccd1 _07206_/B sky130_fd_sc_hd__a21o_1
XFILLER_20_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07136_ _07112_/C _07109_/B _07109_/Y vssd1 vssd1 vccd1 vccd1 _07137_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07067_ _07067_/A _07067_/B vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__or2_1
X_06018_ _06032_/A vssd1 vssd1 vccd1 vccd1 _06018_/X sky130_fd_sc_hd__buf_1
XFILLER_121_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XINSDIODE2_2 _09470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _06593_/Y input42/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _07820_/C _07968_/X _07820_/C _07968_/X vssd1 vssd1 vccd1 vccd1 _07969_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ _06365_/X _06368_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09639_/X sky130_fd_sc_hd__mux2_2
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _10414_/CLK _10414_/D vssd1 vssd1 vccd1 vccd1 _10414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10345_ _10346_/CLK _10345_/D vssd1 vssd1 vccd1 vccd1 _10345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10276_ _10298_/CLK _10276_/D vssd1 vssd1 vccd1 vccd1 _10276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05320_ _10343_/Q _05320_/B vssd1 vssd1 vccd1 vccd1 _05320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05251_ _05263_/A vssd1 vssd1 vccd1 vccd1 _05251_/X sky130_fd_sc_hd__buf_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05182_ _10427_/Q vssd1 vssd1 vccd1 vccd1 _05182_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _08047_/X _07396_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09990_/X sky130_fd_sc_hd__mux2_2
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08941_ _08938_/X _08940_/X _08938_/X _08940_/X vssd1 vssd1 vccd1 vccd1 _08943_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_08872_ _10297_/Q _05782_/X _08840_/X _08871_/X vssd1 vssd1 vccd1 vccd1 _08872_/X
+ sky130_fd_sc_hd__o22a_2
X_07823_ _07823_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07823_/X sky130_fd_sc_hd__or2_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07754_ _07729_/X _07733_/X _07734_/X _07753_/Y vssd1 vssd1 vccd1 vccd1 _07754_/X
+ sky130_fd_sc_hd__o22a_1
X_06705_ _10371_/Q _08719_/A _06703_/Y vssd1 vssd1 vccd1 vccd1 _06811_/B sky130_fd_sc_hd__a21oi_2
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07685_ _07671_/X _07672_/X _07671_/X _07672_/X vssd1 vssd1 vccd1 vccd1 _07685_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_52_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06636_ _10363_/Q vssd1 vssd1 vccd1 vccd1 _06636_/Y sky130_fd_sc_hd__inv_2
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__or2_1
XFILLER_44_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06567_ _08436_/A _06438_/X _06563_/X vssd1 vssd1 vccd1 vccd1 _06567_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_178_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09355_ _09355_/A vssd1 vssd1 vccd1 vccd1 _09356_/B sky130_fd_sc_hd__inv_2
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ _08304_/A _08304_/B _08193_/X _08305_/Y vssd1 vssd1 vccd1 vccd1 _08306_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_193_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09286_ _05922_/X _09418_/A _09423_/A _09285_/Y vssd1 vssd1 vccd1 vccd1 _09286_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06498_ _06498_/A _06498_/B vssd1 vssd1 vccd1 vccd1 _06499_/A sky130_fd_sc_hd__nand2_2
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05518_ _10002_/X _10001_/X _05497_/Y _05574_/A vssd1 vssd1 vccd1 vccd1 _05570_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08237_ _08751_/A _08233_/Y _08219_/X _08241_/B vssd1 vssd1 vccd1 vccd1 _08237_/X
+ sky130_fd_sc_hd__o211a_1
X_05449_ _10319_/Q _05449_/B vssd1 vssd1 vccd1 vccd1 _05449_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08168_ _08599_/A vssd1 vssd1 vccd1 vccd1 _08281_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_180_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08099_ _10206_/Q vssd1 vssd1 vccd1 vccd1 _08307_/A sky130_fd_sc_hd__inv_2
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07119_ _07115_/X _07118_/X _07115_/X _07118_/X vssd1 vssd1 vccd1 vccd1 _07119_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10447_/CLK _10130_/D vssd1 vssd1 vccd1 vccd1 _10130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _10399_/CLK _10061_/D vssd1 vssd1 vccd1 vccd1 _10061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10328_ _10328_/CLK _10328_/D vssd1 vssd1 vccd1 vccd1 _10328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10259_ _10274_/CLK _10259_/D vssd1 vssd1 vccd1 vccd1 _10259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07470_ _09935_/X vssd1 vssd1 vccd1 vccd1 _07537_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_201_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06421_ _10081_/Q vssd1 vssd1 vccd1 vccd1 _06421_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ _09085_/A _09084_/Y _09187_/A vssd1 vssd1 vccd1 vccd1 _09140_/Y sky130_fd_sc_hd__o21ai_1
X_06352_ _06352_/A _06352_/B vssd1 vssd1 vccd1 vccd1 _06353_/A sky130_fd_sc_hd__or2_2
XFILLER_175_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05303_ _05303_/A _05339_/A vssd1 vssd1 vccd1 vccd1 _05334_/A sky130_fd_sc_hd__or2_1
X_09071_ _09037_/X _09039_/X _09024_/X _09040_/X vssd1 vssd1 vccd1 vccd1 _09087_/A
+ sky130_fd_sc_hd__o22a_1
X_06283_ _06283_/A vssd1 vssd1 vccd1 vccd1 _06285_/A sky130_fd_sc_hd__inv_2
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08022_ _08022_/A _08022_/B vssd1 vssd1 vccd1 vccd1 _08023_/B sky130_fd_sc_hd__or2_1
X_05234_ _10368_/Q _05230_/X input32/X _05231_/X _05227_/X vssd1 vssd1 vccd1 vccd1
+ _10368_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05165_ _10431_/Q vssd1 vssd1 vccd1 vccd1 _05165_/Y sky130_fd_sc_hd__inv_2
X_09973_ _09814_/S _08176_/X _10044_/Q vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05096_ _05093_/X _05094_/X _10416_/Q _05095_/X _05086_/X vssd1 vssd1 vccd1 vccd1
+ _10416_/D sky130_fd_sc_hd__a221o_1
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08924_ _08923_/A _08923_/B _08995_/A vssd1 vssd1 vccd1 vccd1 _08926_/B sky130_fd_sc_hd__a21oi_2
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08855_ _08855_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08855_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08786_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__and2_1
X_07806_ _07806_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07806_/X sky130_fd_sc_hd__or2_1
X_05998_ _06028_/A vssd1 vssd1 vccd1 vccd1 _05998_/X sky130_fd_sc_hd__clkbuf_2
X_07737_ _07737_/A _07737_/B vssd1 vssd1 vccd1 vccd1 _07737_/X sky130_fd_sc_hd__or2_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07668_ _10215_/Q _07687_/B _07747_/A vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__and3_1
XFILLER_197_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06619_ _06809_/A vssd1 vssd1 vccd1 vccd1 _06620_/A sky130_fd_sc_hd__inv_2
X_09407_ _10232_/Q _09405_/Y _05933_/X _09232_/Y _09406_/X vssd1 vssd1 vccd1 vccd1
+ _09409_/A sky130_fd_sc_hd__a41o_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07599_ _07585_/X _07587_/X _07585_/X _07587_/X vssd1 vssd1 vccd1 vccd1 _07599_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09338_ _09326_/X _09327_/X _09328_/X _09329_/X vssd1 vssd1 vccd1 vccd1 _09338_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09269_ _09267_/X _09269_/B vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__and2b_1
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10113_ _10334_/CLK _10113_/D vssd1 vssd1 vccd1 vccd1 _10113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10044_ _10450_/CLK _10044_/D vssd1 vssd1 vccd1 vccd1 _10044_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_208_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06970_ _06970_/A vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__inv_2
X_05921_ _10233_/Q vssd1 vssd1 vccd1 vccd1 _09170_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08640_ _08717_/B vssd1 vssd1 vccd1 vccd1 _08713_/B sky130_fd_sc_hd__buf_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05852_ _05853_/A vssd1 vssd1 vccd1 vccd1 _05852_/X sky130_fd_sc_hd__clkbuf_2
X_08571_ _08774_/A _08547_/B _08215_/A _08542_/A vssd1 vssd1 vccd1 vccd1 _08591_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05783_ _10264_/Q vssd1 vssd1 vccd1 vccd1 _05783_/Y sky130_fd_sc_hd__inv_2
X_07522_ _07505_/A _07517_/Y _07514_/X _07518_/X vssd1 vssd1 vccd1 vccd1 _07529_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07453_ _08842_/B vssd1 vssd1 vccd1 vccd1 _07453_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06404_ _06397_/Y _10141_/Q _06399_/A _06401_/X vssd1 vssd1 vccd1 vccd1 _06404_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09123_ _09229_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__clkbuf_2
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__or2_1
X_06335_ _10240_/Q _08370_/A _06322_/Y _06327_/A vssd1 vssd1 vccd1 vccd1 _06335_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06266_ _10200_/Q _08275_/A vssd1 vssd1 vccd1 vccd1 _06267_/B sky130_fd_sc_hd__or2_1
XFILLER_175_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _09053_/A _09053_/B _09100_/A vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__a21o_1
XFILLER_190_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05217_ _10378_/Q _05215_/X input43/X _05216_/X _05206_/X vssd1 vssd1 vccd1 vccd1
+ _10378_/D sky130_fd_sc_hd__o221a_1
X_08005_ _08005_/A vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__inv_2
X_06197_ _06204_/A vssd1 vssd1 vccd1 vccd1 _06197_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05148_ _05157_/A _05148_/B vssd1 vssd1 vccd1 vccd1 _10403_/D sky130_fd_sc_hd__nor2_1
XFILLER_143_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _06616_/D _08265_/A _09981_/S vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__mux2_1
X_05079_ _10424_/Q _05072_/X input23/X _05073_/X _05078_/X vssd1 vssd1 vccd1 vccd1
+ _10424_/D sky130_fd_sc_hd__o221a_1
XFILLER_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08907_ _08860_/X _08909_/B _08860_/X _08909_/B vssd1 vssd1 vccd1 vccd1 _08907_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09887_ _06830_/X _05865_/A _10022_/S vssd1 vssd1 vccd1 vccd1 _09887_/X sky130_fd_sc_hd__mux2_2
X_08838_ _06273_/A _08642_/X _08706_/Y _08837_/X vssd1 vssd1 vccd1 vccd1 _10077_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_106_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08769_ _08215_/A _08767_/X _10186_/Q _08801_/B vssd1 vssd1 vccd1 vccd1 _08769_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput73 _09592_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput62 _09578_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput84 _10028_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[4] sky130_fd_sc_hd__clkbuf_2
X_10027_ _10446_/Q _09547_/X _08350_/Y _09548_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10027_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06120_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06120_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06051_ _09809_/X _06043_/X _10189_/Q _06044_/X _06045_/X vssd1 vssd1 vccd1 vccd1
+ _10189_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05002_ input12/X _05775_/A vssd1 vssd1 vccd1 vccd1 _08329_/C sky130_fd_sc_hd__or2_1
XFILLER_207_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09810_ _08235_/Y _10361_/Q _09814_/S vssd1 vssd1 vccd1 vccd1 _09810_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _06814_/Y _10406_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10072_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06953_ _06940_/X _06952_/X _06940_/X _06952_/X vssd1 vssd1 vccd1 vccd1 _06953_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05904_ _10246_/Q _05902_/X input22/X _05903_/X _05900_/X vssd1 vssd1 vccd1 vccd1
+ _10246_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _10153_/Q _10169_/Q _10175_/Q vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06884_ _06962_/A _07031_/B _07118_/A _09892_/X vssd1 vssd1 vccd1 vccd1 _06884_/X
+ sky130_fd_sc_hd__or4_4
X_08623_ _08623_/A _09937_/X vssd1 vssd1 vccd1 vccd1 _10044_/D sky130_fd_sc_hd__or2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05835_ _10265_/Q _05780_/X _05637_/X _05834_/Y _05764_/X vssd1 vssd1 vccd1 vccd1
+ _10265_/D sky130_fd_sc_hd__o221a_1
X_08554_ _08554_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _08554_/X sky130_fd_sc_hd__or2_1
X_05766_ _07423_/A _05759_/X _09630_/X _05761_/X _05764_/X vssd1 vssd1 vccd1 vccd1
+ _10268_/D sky130_fd_sc_hd__o221a_1
XFILLER_42_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07505_ _07505_/A vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__inv_2
XFILLER_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08485_ _10067_/Q _08485_/B vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__or2_1
XFILLER_195_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05697_ _05771_/A _05694_/Y _05695_/X _08059_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05698_/B sky130_fd_sc_hd__o32a_1
XFILLER_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07436_ _07434_/X _07419_/Y _07428_/B vssd1 vssd1 vccd1 vccd1 _07436_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ _07365_/Y _07366_/X _07365_/Y _07366_/X vssd1 vssd1 vccd1 vccd1 _07367_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_163_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09104_/A _09105_/A _09201_/C _09105_/Y vssd1 vssd1 vccd1 vccd1 _09106_/X
+ sky130_fd_sc_hd__o22a_1
X_06318_ _06313_/A _06317_/X _06313_/A _06317_/X vssd1 vssd1 vccd1 vccd1 _06318_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09036_/A _09036_/B _09083_/B vssd1 vssd1 vccd1 vccd1 _09037_/X sky130_fd_sc_hd__a21o_1
X_07298_ _07283_/X _07296_/Y _07297_/X vssd1 vssd1 vccd1 vccd1 _07299_/A sky130_fd_sc_hd__a21oi_2
X_06249_ _10183_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__or2_1
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _08927_/X _08925_/Y _09986_/S vssd1 vssd1 vccd1 vccd1 _09939_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05620_ _05620_/A vssd1 vssd1 vccd1 vccd1 _05620_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05551_ _05481_/A _05481_/B _05481_/Y vssd1 vssd1 vccd1 vccd1 _05551_/Y sky130_fd_sc_hd__a21oi_2
X_08270_ _08273_/B vssd1 vssd1 vccd1 vccd1 _08270_/Y sky130_fd_sc_hd__inv_2
X_05482_ _10023_/X _10022_/X _10023_/X _10022_/X vssd1 vssd1 vccd1 vccd1 _05482_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07221_ _07063_/A _07212_/B _07223_/A _07218_/B _07220_/Y vssd1 vssd1 vccd1 vccd1
+ _07222_/B sky130_fd_sc_hd__o41a_1
XFILLER_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater92 _09986_/S vssd1 vssd1 vccd1 vccd1 _09994_/S sky130_fd_sc_hd__buf_8
X_07152_ _10218_/Q _07152_/B _10219_/Q _07152_/D vssd1 vssd1 vccd1 vccd1 _07384_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_145_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06103_ _10338_/Q _06101_/X _10166_/Q _06102_/X _06099_/X vssd1 vssd1 vccd1 vccd1
+ _10166_/D sky130_fd_sc_hd__a221o_1
XFILLER_133_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07083_ _07083_/A vssd1 vssd1 vccd1 vccd1 _07083_/Y sky130_fd_sc_hd__inv_2
X_06034_ _10196_/Q vssd1 vssd1 vccd1 vccd1 _06262_/A sky130_fd_sc_hd__buf_2
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07985_ _07940_/X _07975_/X _07940_/X _07975_/X vssd1 vssd1 vccd1 vccd1 _08002_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09724_ _06793_/X _10389_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10055_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06936_ _06961_/A _09894_/X _06935_/X vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__or3b_1
X_09655_ _10121_/Q input20/X _10266_/Q vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06867_ _09668_/X vssd1 vssd1 vccd1 vccd1 _06911_/B sky130_fd_sc_hd__clkbuf_2
X_08606_ _08293_/A _08498_/X _08605_/X vssd1 vssd1 vccd1 vccd1 _08606_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05818_ _07434_/A _05809_/Y _05810_/X _05817_/X vssd1 vssd1 vccd1 vccd1 _05818_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09586_ _08422_/Y _08420_/Y _09600_/S vssd1 vssd1 vccd1 vccd1 _09586_/X sky130_fd_sc_hd__mux2_2
X_06798_ _06802_/A _06798_/B vssd1 vssd1 vccd1 vccd1 _06798_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08765_/A _08574_/B vssd1 vssd1 vccd1 vccd1 _08537_/X sky130_fd_sc_hd__or2_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05749_ _08845_/B _05741_/X _09640_/X _05743_/X _05747_/X vssd1 vssd1 vccd1 vccd1
+ _10278_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08468_ _10050_/Q _08468_/B vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__or2_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _07427_/B vssd1 vssd1 vccd1 vccd1 _07419_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10430_ _10433_/CLK _10430_/D vssd1 vssd1 vccd1 vccd1 _10430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08399_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10361_ _10436_/CLK _10361_/D vssd1 vssd1 vccd1 vccd1 _10361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10292_ _10297_/CLK _10292_/D vssd1 vssd1 vccd1 vccd1 _10292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07770_ _07770_/A vssd1 vssd1 vccd1 vccd1 _07770_/X sky130_fd_sc_hd__buf_1
X_06721_ _10363_/Q _08742_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _06801_/B sky130_fd_sc_hd__a21oi_4
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09440_ _09438_/X _09439_/X _09438_/X _09439_/X vssd1 vssd1 vccd1 vccd1 _09441_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06652_ _08624_/A _10351_/Q vssd1 vssd1 vccd1 vccd1 _06652_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06583_ _06583_/A _06583_/B vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__or2_1
X_09371_ _09462_/C _09312_/Y _09313_/X _09317_/X vssd1 vssd1 vccd1 vccd1 _09430_/B
+ sky130_fd_sc_hd__o22ai_2
X_05603_ _09900_/X _05554_/X _05648_/A vssd1 vssd1 vccd1 vccd1 _05641_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08322_ _09998_/S _09999_/S _08322_/C _08413_/B vssd1 vssd1 vccd1 vccd1 _08839_/A
+ sky130_fd_sc_hd__or4b_4
X_05534_ _05534_/A _05534_/B vssd1 vssd1 vccd1 vccd1 _05534_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05465_ _05465_/A vssd1 vssd1 vccd1 vccd1 _05750_/A sky130_fd_sc_hd__clkbuf_2
X_07204_ _07204_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__or2_1
XFILLER_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _08184_/A _08184_/B vssd1 vssd1 vccd1 vccd1 _08184_/Y sky130_fd_sc_hd__nor2_1
X_05396_ _05396_/A _05404_/A vssd1 vssd1 vccd1 vccd1 _05400_/C sky130_fd_sc_hd__or2_1
XFILLER_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ _07123_/A _07123_/B _07202_/A vssd1 vssd1 vccd1 vccd1 _07138_/A sky130_fd_sc_hd__a21o_1
XFILLER_133_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07066_ _06866_/A _07102_/B _07068_/A _07081_/B _07065_/Y vssd1 vssd1 vccd1 vccd1
+ _07067_/B sky130_fd_sc_hd__o41a_1
X_06017_ _06031_/A vssd1 vssd1 vccd1 vccd1 _06017_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_3 _09408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _07737_/X _07750_/Y _07751_/X _07753_/A vssd1 vssd1 vccd1 vccd1 _07968_/X
+ sky130_fd_sc_hd__a31o_1
X_09707_ _06588_/X input40/X _09709_/S vssd1 vssd1 vccd1 vccd1 _09707_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06919_ _06919_/A _06925_/A vssd1 vssd1 vccd1 vccd1 _06919_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07899_ _07896_/X _07898_/X _07896_/X _07898_/X vssd1 vssd1 vccd1 vccd1 _07899_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09638_ _06356_/X _06358_/X _10175_/Q vssd1 vssd1 vccd1 vccd1 _09638_/X sky130_fd_sc_hd__mux2_2
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ _08395_/Y _09568_/X _09600_/S vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__mux2_2
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10413_ _10422_/CLK _10413_/D vssd1 vssd1 vccd1 vccd1 _10413_/Q sky130_fd_sc_hd__dfxtp_1
X_10344_ _10346_/CLK _10344_/D vssd1 vssd1 vccd1 vccd1 _10344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10275_ _10300_/CLK _10275_/D vssd1 vssd1 vccd1 vccd1 _10275_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05250_ _08753_/A _05263_/A input22/X _05264_/A _05245_/X vssd1 vssd1 vccd1 vccd1
+ _10359_/D sky130_fd_sc_hd__o221a_1
X_05181_ _10395_/Q vssd1 vssd1 vccd1 vccd1 _05181_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ _08918_/Y _08939_/X _08918_/Y _08939_/X vssd1 vssd1 vccd1 vccd1 _08940_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_130_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08871_ _10296_/Q _07453_/Y _08842_/Y _08870_/X vssd1 vssd1 vccd1 vccd1 _08871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ _07814_/A _09915_/X _07815_/A _07837_/B _07821_/Y vssd1 vssd1 vccd1 vccd1
+ _07823_/B sky130_fd_sc_hd__o41a_1
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07753_ _07753_/A vssd1 vssd1 vccd1 vccd1 _07753_/Y sky130_fd_sc_hd__inv_2
X_06704_ _06629_/Y _06703_/Y _08715_/A vssd1 vssd1 vccd1 vccd1 _06812_/B sky130_fd_sc_hd__o21a_1
X_07684_ _07684_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07695_/A sky130_fd_sc_hd__or2_2
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06635_ _10364_/Q vssd1 vssd1 vccd1 vccd1 _06635_/Y sky130_fd_sc_hd__inv_2
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__nand2_1
X_09354_ _09354_/A _09452_/B _09354_/C _09354_/D vssd1 vssd1 vccd1 vccd1 _09355_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_52_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _08309_/B vssd1 vssd1 vccd1 vccd1 _08305_/Y sky130_fd_sc_hd__inv_2
X_06566_ _10104_/Q _06465_/A _08439_/A _06436_/A vssd1 vssd1 vccd1 vccd1 _06566_/X
+ sky130_fd_sc_hd__a22o_1
X_09285_ _09285_/A vssd1 vssd1 vccd1 vccd1 _09285_/Y sky130_fd_sc_hd__inv_2
X_06497_ _08392_/A _06496_/X _08399_/A _06496_/X _06484_/B vssd1 vssd1 vccd1 vccd1
+ _06498_/B sky130_fd_sc_hd__o221a_1
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05517_ _09988_/X _09996_/X _05498_/X _05516_/X vssd1 vssd1 vccd1 vccd1 _05574_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08236_ _08578_/A _08236_/B vssd1 vssd1 vccd1 vccd1 _08241_/B sky130_fd_sc_hd__or2_2
X_05448_ _05448_/A vssd1 vssd1 vccd1 vccd1 _05449_/B sky130_fd_sc_hd__inv_2
XFILLER_60_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08167_ _10200_/Q vssd1 vssd1 vccd1 vccd1 _08599_/A sky130_fd_sc_hd__inv_2
XFILLER_176_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07118_ _07118_/A _07118_/B _07118_/C vssd1 vssd1 vccd1 vccd1 _07118_/X sky130_fd_sc_hd__or3_1
X_05379_ _10323_/Q vssd1 vssd1 vccd1 vccd1 _05390_/A sky130_fd_sc_hd__inv_2
XFILLER_173_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08098_ _08083_/X _08098_/B _08098_/C _08098_/D vssd1 vssd1 vccd1 vccd1 _08176_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_109_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07049_ _07046_/X _07048_/Y _07046_/X _07048_/Y vssd1 vssd1 vccd1 vccd1 _07049_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10060_ _10426_/CLK _10060_/D vssd1 vssd1 vccd1 vccd1 _10060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10327_ _10328_/CLK _10327_/D vssd1 vssd1 vccd1 vccd1 _10327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10258_ _10274_/CLK _10258_/D vssd1 vssd1 vccd1 vccd1 _10258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _10426_/CLK _10189_/D vssd1 vssd1 vccd1 vccd1 _10189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06420_ _06420_/A vssd1 vssd1 vccd1 vccd1 _06443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06351_ _06351_/A _10136_/Q vssd1 vssd1 vccd1 vccd1 _06352_/B sky130_fd_sc_hd__nor2_1
XFILLER_187_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09070_ _09070_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _09104_/A sky130_fd_sc_hd__or2_2
X_05302_ _05302_/A _05343_/A vssd1 vssd1 vccd1 vccd1 _05339_/A sky130_fd_sc_hd__or2_1
X_06282_ _10236_/Q _08343_/A _06281_/Y _10129_/Q vssd1 vssd1 vccd1 vccd1 _06283_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05233_ _10369_/Q _05230_/X input33/X _05231_/X _05227_/X vssd1 vssd1 vccd1 vccd1
+ _10369_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__or2_1
XFILLER_190_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05164_ _10399_/Q vssd1 vssd1 vccd1 vccd1 _06616_/D sky130_fd_sc_hd__inv_2
XFILLER_162_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05095_ _05095_/A vssd1 vssd1 vccd1 vccd1 _05095_/X sky130_fd_sc_hd__clkbuf_2
X_09972_ _09971_/X _07878_/C _10000_/S vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08923_ _08923_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__nor2_2
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08854_ _10286_/Q vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__inv_2
X_08785_ _08629_/X _08784_/X _08629_/X _08784_/X vssd1 vssd1 vccd1 vccd1 _08788_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_05997_ _06067_/A vssd1 vssd1 vccd1 vccd1 _06028_/A sky130_fd_sc_hd__clkbuf_4
X_07805_ _09915_/X vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07736_ _07699_/A _07699_/B _07721_/B vssd1 vssd1 vccd1 vccd1 _07737_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__or2_1
XFILLER_197_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _09452_/A _09474_/B _09470_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09406_/X
+ sky130_fd_sc_hd__o22a_1
X_06618_ _06605_/X _06608_/X _06613_/Y _06617_/X vssd1 vssd1 vccd1 vccd1 _06809_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07598_ _07588_/X _07589_/X _07596_/X _07597_/X vssd1 vssd1 vccd1 vccd1 _07598_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06549_ _10101_/Q vssd1 vssd1 vccd1 vccd1 _08432_/A sky130_fd_sc_hd__inv_2
X_09337_ _09336_/A _09336_/B _09457_/A vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09268_ _09268_/A _09268_/B vssd1 vssd1 vccd1 vccd1 _09269_/B sky130_fd_sc_hd__or2_1
XFILLER_138_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08219_ _08264_/A vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__buf_2
XFILLER_138_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ _09252_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10112_ _10334_/CLK _10112_/D vssd1 vssd1 vccd1 vccd1 _10112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10043_ _10442_/CLK _10043_/D vssd1 vssd1 vccd1 vccd1 _10043_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_102_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05920_ _10234_/Q _05910_/A input19/X _05911_/A _05918_/X vssd1 vssd1 vccd1 vccd1
+ _10234_/D sky130_fd_sc_hd__o221a_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05851_ _05871_/A vssd1 vssd1 vccd1 vccd1 _05851_/X sky130_fd_sc_hd__clkbuf_2
X_08570_ _08772_/A _08545_/B _08551_/Y _08568_/X _08569_/Y vssd1 vssd1 vccd1 vccd1
+ _08570_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07521_ _07521_/A vssd1 vssd1 vccd1 vccd1 _07523_/A sky130_fd_sc_hd__inv_2
X_05782_ _07854_/A vssd1 vssd1 vccd1 vccd1 _05782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07452_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__buf_2
XFILLER_179_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06403_ _06399_/X _06400_/X _06399_/X _06400_/X vssd1 vssd1 vccd1 vccd1 _06403_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_07383_ _06942_/A _07235_/B _06942_/C _06824_/X vssd1 vssd1 vccd1 vccd1 _07384_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_210_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09122_ _09122_/A vssd1 vssd1 vccd1 vccd1 _09174_/C sky130_fd_sc_hd__inv_2
X_06334_ _06332_/Y _06333_/X _06332_/Y _06333_/X vssd1 vssd1 vccd1 vccd1 _06334_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_194_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06265_ _06265_/A _06265_/B vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__or2_1
XFILLER_175_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _09053_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09100_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06196_ _06203_/A vssd1 vssd1 vccd1 vccd1 _06196_/X sky130_fd_sc_hd__clkbuf_2
X_05216_ _05240_/A vssd1 vssd1 vccd1 vccd1 _05216_/X sky130_fd_sc_hd__clkbuf_2
X_08004_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__inv_2
X_05147_ _05129_/X _06615_/D _05146_/Y _05138_/X vssd1 vssd1 vccd1 vccd1 _05148_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09955_ _09954_/X _06631_/Y _09982_/S vssd1 vssd1 vccd1 vccd1 _09955_/X sky130_fd_sc_hd__mux2_2
X_05078_ _05189_/A vssd1 vssd1 vccd1 vccd1 _05078_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08906_ _08855_/A _08855_/B _08855_/Y vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09886_ _06825_/Y _06411_/Y _10022_/S vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__mux2_1
X_08837_ _06272_/A _08708_/X _06000_/A _08642_/X _08836_/X vssd1 vssd1 vccd1 vccd1
+ _08837_/X sky130_fd_sc_hd__o221a_1
X_08768_ _08763_/A _08763_/B _08763_/Y vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__a21oi_1
XFILLER_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08699_ _08694_/B _08698_/Y _08688_/X vssd1 vssd1 vccd1 vccd1 _08699_/X sky130_fd_sc_hd__o21ba_1
XFILLER_198_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07719_ _07652_/B _07718_/Y _07652_/B _07718_/Y vssd1 vssd1 vccd1 vccd1 _07719_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_198_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 _09593_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput63 _09581_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _10029_/X vssd1 vssd1 vccd1 vccd1 io_wb_dat_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10026_ _10445_/Q _09543_/X _08344_/Y _09545_/X _09490_/X _09600_/S vssd1 vssd1 vccd1
+ vccd1 _10026_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06050_ _09813_/X _06043_/X _08751_/A _06044_/X _06045_/X vssd1 vssd1 vccd1 vccd1
+ _10190_/D sky130_fd_sc_hd__o221a_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05001_ input13/X input15/X input14/X vssd1 vssd1 vccd1 vccd1 _05775_/A sky130_fd_sc_hd__or3_4
XFILLER_153_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09740_ _06813_/Y _10405_/Q _09745_/S vssd1 vssd1 vccd1 vccd1 _10071_/D sky130_fd_sc_hd__mux2_1
X_06952_ _06943_/X _06947_/X _06950_/X _06951_/X vssd1 vssd1 vccd1 vccd1 _06952_/X
+ sky130_fd_sc_hd__o22a_1
.ends

