* NGSPICE file created from cic_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt cic_block io_adr_i[0] io_adr_i[1] io_cs_i io_dat_i[0] io_dat_i[10] io_dat_i[11]
+ io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[1] io_dat_i[2] io_dat_i[3]
+ io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7] io_dat_i[8] io_dat_i[9] io_dat_o[0]
+ io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13] io_dat_o[14] io_dat_o[15] io_dat_o[1]
+ io_dat_o[2] io_dat_o[3] io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8]
+ io_dat_o[9] io_eo[0] io_eo[10] io_eo[11] io_eo[12] io_eo[13] io_eo[14] io_eo[15]
+ io_eo[16] io_eo[17] io_eo[18] io_eo[19] io_eo[1] io_eo[20] io_eo[21] io_eo[22] io_eo[23]
+ io_eo[24] io_eo[25] io_eo[26] io_eo[27] io_eo[28] io_eo[29] io_eo[2] io_eo[30] io_eo[31]
+ io_eo[32] io_eo[33] io_eo[34] io_eo[35] io_eo[36] io_eo[37] io_eo[38] io_eo[39]
+ io_eo[3] io_eo[40] io_eo[41] io_eo[42] io_eo[43] io_eo[44] io_eo[45] io_eo[46] io_eo[47]
+ io_eo[48] io_eo[49] io_eo[4] io_eo[50] io_eo[51] io_eo[52] io_eo[53] io_eo[54] io_eo[55]
+ io_eo[56] io_eo[57] io_eo[58] io_eo[59] io_eo[5] io_eo[60] io_eo[61] io_eo[62] io_eo[63]
+ io_eo[6] io_eo[7] io_eo[8] io_eo[9] io_i_0_ci io_i_0_in1[0] io_i_0_in1[1] io_i_0_in1[2]
+ io_i_0_in1[3] io_i_0_in1[4] io_i_0_in1[5] io_i_0_in1[6] io_i_0_in1[7] io_i_1_ci
+ io_i_1_in1[0] io_i_1_in1[1] io_i_1_in1[2] io_i_1_in1[3] io_i_1_in1[4] io_i_1_in1[5]
+ io_i_1_in1[6] io_i_1_in1[7] io_i_2_ci io_i_2_in1[0] io_i_2_in1[1] io_i_2_in1[2]
+ io_i_2_in1[3] io_i_2_in1[4] io_i_2_in1[5] io_i_2_in1[6] io_i_2_in1[7] io_i_3_ci
+ io_i_3_in1[0] io_i_3_in1[1] io_i_3_in1[2] io_i_3_in1[3] io_i_3_in1[4] io_i_3_in1[5]
+ io_i_3_in1[6] io_i_3_in1[7] io_i_4_ci io_i_4_in1[0] io_i_4_in1[1] io_i_4_in1[2]
+ io_i_4_in1[3] io_i_4_in1[4] io_i_4_in1[5] io_i_4_in1[6] io_i_4_in1[7] io_i_5_ci
+ io_i_5_in1[0] io_i_5_in1[1] io_i_5_in1[2] io_i_5_in1[3] io_i_5_in1[4] io_i_5_in1[5]
+ io_i_5_in1[6] io_i_5_in1[7] io_i_6_ci io_i_6_in1[0] io_i_6_in1[1] io_i_6_in1[2]
+ io_i_6_in1[3] io_i_6_in1[4] io_i_6_in1[5] io_i_6_in1[6] io_i_6_in1[7] io_i_7_ci
+ io_i_7_in1[0] io_i_7_in1[1] io_i_7_in1[2] io_i_7_in1[3] io_i_7_in1[4] io_i_7_in1[5]
+ io_i_7_in1[6] io_i_7_in1[7] io_o_0_co io_o_0_out[0] io_o_0_out[1] io_o_0_out[2]
+ io_o_0_out[3] io_o_0_out[4] io_o_0_out[5] io_o_0_out[6] io_o_0_out[7] io_o_1_co
+ io_o_1_out[0] io_o_1_out[1] io_o_1_out[2] io_o_1_out[3] io_o_1_out[4] io_o_1_out[5]
+ io_o_1_out[6] io_o_1_out[7] io_o_2_co io_o_2_out[0] io_o_2_out[1] io_o_2_out[2]
+ io_o_2_out[3] io_o_2_out[4] io_o_2_out[5] io_o_2_out[6] io_o_2_out[7] io_o_3_co
+ io_o_3_out[0] io_o_3_out[1] io_o_3_out[2] io_o_3_out[3] io_o_3_out[4] io_o_3_out[5]
+ io_o_3_out[6] io_o_3_out[7] io_o_4_co io_o_4_out[0] io_o_4_out[1] io_o_4_out[2]
+ io_o_4_out[3] io_o_4_out[4] io_o_4_out[5] io_o_4_out[6] io_o_4_out[7] io_o_5_co
+ io_o_5_out[0] io_o_5_out[1] io_o_5_out[2] io_o_5_out[3] io_o_5_out[4] io_o_5_out[5]
+ io_o_5_out[6] io_o_5_out[7] io_o_6_co io_o_6_out[0] io_o_6_out[1] io_o_6_out[2]
+ io_o_6_out[3] io_o_6_out[4] io_o_6_out[5] io_o_6_out[6] io_o_6_out[7] io_o_7_co
+ io_o_7_out[0] io_o_7_out[1] io_o_7_out[2] io_o_7_out[3] io_o_7_out[4] io_o_7_out[5]
+ io_o_7_out[6] io_o_7_out[7] io_vci io_vco io_vi io_we_i io_wo[0] io_wo[10] io_wo[11]
+ io_wo[12] io_wo[13] io_wo[14] io_wo[15] io_wo[16] io_wo[17] io_wo[18] io_wo[19]
+ io_wo[1] io_wo[20] io_wo[21] io_wo[22] io_wo[23] io_wo[24] io_wo[25] io_wo[26] io_wo[27]
+ io_wo[28] io_wo[29] io_wo[2] io_wo[30] io_wo[31] io_wo[32] io_wo[33] io_wo[34] io_wo[35]
+ io_wo[36] io_wo[37] io_wo[38] io_wo[39] io_wo[3] io_wo[40] io_wo[41] io_wo[42] io_wo[43]
+ io_wo[44] io_wo[45] io_wo[46] io_wo[47] io_wo[48] io_wo[49] io_wo[4] io_wo[50] io_wo[51]
+ io_wo[52] io_wo[53] io_wo[54] io_wo[55] io_wo[56] io_wo[57] io_wo[58] io_wo[59]
+ io_wo[5] io_wo[60] io_wo[61] io_wo[62] io_wo[63] io_wo[6] io_wo[7] io_wo[8] io_wo[9]
+ wb_clk_i wb_rst_i vccd1 vssd1
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3155_ _3189_/CLK _3155_/D vssd1 vssd1 vccd1 vccd1 _3155_/Q sky130_fd_sc_hd__dfxtp_4
X_3086_ _3110_/CLK _3086_/D vssd1 vssd1 vccd1 vccd1 _3086_/Q sky130_fd_sc_hd__dfxtp_1
X_2106_ _3047_/Q _2996_/X _2106_/S vssd1 vssd1 vccd1 vccd1 _3047_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2037_ _2034_/Y _2035_/Y _2094_/A vssd1 vssd1 vccd1 vccd1 _2037_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2939_ _2387_/Y _1923_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2939_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2724_ _2727_/X _3140_/Q _3200_/Q vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__mux2_1
X_2655_ _3030_/Q vssd1 vssd1 vccd1 vccd1 _2655_/Y sky130_fd_sc_hd__inv_2
X_1606_ input6/X _1606_/B _2608_/A vssd1 vssd1 vccd1 vccd1 _1606_/Y sky130_fd_sc_hd__nor3_2
X_2586_ _3175_/Q _1544_/B _2582_/Y _2585_/Y vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__a211o_1
X_1537_ input2/X vssd1 vssd1 vccd1 vccd1 _2598_/A sky130_fd_sc_hd__clkbuf_2
X_1468_ _1472_/A _1633_/B vssd1 vssd1 vccd1 vccd1 _1468_/Y sky130_fd_sc_hd__nand2_1
X_3207_ _3209_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_4
X_3138_ _3138_/CLK _3138_/D vssd1 vssd1 vccd1 vccd1 _3138_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3069_ _3211_/CLK _3069_/D vssd1 vssd1 vccd1 vccd1 _3069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2440_ _3079_/Q vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__inv_2
X_2371_ _2371_/A vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2707_ _2707_/A vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__clkbuf_2
Xoutput242 _3041_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput231 _3055_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput220 _3094_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput253 _2673_/X vssd1 vssd1 vccd1 vccd1 io_wo[13] sky130_fd_sc_hd__clkbuf_2
X_2638_ _2646_/A _2981_/X vssd1 vssd1 vccd1 vccd1 _2638_/Y sky130_fd_sc_hd__nand2_1
Xoutput264 _2683_/X vssd1 vssd1 vccd1 vccd1 io_wo[23] sky130_fd_sc_hd__clkbuf_2
Xoutput275 _2693_/X vssd1 vssd1 vccd1 vccd1 io_wo[33] sky130_fd_sc_hd__clkbuf_2
X_2569_ _2600_/A _2600_/B _3156_/Q vssd1 vssd1 vccd1 vccd1 _2569_/Y sky130_fd_sc_hd__nand3_2
Xoutput286 _2703_/X vssd1 vssd1 vccd1 vccd1 io_wo[43] sky130_fd_sc_hd__clkbuf_2
Xoutput297 _2713_/X vssd1 vssd1 vccd1 vccd1 io_wo[53] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_4 _3015_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1940_ _1887_/Y _1882_/X _1886_/Y _2026_/A vssd1 vssd1 vccd1 vccd1 _1940_/Y sky130_fd_sc_hd__o31ai_2
X_1871_ _1868_/X _1869_/Y _1659_/X _1870_/Y vssd1 vssd1 vccd1 vccd1 _3103_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2423_ _2427_/A _2759_/X vssd1 vssd1 vccd1 vccd1 _2423_/Y sky130_fd_sc_hd__nand2_1
X_2354_ _3139_/Q vssd1 vssd1 vccd1 vccd1 _2354_/Y sky130_fd_sc_hd__inv_2
X_2285_ _2285_/A _2285_/B vssd1 vssd1 vccd1 vccd1 _2285_/X sky130_fd_sc_hd__xor2_1
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2070_ _2070_/A _2070_/B vssd1 vssd1 vccd1 vccd1 _2072_/C sky130_fd_sc_hd__nor2_1
XFILLER_75_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _2308_/Y _2307_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1923_ _3092_/Q vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__inv_2
X_1854_ _1862_/S _1851_/X _1853_/X vssd1 vssd1 vccd1 vccd1 _3108_/D sky130_fd_sc_hd__o21bai_1
X_1785_ _1785_/A _1785_/B vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__xor2_1
X_2406_ _3178_/Q vssd1 vssd1 vccd1 vccd1 _2406_/Y sky130_fd_sc_hd__inv_2
X_2337_ _2361_/A _3003_/X vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2268_ _2268_/A vssd1 vssd1 vccd1 vccd1 _2268_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2199_ _2199_/A vssd1 vssd1 vccd1 vccd1 _2253_/C sky130_fd_sc_hd__inv_2
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3171_ _3189_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2122_ _2815_/X vssd1 vssd1 vccd1 vccd1 _2123_/B sky130_fd_sc_hd__inv_2
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _2994_/X _2977_/X vssd1 vssd1 vccd1 vccd1 _2070_/A sky130_fd_sc_hd__nor2_1
X_2955_ _2361_/Y _2954_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__mux2_2
X_2886_ _2457_/Y _2885_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2886_/X sky130_fd_sc_hd__mux2_1
X_1906_ _1920_/A _1906_/B _1920_/B vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__nand3_4
X_1837_ _1831_/Y _1833_/Y _1836_/Y vssd1 vssd1 vccd1 vccd1 _1837_/Y sky130_fd_sc_hd__a21boi_1
X_1768_ _1769_/A _1769_/B _1769_/C vssd1 vssd1 vccd1 vccd1 _1768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1699_ _1699_/A _1699_/B vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__xor2_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput120 io_i_4_ci vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__clkbuf_1
Xinput153 io_i_7_in1[5] vssd1 vssd1 vccd1 vccd1 _2418_/A sky130_fd_sc_hd__buf_1
Xinput131 io_i_5_in1[1] vssd1 vssd1 vccd1 vccd1 _2368_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput142 io_i_6_in1[3] vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__buf_1
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ _2305_/Y _2242_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__mux2_1
X_2671_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__clkbuf_1
X_1622_ _3160_/Q _1613_/X _1583_/X _1621_/Y vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__o211a_1
X_1553_ _3182_/Q _1540_/X _1541_/X _1552_/Y vssd1 vssd1 vccd1 vccd1 _3182_/D sky130_fd_sc_hd__o211a_1
X_1484_ _1535_/B vssd1 vssd1 vccd1 vccd1 _1498_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3154_ _3189_/CLK _3154_/D vssd1 vssd1 vccd1 vccd1 _3154_/Q sky130_fd_sc_hd__dfxtp_4
X_2105_ _3048_/Q _2997_/X _2106_/S vssd1 vssd1 vccd1 vccd1 _3048_/D sky130_fd_sc_hd__mux2_1
X_3085_ _3110_/CLK _3085_/D vssd1 vssd1 vccd1 vccd1 _3085_/Q sky130_fd_sc_hd__dfxtp_1
X_2036_ _2988_/X _2965_/X vssd1 vssd1 vccd1 vccd1 _2094_/A sky130_fd_sc_hd__nor2_4
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ _3007_/A3 _3107_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__mux2_1
X_2869_ input99/X _3020_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2723_ _2723_/A vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__clkbuf_2
X_2654_ _2654_/A _2987_/X vssd1 vssd1 vccd1 vccd1 _2654_/Y sky130_fd_sc_hd__nand2_1
X_1605_ _3165_/Q vssd1 vssd1 vccd1 vccd1 _1605_/Y sky130_fd_sc_hd__inv_2
X_2585_ _2585_/A _2585_/B vssd1 vssd1 vccd1 vccd1 _2585_/Y sky130_fd_sc_hd__nand2_1
X_1536_ _3186_/Q _1522_/A _1525_/X _1535_/Y vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__o211a_1
X_1467_ _1467_/A vssd1 vssd1 vccd1 vccd1 _1633_/B sky130_fd_sc_hd__inv_2
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _3209_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_4
X_3137_ _3138_/CLK _3137_/D vssd1 vssd1 vccd1 vccd1 _3137_/Q sky130_fd_sc_hd__dfxtp_2
X_3068_ _3209_/CLK _3068_/D vssd1 vssd1 vccd1 vccd1 _3068_/Q sky130_fd_sc_hd__dfxtp_1
X_2019_ _2019_/A vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2370_ _3048_/Q vssd1 vssd1 vccd1 vccd1 _2370_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3211_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _2706_/A vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__clkbuf_2
Xoutput210 _3109_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[6] sky130_fd_sc_hd__clkbuf_2
X_2637_ _3184_/Q vssd1 vssd1 vccd1 vccd1 _2637_/Y sky130_fd_sc_hd__inv_2
Xoutput232 _3056_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput221 _2535_/Y vssd1 vssd1 vccd1 vccd1 io_o_5_co sky130_fd_sc_hd__clkbuf_2
Xoutput243 _3042_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput254 _2674_/X vssd1 vssd1 vccd1 vccd1 io_wo[14] sky130_fd_sc_hd__clkbuf_2
Xoutput265 _2684_/X vssd1 vssd1 vccd1 vccd1 io_wo[24] sky130_fd_sc_hd__clkbuf_2
Xoutput276 _2694_/X vssd1 vssd1 vccd1 vccd1 io_wo[34] sky130_fd_sc_hd__clkbuf_2
X_2568_ _3204_/Q _2610_/B _2626_/C vssd1 vssd1 vccd1 vccd1 _2568_/Y sky130_fd_sc_hd__nand3_2
Xoutput298 _2714_/X vssd1 vssd1 vccd1 vccd1 io_wo[54] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_5 _3016_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2499_ _3134_/Q vssd1 vssd1 vccd1 vccd1 _2499_/Y sky130_fd_sc_hd__inv_2
Xoutput287 _2704_/X vssd1 vssd1 vccd1 vccd1 io_wo[44] sky130_fd_sc_hd__clkbuf_2
X_1519_ _1535_/B vssd1 vssd1 vccd1 vccd1 _1530_/B sky130_fd_sc_hd__buf_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ _3103_/Q vssd1 vssd1 vccd1 vccd1 _1870_/Y sky130_fd_sc_hd__inv_2
X_2422_ _2422_/A vssd1 vssd1 vccd1 vccd1 _2422_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2353_ _3107_/Q vssd1 vssd1 vccd1 vccd1 _2353_/Y sky130_fd_sc_hd__inv_2
X_2284_ _2284_/A _2284_/B vssd1 vssd1 vccd1 vccd1 _2285_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1999_ _3000_/X _2957_/X _1998_/Y vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__o21a_1
XFILLER_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ _2313_/Y _2970_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__mux2_2
X_1922_ _1670_/X _1917_/Y _1921_/Y vssd1 vssd1 vccd1 vccd1 _3093_/D sky130_fd_sc_hd__o21ai_1
X_1853_ _1955_/S _3108_/Q vssd1 vssd1 vccd1 vccd1 _1853_/X sky130_fd_sc_hd__and2b_1
X_1784_ _1783_/Y _3122_/Q _1786_/S vssd1 vssd1 vccd1 vccd1 _3122_/D sky130_fd_sc_hd__mux2_1
X_2405_ _3063_/Q vssd1 vssd1 vccd1 vccd1 _2405_/Y sky130_fd_sc_hd__inv_2
X_2336_ _2372_/A vssd1 vssd1 vccd1 vccd1 _2361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2267_ _2267_/A _2289_/A vssd1 vssd1 vccd1 vccd1 _2268_/A sky130_fd_sc_hd__and2_1
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2198_ _3010_/X _2839_/X vssd1 vssd1 vccd1 vccd1 _2199_/A sky130_fd_sc_hd__and2b_1
XFILLER_37_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3170_ _3189_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
X_2121_ _2982_/X vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__inv_2
XFILLER_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2052_ _2082_/B _2082_/A _2078_/A vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__nand3_4
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2954_ _2362_/Y _2309_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2954_/X sky130_fd_sc_hd__mux2_1
X_2885_ _2458_/Y _2312_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__mux2_1
X_1905_ _1905_/A _1905_/B vssd1 vssd1 vccd1 vccd1 _1920_/B sky130_fd_sc_hd__nor2_4
X_1836_ _1836_/A _2526_/A vssd1 vssd1 vccd1 vccd1 _1836_/Y sky130_fd_sc_hd__nor2_1
X_1767_ _1767_/A _1767_/B vssd1 vssd1 vccd1 vccd1 _1769_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1698_ _1697_/Y _3138_/Q _2290_/S vssd1 vssd1 vccd1 vccd1 _3138_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2319_ _3121_/Q vssd1 vssd1 vccd1 vccd1 _2319_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput110 io_i_2_in1[7] vssd1 vssd1 vccd1 vccd1 _2899_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput154 io_i_7_in1[6] vssd1 vssd1 vccd1 vccd1 _2414_/A sky130_fd_sc_hd__buf_1
Xinput132 io_i_5_in1[2] vssd1 vssd1 vccd1 vccd1 _2363_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput121 io_i_4_in1[0] vssd1 vssd1 vccd1 vccd1 _3011_/A3 sky130_fd_sc_hd__buf_1
Xinput143 io_i_6_in1[4] vssd1 vssd1 vccd1 vccd1 _2303_/A sky130_fd_sc_hd__buf_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2670_ _2670_/A vssd1 vssd1 vccd1 vccd1 _2670_/X sky130_fd_sc_hd__clkbuf_1
X_1621_ _1627_/A _1621_/B vssd1 vssd1 vccd1 vccd1 _1621_/Y sky130_fd_sc_hd__nand2_1
X_1552_ _1551_/X _1558_/B _1648_/B vssd1 vssd1 vccd1 vccd1 _1552_/Y sky130_fd_sc_hd__nand3b_1
X_1483_ _2596_/A _2611_/A vssd1 vssd1 vccd1 vccd1 _1535_/B sky130_fd_sc_hd__nor2b_4
X_3153_ _3211_/CLK _3153_/D vssd1 vssd1 vccd1 vccd1 _3153_/Q sky130_fd_sc_hd__dfxtp_4
X_2104_ _3049_/Q _2998_/X _2106_/S vssd1 vssd1 vccd1 vccd1 _3049_/D sky130_fd_sc_hd__mux2_1
X_3084_ _3110_/CLK _3084_/D vssd1 vssd1 vccd1 vccd1 _3084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2035_ _2823_/X vssd1 vssd1 vccd1 vccd1 _2035_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2937_ _2389_/Y _2936_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2937_/X sky130_fd_sc_hd__mux2_4
X_2868_ _2478_/Y _2867_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__mux2_1
X_1819_ _2427_/B _2910_/X _2755_/X _2907_/X vssd1 vssd1 vccd1 vccd1 _1819_/X sky130_fd_sc_hd__a211o_1
X_2799_ _2474_/Y _2798_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2799_/X sky130_fd_sc_hd__mux2_2
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2722_ _2722_/A vssd1 vssd1 vccd1 vccd1 _2722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653_ _3029_/Q vssd1 vssd1 vccd1 vccd1 _2653_/Y sky130_fd_sc_hd__inv_2
X_1604_ _1587_/X _1602_/Y _1655_/A _1603_/Y vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__a211oi_1
X_2584_ _3207_/Q _2627_/B _2593_/C vssd1 vssd1 vccd1 vccd1 _2585_/B sky130_fd_sc_hd__nand3_1
X_1535_ _1532_/X _1535_/B _1636_/B vssd1 vssd1 vccd1 vccd1 _1535_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1466_ _2493_/A _1458_/X _1459_/X _1465_/Y vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__o211a_1
X_3205_ _3205_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3136_ _3138_/CLK _3136_/D vssd1 vssd1 vccd1 vccd1 _3136_/Q sky130_fd_sc_hd__dfxtp_2
X_3067_ _3123_/CLK _3067_/D vssd1 vssd1 vccd1 vccd1 _3067_/Q sky130_fd_sc_hd__dfxtp_1
X_2018_ _3071_/Q vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2705_ _2705_/A vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__clkbuf_2
Xoutput200 _3124_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[5] sky130_fd_sc_hd__clkbuf_2
X_2636_ _3023_/Q vssd1 vssd1 vccd1 vccd1 _2636_/Y sky130_fd_sc_hd__inv_2
Xoutput233 _3057_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput222 _3071_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput244 _3043_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput211 _3110_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput255 _2675_/X vssd1 vssd1 vccd1 vccd1 io_wo[15] sky130_fd_sc_hd__clkbuf_2
Xoutput266 _2685_/X vssd1 vssd1 vccd1 vccd1 io_wo[25] sky130_fd_sc_hd__clkbuf_2
Xoutput277 _2695_/X vssd1 vssd1 vccd1 vccd1 io_wo[35] sky130_fd_sc_hd__clkbuf_2
X_2567_ _2605_/C vssd1 vssd1 vccd1 vccd1 _2610_/B sky130_fd_sc_hd__buf_2
Xoutput299 _2715_/X vssd1 vssd1 vccd1 vccd1 io_wo[55] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2498_ _2498_/A _2506_/B vssd1 vssd1 vccd1 vccd1 _2498_/Y sky130_fd_sc_hd__nand2_1
Xoutput288 _2705_/X vssd1 vssd1 vccd1 vccd1 io_wo[45] sky130_fd_sc_hd__clkbuf_2
X_1518_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__buf_1
X_1449_ _2439_/A _1435_/X _1438_/X _1448_/Y vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3119_ _3123_/CLK _3119_/D vssd1 vssd1 vccd1 vccd1 _3119_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2421_ _2914_/X vssd1 vssd1 vccd1 vccd1 _2421_/Y sky130_fd_sc_hd__inv_2
X_2352_ _2352_/A vssd1 vssd1 vccd1 vccd1 _2352_/Y sky130_fd_sc_hd__inv_2
X_2283_ _1796_/S _2263_/Y _2282_/Y vssd1 vssd1 vccd1 vccd1 _3014_/D sky130_fd_sc_hd__o21ai_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1998_ _1998_/A _1998_/B vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__nand2_1
X_2619_ _3150_/Q _2627_/B _2627_/C vssd1 vssd1 vccd1 vccd1 _2619_/Y sky130_fd_sc_hd__nand3_2
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _2315_/Y _2314_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__mux2_1
X_1921_ _1919_/Y _1920_/X _1937_/S vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__o21bai_1
X_1852_ _2749_/X vssd1 vssd1 vccd1 vccd1 _1955_/S sky130_fd_sc_hd__clkbuf_2
X_1783_ _1783_/A _1783_/B vssd1 vssd1 vccd1 vccd1 _1783_/Y sky130_fd_sc_hd__xnor2_1
X_2404_ _2404_/A _2733_/X vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__nand2_1
X_2335_ _2348_/A _3186_/Q vssd1 vssd1 vccd1 vccd1 _2335_/Y sky130_fd_sc_hd__nand2_1
X_2266_ _2266_/A _2266_/B vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2197_ _2835_/X _2257_/A _2196_/Y vssd1 vssd1 vccd1 vccd1 _2253_/B sky130_fd_sc_hd__o21ai_2
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2120_ _2114_/X _2118_/Y _2119_/Y vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__o21bai_4
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2051_ _2056_/A _2051_/B vssd1 vssd1 vccd1 vccd1 _2078_/A sky130_fd_sc_hd__nor2_4
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _2366_/Y _2952_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__mux2_2
X_1904_ _2743_/X _2940_/X _2741_/X _2937_/X vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__a211oi_4
X_2884_ _2884_/A0 _3137_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__mux2_1
X_1835_ _2765_/X _2922_/X vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__and2_1
X_1766_ _3125_/Q vssd1 vssd1 vccd1 vccd1 _1766_/Y sky130_fd_sc_hd__inv_2
X_1697_ _1697_/A _1697_/B vssd1 vssd1 vccd1 vccd1 _1697_/Y sky130_fd_sc_hd__xnor2_1
X_2318_ _3089_/Q vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2249_ _2249_/A _2249_/B vssd1 vssd1 vccd1 vccd1 _2249_/X sky130_fd_sc_hd__xor2_1
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput111 io_i_3_ci vssd1 vssd1 vccd1 vccd1 _2442_/A sky130_fd_sc_hd__buf_1
Xinput100 io_i_1_in1[6] vssd1 vssd1 vccd1 vccd1 _2872_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput122 io_i_4_in1[1] vssd1 vssd1 vccd1 vccd1 _3010_/A3 sky130_fd_sc_hd__buf_1
Xinput133 io_i_5_in1[3] vssd1 vssd1 vccd1 vccd1 _2358_/A sky130_fd_sc_hd__clkbuf_1
Xinput144 io_i_6_in1[5] vssd1 vssd1 vccd1 vccd1 _2299_/A sky130_fd_sc_hd__buf_1
Xinput155 io_i_7_in1[7] vssd1 vssd1 vccd1 vccd1 _2409_/A sky130_fd_sc_hd__buf_1
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1620_ _3161_/Q _1613_/X _1583_/X _1619_/Y vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__o211a_1
X_1551_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__buf_1
X_1482_ input2/X vssd1 vssd1 vccd1 vccd1 _2611_/A sky130_fd_sc_hd__clkbuf_2
X_3152_ _3211_/CLK _3152_/D vssd1 vssd1 vccd1 vccd1 _3152_/Q sky130_fd_sc_hd__dfxtp_4
X_2103_ _3050_/Q _2361_/B _2106_/S vssd1 vssd1 vccd1 vccd1 _3050_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _3122_/CLK _3083_/D vssd1 vssd1 vccd1 vccd1 _3083_/Q sky130_fd_sc_hd__dfxtp_1
X_2034_ _2988_/X _2965_/X vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__nand2_2
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2936_ _2390_/Y _2304_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2867_ _2479_/Y _2347_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__mux2_1
X_1818_ _1818_/A _1818_/B vssd1 vssd1 vccd1 vccd1 _1859_/A sky130_fd_sc_hd__nor2_2
X_2798_ _2414_/Y _2339_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2798_/X sky130_fd_sc_hd__mux2_1
X_1749_ _1779_/B _1779_/A _1775_/A vssd1 vssd1 vccd1 vccd1 _1769_/A sky130_fd_sc_hd__nand3_4
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2721_ _2721_/A vssd1 vssd1 vccd1 vccd1 _2721_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2652_ _2654_/A _2986_/X vssd1 vssd1 vccd1 vccd1 _2652_/Y sky130_fd_sc_hd__nand2_1
X_1603_ input7/X _1606_/B _1603_/C vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__nor3_1
X_2583_ _2548_/A _3191_/Q _2631_/C vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__nand3b_1
X_1534_ _3187_/Q _1522_/X _1525_/X _1533_/Y vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__o211a_1
X_1465_ _1472_/A _1631_/B vssd1 vssd1 vccd1 vccd1 _1465_/Y sky130_fd_sc_hd__nand2_1
X_3204_ _3205_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_4
X_3135_ _3138_/CLK _3135_/D vssd1 vssd1 vccd1 vccd1 _3135_/Q sky130_fd_sc_hd__dfxtp_2
X_3066_ _3123_/CLK _3066_/D vssd1 vssd1 vccd1 vccd1 _3066_/Q sky130_fd_sc_hd__dfxtp_1
X_2017_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2102_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2919_ _2415_/Y _2918_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _2704_/A vssd1 vssd1 vccd1 vccd1 _2704_/X sky130_fd_sc_hd__clkbuf_2
Xoutput201 _3125_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[6] sky130_fd_sc_hd__clkbuf_2
X_2635_ _2646_/A _2980_/X vssd1 vssd1 vccd1 vccd1 _2635_/Y sky130_fd_sc_hd__nand2_1
Xoutput223 _3072_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput212 _2536_/Y vssd1 vssd1 vccd1 vccd1 io_o_4_co sky130_fd_sc_hd__clkbuf_2
Xoutput234 _3058_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput245 _3044_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput256 _2676_/X vssd1 vssd1 vccd1 vccd1 io_wo[16] sky130_fd_sc_hd__clkbuf_2
Xoutput267 _2686_/X vssd1 vssd1 vccd1 vccd1 io_wo[26] sky130_fd_sc_hd__clkbuf_2
X_2566_ _2593_/B _3188_/Q _2632_/C vssd1 vssd1 vccd1 vccd1 _2566_/Y sky130_fd_sc_hd__nand3b_4
X_1517_ _3193_/Q _1506_/X _1510_/X _1516_/Y vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__o211a_1
X_2497_ _3202_/Q vssd1 vssd1 vccd1 vccd1 _2506_/B sky130_fd_sc_hd__clkbuf_2
Xoutput278 _2696_/X vssd1 vssd1 vccd1 vccd1 io_wo[36] sky130_fd_sc_hd__clkbuf_2
Xoutput289 _2706_/X vssd1 vssd1 vccd1 vccd1 io_wo[46] sky130_fd_sc_hd__clkbuf_2
X_1448_ _1451_/A _1621_/B vssd1 vssd1 vccd1 vccd1 _1448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3118_ _3205_/CLK _3118_/D vssd1 vssd1 vccd1 vccd1 _3118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3049_ _3110_/CLK _3049_/D vssd1 vssd1 vccd1 vccd1 _3049_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2420_ _3084_/Q vssd1 vssd1 vccd1 vccd1 _2420_/Y sky130_fd_sc_hd__inv_2
X_2351_ _3052_/Q vssd1 vssd1 vccd1 vccd1 _2351_/Y sky130_fd_sc_hd__inv_2
X_2282_ _2280_/Y _2281_/X _1693_/A vssd1 vssd1 vccd1 vccd1 _2282_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _1657_/X _1992_/Y _1996_/Y vssd1 vssd1 vccd1 vccd1 _3077_/D sky130_fd_sc_hd__o21ai_1
X_2618_ _2596_/X _3198_/Q _2618_/C vssd1 vssd1 vccd1 vccd1 _2618_/Y sky130_fd_sc_hd__nand3b_4
X_2549_ _2598_/A vssd1 vssd1 vccd1 vccd1 _2626_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1920_ _1920_/A _1920_/B _1920_/C vssd1 vssd1 vccd1 vccd1 _1920_/X sky130_fd_sc_hd__and3_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1851_ _1851_/A _1851_/B vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__xor2_1
X_1782_ _1785_/B _1785_/A _1781_/Y vssd1 vssd1 vccd1 vccd1 _1783_/B sky130_fd_sc_hd__a21oi_1
X_2403_ _2926_/X vssd1 vssd1 vccd1 vccd1 _2403_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2334_ _2348_/A _3188_/Q vssd1 vssd1 vccd1 vccd1 _2334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2265_ _2797_/X _2868_/X vssd1 vssd1 vccd1 vccd1 _2266_/B sky130_fd_sc_hd__and2_1
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2196_ _2837_/X _3011_/X vssd1 vssd1 vccd1 vccd1 _2196_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2050_ _2993_/X _2975_/X vssd1 vssd1 vccd1 vccd1 _2051_/B sky130_fd_sc_hd__and2_1
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2952_ _2367_/Y _2316_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2952_/X sky130_fd_sc_hd__mux2_1
X_1903_ _1918_/A vssd1 vssd1 vccd1 vccd1 _1906_/B sky130_fd_sc_hd__inv_2
X_2883_ _2460_/Y _2882_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2883_/X sky130_fd_sc_hd__mux2_2
X_1834_ _2765_/X _2922_/X vssd1 vssd1 vccd1 vccd1 _1836_/A sky130_fd_sc_hd__nor2_4
X_1765_ _1661_/X _1729_/Y _1764_/Y vssd1 vssd1 vccd1 vccd1 _3126_/D sky130_fd_sc_hd__o21ai_1
X_1696_ _1699_/B _1699_/A _1695_/Y vssd1 vssd1 vccd1 vccd1 _1697_/B sky130_fd_sc_hd__a21oi_1
X_2317_ _2317_/A vssd1 vssd1 vccd1 vccd1 _2317_/Y sky130_fd_sc_hd__inv_2
X_2248_ _2508_/A _2841_/X _2247_/Y vssd1 vssd1 vccd1 vccd1 _2249_/B sky130_fd_sc_hd__o21bai_1
X_2179_ _3035_/Q _2992_/X _2183_/S vssd1 vssd1 vccd1 vccd1 _3035_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput101 io_i_1_in1[7] vssd1 vssd1 vccd1 vccd1 _2875_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput123 io_i_4_in1[2] vssd1 vssd1 vccd1 vccd1 _3009_/A3 sky130_fd_sc_hd__buf_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput112 io_i_3_in1[0] vssd1 vssd1 vccd1 vccd1 _2902_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput145 io_i_6_in1[6] vssd1 vssd1 vccd1 vccd1 _2295_/A sky130_fd_sc_hd__buf_1
Xinput134 io_i_5_in1[4] vssd1 vssd1 vccd1 vccd1 _2352_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput156 io_vci vssd1 vssd1 vccd1 vccd1 _2802_/A0 sky130_fd_sc_hd__buf_2
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _3183_/Q _1540_/X _1541_/X _1549_/Y vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3209_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1481_ input1/X vssd1 vssd1 vccd1 vccd1 _2596_/A sky130_fd_sc_hd__clkbuf_2
X_3151_ _3211_/CLK _3151_/D vssd1 vssd1 vccd1 vccd1 _3151_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2102_ _3051_/Q _3000_/X _2102_/S vssd1 vssd1 vccd1 vccd1 _3051_/D sky130_fd_sc_hd__mux2_1
X_3082_ _3122_/CLK _3082_/D vssd1 vssd1 vccd1 vccd1 _3082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2033_ _2989_/X _2967_/X vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__and2_2
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _3008_/A3 _3106_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2935_/X sky130_fd_sc_hd__mux2_1
X_2866_ input98/X _3019_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__mux2_1
X_1817_ _2757_/X _2910_/X vssd1 vssd1 vccd1 vccd1 _1818_/B sky130_fd_sc_hd__and2_1
X_2797_ _2477_/Y _2796_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__mux2_1
X_1748_ _1753_/A _1748_/B vssd1 vssd1 vccd1 vccd1 _1775_/A sky130_fd_sc_hd__nor2_4
X_1679_ _2787_/X _2853_/X vssd1 vssd1 vccd1 vccd1 _1679_/Y sky130_fd_sc_hd__nor2_4
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _2720_/A vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2651_ _3044_/Q vssd1 vssd1 vccd1 vccd1 _2651_/Y sky130_fd_sc_hd__inv_2
X_1602_ _3166_/Q vssd1 vssd1 vccd1 vccd1 _1602_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2582_ _2620_/C _2616_/C _3159_/Q vssd1 vssd1 vccd1 vccd1 _2582_/Y sky130_fd_sc_hd__nor3b_2
X_1533_ _1532_/X _1535_/B _1633_/B vssd1 vssd1 vccd1 vccd1 _1533_/Y sky130_fd_sc_hd__nand3b_1
X_1464_ _1464_/A vssd1 vssd1 vccd1 vccd1 _1631_/B sky130_fd_sc_hd__clkinv_4
X_3203_ _3205_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3134_ _3205_/CLK _3134_/D vssd1 vssd1 vccd1 vccd1 _3134_/Q sky130_fd_sc_hd__dfxtp_1
X_3065_ _3123_/CLK _3065_/D vssd1 vssd1 vccd1 vccd1 _3065_/Q sky130_fd_sc_hd__dfxtp_1
X_2016_ _1657_/X _2012_/Y _2013_/X _2015_/Y vssd1 vssd1 vccd1 vccd1 _3072_/D sky130_fd_sc_hd__o22ai_1
X_2918_ _2416_/Y _1842_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2918_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2849_ _2500_/Y _2848_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2703_ _2703_/A vssd1 vssd1 vccd1 vccd1 _2703_/X sky130_fd_sc_hd__clkbuf_1
X_2634_ _2654_/A vssd1 vssd1 vccd1 vccd1 _2646_/A sky130_fd_sc_hd__buf_2
Xoutput224 _3073_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput213 _3087_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput235 _3059_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput202 _3126_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[7] sky130_fd_sc_hd__clkbuf_2
X_2565_ _3171_/Q _1544_/B _2558_/Y _2564_/Y vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__a211o_1
Xoutput246 _3045_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput257 _2677_/X vssd1 vssd1 vccd1 vccd1 io_wo[17] sky130_fd_sc_hd__clkbuf_2
Xoutput268 _2687_/X vssd1 vssd1 vccd1 vccd1 io_wo[27] sky130_fd_sc_hd__clkbuf_2
X_1516_ _1501_/X _1516_/B _1619_/B vssd1 vssd1 vccd1 vccd1 _1516_/Y sky130_fd_sc_hd__nand3b_1
X_2496_ _2496_/A vssd1 vssd1 vccd1 vccd1 _2496_/Y sky130_fd_sc_hd__inv_2
Xoutput279 _2697_/X vssd1 vssd1 vccd1 vccd1 io_wo[37] sky130_fd_sc_hd__clkbuf_2
X_1447_ _1447_/A vssd1 vssd1 vccd1 vccd1 _1621_/B sky130_fd_sc_hd__inv_2
X_3117_ _3139_/CLK _3117_/D vssd1 vssd1 vccd1 vccd1 _3117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3048_ _3110_/CLK _3048_/D vssd1 vssd1 vccd1 vccd1 _3048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2350_ _2361_/A _3001_/X vssd1 vssd1 vccd1 vccd1 _2350_/Y sky130_fd_sc_hd__nand2_1
X_2281_ _2799_/X _2871_/X _2279_/Y _2521_/A vssd1 vssd1 vccd1 vccd1 _2281_/X sky130_fd_sc_hd__o211a_1
XFILLER_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _1994_/Y _1995_/X _2011_/S vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__o21bai_1
X_2617_ _1605_/Y _2608_/X _2614_/Y _2615_/Y _2616_/Y vssd1 vssd1 vccd1 vccd1 _2617_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_2548_ _2548_/A vssd1 vssd1 vccd1 vccd1 _2630_/C sky130_fd_sc_hd__clkbuf_4
X_2479_ _3116_/Q vssd1 vssd1 vccd1 vccd1 _2479_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3193_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1850_ _1855_/B _1855_/A _1849_/Y vssd1 vssd1 vccd1 vccd1 _1851_/B sky130_fd_sc_hd__a21oi_1
X_1781_ _2773_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _1781_/Y sky130_fd_sc_hd__nor2_1
X_2402_ _3064_/Q vssd1 vssd1 vccd1 vccd1 _2402_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2333_ _2541_/A vssd1 vssd1 vccd1 vccd1 _2348_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2264_ _2478_/B _2868_/X vssd1 vssd1 vccd1 vccd1 _2266_/A sky130_fd_sc_hd__nor2_1
X_2195_ _3011_/X _2837_/X vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__and2b_1
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1979_ _3001_/X _2959_/X _3000_/X _2957_/X vssd1 vssd1 vccd1 vccd1 _1980_/B sky130_fd_sc_hd__a211oi_4
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2951_ _2369_/Y _2950_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__mux2_1
X_1902_ _2745_/X _2943_/X vssd1 vssd1 vccd1 vccd1 _1918_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2882_ _2461_/Y _2319_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2882_/X sky130_fd_sc_hd__mux2_1
X_1833_ _1843_/B vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__inv_2
X_1764_ _1760_/Y _1761_/X _1786_/S vssd1 vssd1 vccd1 vccd1 _1764_/Y sky130_fd_sc_hd__o21bai_1
X_1695_ _2791_/X _2859_/X vssd1 vssd1 vccd1 vccd1 _1695_/Y sky130_fd_sc_hd__nor2_1
X_2316_ _3073_/Q vssd1 vssd1 vccd1 vccd1 _2316_/Y sky130_fd_sc_hd__inv_2
X_2247_ _2251_/A _2251_/B vssd1 vssd1 vccd1 vccd1 _2247_/Y sky130_fd_sc_hd__nor2_1
X_2178_ _2727_/X vssd1 vssd1 vccd1 vccd1 _2183_/S sky130_fd_sc_hd__buf_2
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 io_i_2_ci vssd1 vssd1 vccd1 vccd1 _2469_/A sky130_fd_sc_hd__clkbuf_1
Xinput113 io_i_3_in1[1] vssd1 vssd1 vccd1 vccd1 _2905_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput124 io_i_4_in1[3] vssd1 vssd1 vccd1 vccd1 _3008_/A3 sky130_fd_sc_hd__buf_1
Xinput135 io_i_5_in1[5] vssd1 vssd1 vccd1 vccd1 _2345_/A sky130_fd_sc_hd__clkbuf_1
Xinput157 io_vi vssd1 vssd1 vccd1 vccd1 _2332_/A sky130_fd_sc_hd__buf_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput146 io_i_6_in1[7] vssd1 vssd1 vccd1 vccd1 _2291_/A sky130_fd_sc_hd__buf_1
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1611_/C vssd1 vssd1 vccd1 vccd1 _1609_/B sky130_fd_sc_hd__buf_1
X_3150_ _3166_/CLK _3150_/D vssd1 vssd1 vccd1 vccd1 _3150_/Q sky130_fd_sc_hd__dfxtp_4
X_3081_ _3122_/CLK _3081_/D vssd1 vssd1 vccd1 vccd1 _3081_/Q sky130_fd_sc_hd__dfxtp_1
X_2101_ _3052_/Q _3001_/X _2102_/S vssd1 vssd1 vccd1 vccd1 _3052_/D sky130_fd_sc_hd__mux2_1
X_2032_ _3062_/Q vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2934_ _2393_/Y _2933_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__mux2_2
X_2865_ _2481_/Y _2864_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__mux2_2
X_1816_ _2427_/B _2910_/X vssd1 vssd1 vccd1 vccd1 _1818_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2796_ _2418_/Y _2345_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2796_/X sky130_fd_sc_hd__mux2_1
X_1747_ _2779_/X _2892_/X vssd1 vssd1 vccd1 vccd1 _1748_/B sky130_fd_sc_hd__and2_1
X_1678_ _2833_/X vssd1 vssd1 vccd1 vccd1 _1678_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2650_ _3028_/Q vssd1 vssd1 vccd1 vccd1 _2650_/Y sky130_fd_sc_hd__inv_2
X_1601_ _1587_/X _1598_/Y _1655_/A _1600_/Y vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__a211oi_1
X_2581_ _2603_/B vssd1 vssd1 vccd1 vccd1 _2620_/C sky130_fd_sc_hd__buf_2
X_1532_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1532_/X sky130_fd_sc_hd__buf_1
X_1463_ _3204_/Q vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__buf_2
X_3202_ _3205_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3133_ _3205_/CLK _3133_/D vssd1 vssd1 vccd1 vccd1 _3133_/Q sky130_fd_sc_hd__dfxtp_1
X_3064_ _3123_/CLK _3064_/D vssd1 vssd1 vccd1 vccd1 _3064_/Q sky130_fd_sc_hd__dfxtp_1
X_2015_ _1962_/Y _1957_/X _1961_/Y _2106_/S vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _2917_/A0 _3124_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2917_/X sky130_fd_sc_hd__mux2_1
X_2848_ _2501_/Y _2382_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__mux2_1
X_2779_ _2450_/Y _2778_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__mux2_4
XFILLER_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _2702_/A vssd1 vssd1 vccd1 vccd1 _2702_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2633_ _1588_/Y _1603_/C _2630_/Y _2631_/Y _2632_/Y vssd1 vssd1 vccd1 vccd1 _2633_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput214 _3088_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput203 _2537_/Y vssd1 vssd1 vccd1 vccd1 io_o_3_co sky130_fd_sc_hd__clkbuf_2
Xoutput225 _3074_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[3] sky130_fd_sc_hd__clkbuf_2
X_2564_ _2564_/A _2564_/B vssd1 vssd1 vccd1 vccd1 _2564_/Y sky130_fd_sc_hd__nand2_1
X_1515_ _3194_/Q _1506_/X _1510_/X _1514_/Y vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__o211a_1
Xoutput236 _3060_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput247 _3046_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput258 _2678_/X vssd1 vssd1 vccd1 vccd1 io_wo[18] sky130_fd_sc_hd__clkbuf_2
X_2495_ _3172_/Q vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__inv_2
Xoutput269 _2688_/X vssd1 vssd1 vccd1 vccd1 io_wo[28] sky130_fd_sc_hd__clkbuf_2
X_1446_ _3208_/Q vssd1 vssd1 vccd1 vccd1 _2439_/A sky130_fd_sc_hd__buf_2
X_3116_ _3139_/CLK _3116_/D vssd1 vssd1 vccd1 vccd1 _3116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _3110_/CLK _3047_/D vssd1 vssd1 vccd1 vccd1 _3047_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2280_ _2521_/A _2521_/B _2279_/Y vssd1 vssd1 vccd1 vccd1 _2280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _1995_/A _1995_/B _1995_/C vssd1 vssd1 vccd1 vccd1 _1995_/X sky130_fd_sc_hd__and3_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2616_ _3153_/Q _2632_/B _2616_/C vssd1 vssd1 vccd1 vccd1 _2616_/Y sky130_fd_sc_hd__nand3_2
X_2547_ _2596_/A vssd1 vssd1 vccd1 vccd1 _2548_/A sky130_fd_sc_hd__buf_1
X_2478_ _2484_/A _2478_/B vssd1 vssd1 vccd1 vccd1 _2478_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1780_ _1779_/X _3123_/Q _1786_/S vssd1 vssd1 vccd1 vccd1 _3123_/D sky130_fd_sc_hd__mux2_1
X_2401_ _2404_/A _2735_/X vssd1 vssd1 vccd1 vccd1 _2401_/Y sky130_fd_sc_hd__nand2_1
X_2332_ _2332_/A vssd1 vssd1 vccd1 vccd1 _2541_/A sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2263_ _3014_/Q vssd1 vssd1 vccd1 vccd1 _2263_/Y sky130_fd_sc_hd__inv_2
X_2194_ _2194_/A vssd1 vssd1 vccd1 vccd1 _2251_/A sky130_fd_sc_hd__inv_2
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1978_ _1993_/A vssd1 vssd1 vccd1 vccd1 _1981_/B sky130_fd_sc_hd__inv_2
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2950_ _2370_/Y _2012_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__mux2_1
X_2881_ _2881_/A0 _3136_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2881_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1901_ _1930_/B _1930_/A _1926_/A vssd1 vssd1 vccd1 vccd1 _1920_/A sky130_fd_sc_hd__nand3_4
X_1832_ _2763_/X _2919_/X vssd1 vssd1 vccd1 vccd1 _1843_/B sky130_fd_sc_hd__and2_1
X_1763_ _1763_/A vssd1 vssd1 vccd1 vccd1 _1786_/S sky130_fd_sc_hd__buf_2
X_1694_ _1691_/X _3139_/Q _2290_/S vssd1 vssd1 vccd1 vccd1 _3139_/D sky130_fd_sc_hd__mux2_1
X_2315_ _3034_/Q vssd1 vssd1 vccd1 vccd1 _2315_/Y sky130_fd_sc_hd__inv_2
X_2246_ _3008_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _2249_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2177_ _3036_/Q _2993_/X _2177_/S vssd1 vssd1 vccd1 vccd1 _3036_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput114 io_i_3_in1[2] vssd1 vssd1 vccd1 vccd1 _2908_/A0 sky130_fd_sc_hd__buf_1
Xinput103 io_i_2_in1[0] vssd1 vssd1 vccd1 vccd1 _2878_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput136 io_i_5_in1[6] vssd1 vssd1 vccd1 vccd1 _2339_/A sky130_fd_sc_hd__clkbuf_1
Xinput125 io_i_4_in1[4] vssd1 vssd1 vccd1 vccd1 _3007_/A3 sky130_fd_sc_hd__buf_1
Xinput158 io_we_i vssd1 vssd1 vccd1 vccd1 _1432_/A sky130_fd_sc_hd__buf_1
Xinput147 io_i_7_ci vssd1 vssd1 vccd1 vccd1 _2515_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3080_ _3138_/CLK _3080_/D vssd1 vssd1 vccd1 vccd1 _3080_/Q sky130_fd_sc_hd__dfxtp_1
X_2100_ _3053_/Q _3002_/X _2102_/S vssd1 vssd1 vccd1 vccd1 _3053_/D sky130_fd_sc_hd__mux2_1
X_2031_ _3063_/Q _2733_/X _2031_/S vssd1 vssd1 vccd1 vccd1 _3063_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2933_ _2394_/Y _2311_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2933_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2864_ _2482_/Y _2354_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1815_ _2757_/X vssd1 vssd1 vccd1 vccd1 _2427_/B sky130_fd_sc_hd__buf_1
X_2795_ _2480_/Y _2794_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__mux2_2
X_1746_ _2779_/X _2892_/X vssd1 vssd1 vccd1 vccd1 _1753_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1677_ _2787_/X _2853_/X vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__nand2_2
XFILLER_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2229_ _2252_/S _3022_/Q vssd1 vssd1 vccd1 vccd1 _2230_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1600_ input8/X _1606_/B _1603_/C vssd1 vssd1 vccd1 vccd1 _1600_/Y sky130_fd_sc_hd__nor3_1
X_2580_ _2468_/Y _2542_/Y _2577_/Y _2578_/Y _2579_/Y vssd1 vssd1 vccd1 vccd1 _2580_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_1531_ _3188_/Q _1522_/X _1525_/X _1530_/Y vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__o211a_1
X_1462_ _3205_/Q _1458_/X _1459_/X _1461_/Y vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__o211a_1
X_3201_ _3201_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3132_ _3205_/CLK _3132_/D vssd1 vssd1 vccd1 vccd1 _3132_/Q sky130_fd_sc_hd__dfxtp_1
X_3063_ _3123_/CLK _3063_/D vssd1 vssd1 vccd1 vccd1 _3063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2014_ _2729_/X vssd1 vssd1 vccd1 vccd1 _2106_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _2419_/Y _2915_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2916_/X sky130_fd_sc_hd__mux2_2
X_2847_ _2502_/Y _2846_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__mux2_2
X_2778_ _2236_/Y _2299_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2778_/X sky130_fd_sc_hd__mux2_1
X_1729_ _3126_/Q vssd1 vssd1 vccd1 vccd1 _1729_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2701_ _2701_/A vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2632_ _3149_/Q _2632_/B _2632_/C vssd1 vssd1 vccd1 vccd1 _2632_/Y sky130_fd_sc_hd__nand3_2
Xoutput215 _3089_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput204 _3103_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput226 _3075_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[4] sky130_fd_sc_hd__clkbuf_2
X_2563_ _3203_/Q _2627_/B _2593_/C vssd1 vssd1 vccd1 vccd1 _2564_/B sky130_fd_sc_hd__nand3_1
X_1514_ _1501_/X _1516_/B _1617_/B vssd1 vssd1 vccd1 vccd1 _1514_/Y sky130_fd_sc_hd__nand3b_1
Xoutput248 _2725_/X vssd1 vssd1 vccd1 vccd1 io_vco sky130_fd_sc_hd__clkbuf_2
Xoutput237 _3061_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput259 _2679_/X vssd1 vssd1 vccd1 vccd1 io_wo[19] sky130_fd_sc_hd__clkbuf_2
X_2494_ _3111_/Q vssd1 vssd1 vccd1 vccd1 _2494_/Y sky130_fd_sc_hd__inv_2
X_1445_ _3209_/Q _1435_/X _1438_/X _1444_/Y vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__o211a_1
X_3115_ _3139_/CLK _3115_/D vssd1 vssd1 vccd1 vccd1 _3115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3166_/CLK _3046_/D vssd1 vssd1 vccd1 vccd1 _3046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _1995_/A _1995_/B _1995_/C vssd1 vssd1 vccd1 vccd1 _1994_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2615_ _2596_/X _3197_/Q _2627_/C vssd1 vssd1 vccd1 vccd1 _2615_/Y sky130_fd_sc_hd__nand3b_2
X_2546_ _2593_/B _3186_/Q _2632_/C vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__nand3b_4
X_2477_ _2869_/X vssd1 vssd1 vccd1 vccd1 _2477_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _3166_/CLK _3029_/D vssd1 vssd1 vccd1 vccd1 _3029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2400_ _3016_/Q vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2331_ _2331_/A vssd1 vssd1 vccd1 vccd1 _2331_/Y sky130_fd_sc_hd__inv_2
X_2262_ _2259_/X _2260_/Y _1666_/X _2261_/Y vssd1 vssd1 vccd1 vccd1 _3015_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2193_ _3009_/X _2841_/X vssd1 vssd1 vccd1 vccd1 _2194_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1977_ _3002_/X _2961_/X vssd1 vssd1 vccd1 vccd1 _1993_/A sky130_fd_sc_hd__nor2_1
X_2529_ _1906_/Y _2528_/Y _1908_/Y _1911_/A vssd1 vssd1 vccd1 vccd1 _2536_/A sky130_fd_sc_hd__a31oi_4
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2880_ _2463_/Y _2879_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ _1905_/A _1900_/B vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__nor2_4
X_1831_ _1845_/A _1831_/B _1845_/B vssd1 vssd1 vccd1 vccd1 _1831_/Y sky130_fd_sc_hd__nand3_4
X_1762_ _2767_/X vssd1 vssd1 vccd1 vccd1 _1763_/A sky130_fd_sc_hd__inv_2
X_1693_ _1693_/A vssd1 vssd1 vccd1 vccd1 _2290_/S sky130_fd_sc_hd__buf_2
X_2314_ _3058_/Q vssd1 vssd1 vccd1 vccd1 _2314_/Y sky130_fd_sc_hd__inv_2
X_2245_ _1666_/X _2242_/Y _2244_/Y vssd1 vssd1 vccd1 vccd1 _3019_/D sky130_fd_sc_hd__o21ai_1
X_2176_ _3037_/Q _2994_/X _2177_/S vssd1 vssd1 vccd1 vccd1 _3037_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput104 io_i_2_in1[1] vssd1 vssd1 vccd1 vccd1 _2881_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput115 io_i_3_in1[3] vssd1 vssd1 vccd1 vccd1 _2911_/A0 sky130_fd_sc_hd__buf_1
Xinput126 io_i_4_in1[5] vssd1 vssd1 vccd1 vccd1 _3006_/A3 sky130_fd_sc_hd__buf_1
Xinput159 wb_rst_i vssd1 vssd1 vccd1 vccd1 _1599_/A sky130_fd_sc_hd__clkbuf_2
Xinput148 io_i_7_in1[0] vssd1 vssd1 vccd1 vccd1 _2438_/A sky130_fd_sc_hd__buf_1
Xinput137 io_i_5_in1[7] vssd1 vssd1 vccd1 vccd1 _2331_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2030_ _3064_/Q _2735_/X _2031_/S vssd1 vssd1 vccd1 vccd1 _3064_/D sky130_fd_sc_hd__mux2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2932_ _3009_/A3 _3105_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2932_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ input97/X _3018_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1814_ _2755_/X _2907_/X vssd1 vssd1 vccd1 vccd1 _1861_/A sky130_fd_sc_hd__xor2_4
X_2794_ _2422_/Y _2352_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2794_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1745_ _2777_/X _2889_/X vssd1 vssd1 vccd1 vccd1 _1779_/A sky130_fd_sc_hd__xor2_4
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1676_ _2789_/X _2856_/X vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__and2_1
X_2228_ _2803_/X vssd1 vssd1 vccd1 vccd1 _2252_/S sky130_fd_sc_hd__inv_2
X_2159_ _2158_/X _3043_/Q _2164_/S vssd1 vssd1 vccd1 vccd1 _3043_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1530_ _1518_/X _1530_/B _1631_/B vssd1 vssd1 vccd1 vccd1 _1530_/Y sky130_fd_sc_hd__nand3b_1
X_1461_ _1472_/A _1629_/B vssd1 vssd1 vccd1 vccd1 _1461_/Y sky130_fd_sc_hd__nand2_1
X_3200_ _3201_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_2
X_3131_ _3205_/CLK _3131_/D vssd1 vssd1 vccd1 vccd1 _3131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3062_ _3166_/CLK _3062_/D vssd1 vssd1 vccd1 vccd1 _3062_/Q sky130_fd_sc_hd__dfxtp_1
X_2013_ _1962_/Y _1957_/X _1961_/Y vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2915_ _2420_/Y _2346_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2846_ _2503_/Y _2236_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2777_ _2453_/Y _2776_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2777_/X sky130_fd_sc_hd__mux2_4
X_1728_ _3127_/Q _2512_/A _1728_/S vssd1 vssd1 vccd1 vccd1 _3127_/D sky130_fd_sc_hd__mux2_1
X_1659_ _2749_/X vssd1 vssd1 vccd1 vccd1 _1659_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3205_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__clkbuf_1
X_2631_ _2603_/B _3201_/Q _2631_/C vssd1 vssd1 vccd1 vccd1 _2631_/Y sky130_fd_sc_hd__nand3b_2
Xoutput205 _3104_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput216 _3090_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[3] sky130_fd_sc_hd__clkbuf_2
X_2562_ _2598_/A vssd1 vssd1 vccd1 vccd1 _2593_/C sky130_fd_sc_hd__clkbuf_2
X_1513_ _3195_/Q _1506_/X _1510_/X _1512_/Y vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__o211a_1
Xoutput227 _3076_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput238 _3062_/Q vssd1 vssd1 vccd1 vccd1 io_o_6_out[7] sky130_fd_sc_hd__clkbuf_2
Xoutput249 _2660_/X vssd1 vssd1 vccd1 vccd1 io_wo[0] sky130_fd_sc_hd__clkbuf_2
X_2493_ _2493_/A _2787_/X vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1444_ _1451_/A _1619_/B vssd1 vssd1 vccd1 vccd1 _1444_/Y sky130_fd_sc_hd__nand2_1
X_3114_ _3139_/CLK _3114_/D vssd1 vssd1 vccd1 vccd1 _3114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3045_ _3166_/CLK _3045_/D vssd1 vssd1 vccd1 vccd1 _3045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2829_ _2441_/Y _2828_/X _3177_/Q vssd1 vssd1 vccd1 vccd1 _2829_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _1993_/A _1993_/B vssd1 vssd1 vccd1 vccd1 _1995_/C sky130_fd_sc_hd__nor2_1
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2614_ _2611_/X _3181_/Q _2630_/C vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__nand3b_2
X_2545_ _2603_/C vssd1 vssd1 vccd1 vccd1 _2632_/C sky130_fd_sc_hd__clkbuf_4
X_2476_ _3117_/Q vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _3075_/CLK _3028_/D vssd1 vssd1 vccd1 vccd1 _3028_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2330_ _2330_/A vssd1 vssd1 vccd1 vccd1 _2330_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2261_ _3015_/Q vssd1 vssd1 vccd1 vccd1 _2261_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2192_ _3023_/Q _2980_/X _2192_/S vssd1 vssd1 vccd1 vccd1 _3023_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1976_ _1998_/A _1998_/B _2000_/A vssd1 vssd1 vccd1 vccd1 _1995_/A sky130_fd_sc_hd__nand3_4
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2528_ _2528_/A vssd1 vssd1 vccd1 vccd1 _2528_/Y sky130_fd_sc_hd__inv_2
X_2459_ _2884_/X vssd1 vssd1 vccd1 vccd1 _2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1830_ _1830_/A _1830_/B vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__nor2_4
X_1761_ _2524_/A _1759_/A _1756_/Y _1754_/Y vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__o211a_1
X_1692_ _2785_/X vssd1 vssd1 vccd1 vccd1 _1693_/A sky130_fd_sc_hd__inv_2
X_2313_ _2313_/A _2313_/B vssd1 vssd1 vccd1 vccd1 _2313_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3189_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2244_ _2244_/A _2244_/B _2244_/C vssd1 vssd1 vccd1 vccd1 _2244_/Y sky130_fd_sc_hd__nand3_1
X_2175_ _3038_/Q _2995_/X _2177_/S vssd1 vssd1 vccd1 vccd1 _3038_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1959_ _2825_/X vssd1 vssd1 vccd1 vccd1 _1959_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput105 io_i_2_in1[2] vssd1 vssd1 vccd1 vccd1 _2884_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput116 io_i_3_in1[4] vssd1 vssd1 vccd1 vccd1 _2914_/A0 sky130_fd_sc_hd__buf_1
Xinput127 io_i_4_in1[6] vssd1 vssd1 vccd1 vccd1 _3005_/A3 sky130_fd_sc_hd__buf_1
XFILLER_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput149 io_i_7_in1[1] vssd1 vssd1 vccd1 vccd1 _2434_/A sky130_fd_sc_hd__buf_1
Xinput138 io_i_6_ci vssd1 vssd1 vccd1 vccd1 _2330_/A sky130_fd_sc_hd__buf_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2931_ _2397_/Y _2930_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__mux2_2
X_2862_ _2484_/Y _2861_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2793_ _2483_/Y _2792_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__mux2_1
X_1813_ _1807_/X _1811_/Y _1812_/Y vssd1 vssd1 vccd1 vccd1 _1861_/B sky130_fd_sc_hd__o21bai_2
X_1744_ _1785_/B _1785_/A _1783_/A _1743_/Y vssd1 vssd1 vccd1 vccd1 _1779_/B sky130_fd_sc_hd__a31o_2
XFILLER_7_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1675_ _2267_/A vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__inv_2
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2227_ _2227_/A _2244_/B vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2158_ _2158_/A _2158_/B vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__xor2_1
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2089_ _2088_/X _3057_/Q _2089_/S vssd1 vssd1 vccd1 vccd1 _3057_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1460_ _1460_/A vssd1 vssd1 vccd1 vccd1 _1629_/B sky130_fd_sc_hd__clkinv_4
X_3130_ _3139_/CLK _3130_/D vssd1 vssd1 vccd1 vccd1 _3130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3061_ _3075_/CLK _3061_/D vssd1 vssd1 vccd1 vccd1 _3061_/Q sky130_fd_sc_hd__dfxtp_1
X_2012_ _3072_/Q vssd1 vssd1 vccd1 vccd1 _2012_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2914_ _2914_/A0 _3123_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_2845_ _2504_/Y _2844_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__mux2_2
X_2776_ _2242_/Y _2303_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2776_/X sky130_fd_sc_hd__mux2_1
X_1727_ _3011_/X vssd1 vssd1 vccd1 vccd1 _2512_/A sky130_fd_sc_hd__inv_2
X_1658_ _1667_/A _1657_/X vssd1 vssd1 vccd1 vccd1 _3147_/D sky130_fd_sc_hd__nor2b_1
X_1589_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1673_/A sky130_fd_sc_hd__buf_2
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _2603_/C _3185_/Q _2630_/C vssd1 vssd1 vccd1 vccd1 _2630_/Y sky130_fd_sc_hd__nand3b_2
Xoutput206 _3105_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput217 _3091_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[4] sky130_fd_sc_hd__clkbuf_2
X_2561_ _2605_/C vssd1 vssd1 vccd1 vccd1 _2627_/B sky130_fd_sc_hd__buf_2
X_2492_ _2854_/X vssd1 vssd1 vccd1 vccd1 _2492_/Y sky130_fd_sc_hd__inv_2
Xoutput239 _2657_/Y vssd1 vssd1 vccd1 vccd1 io_o_7_co sky130_fd_sc_hd__clkbuf_2
Xoutput228 _3077_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[6] sky130_fd_sc_hd__clkbuf_2
X_1512_ _1501_/X _1516_/B _2658_/B vssd1 vssd1 vccd1 vccd1 _1512_/Y sky130_fd_sc_hd__nand3b_1
X_1443_ _1443_/A vssd1 vssd1 vccd1 vccd1 _1619_/B sky130_fd_sc_hd__inv_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3113_ _3138_/CLK _3113_/D vssd1 vssd1 vccd1 vccd1 _3113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _3075_/CLK _3044_/D vssd1 vssd1 vccd1 vccd1 _3044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2828_ _2442_/Y _2538_/A _3176_/Q vssd1 vssd1 vccd1 vccd1 _2828_/X sky130_fd_sc_hd__mux2_1
X_2759_ _2421_/Y _2758_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__mux2_8
XFILLER_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ _3077_/Q vssd1 vssd1 vccd1 vccd1 _1992_/Y sky130_fd_sc_hd__inv_2
X_2613_ _1608_/Y _2608_/X _2609_/Y _2610_/Y _2612_/Y vssd1 vssd1 vccd1 vccd1 _2613_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_2544_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2603_/C sky130_fd_sc_hd__buf_1
X_2475_ _2484_/A _2799_/X vssd1 vssd1 vccd1 vccd1 _2475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3027_ _3075_/CLK _3027_/D vssd1 vssd1 vccd1 vccd1 _3027_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2260_ _2257_/Y _2258_/Y _2196_/Y _2252_/S vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__a31oi_1
X_2191_ _3024_/Q _2981_/X _2192_/S vssd1 vssd1 vccd1 vccd1 _3024_/D sky130_fd_sc_hd__mux2_1
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1980_/A _1975_/B vssd1 vssd1 vccd1 vccd1 _2000_/A sky130_fd_sc_hd__nor2_4
X_2527_ _1831_/Y _2526_/Y _1833_/Y _1836_/A vssd1 vssd1 vccd1 vccd1 _2537_/A sky130_fd_sc_hd__a31oi_4
X_2458_ _3098_/Q vssd1 vssd1 vccd1 vccd1 _2458_/Y sky130_fd_sc_hd__inv_2
X_2389_ _2393_/A _2741_/X vssd1 vssd1 vccd1 vccd1 _2389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1760_ _1754_/Y _1756_/Y _1759_/Y vssd1 vssd1 vccd1 vccd1 _1760_/Y sky130_fd_sc_hd__a21boi_1
X_1691_ _1691_/A _1691_/B vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__xor2_1
X_2312_ _3122_/Q vssd1 vssd1 vccd1 vccd1 _2312_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2243_ _2208_/A _2208_/C _2208_/B vssd1 vssd1 vccd1 vccd1 _2244_/A sky130_fd_sc_hd__a21o_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2174_ _2184_/S _2170_/Y _2172_/X _2173_/Y vssd1 vssd1 vccd1 vccd1 _3039_/D sky130_fd_sc_hd__o22ai_1
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1958_ _2996_/X _2949_/X vssd1 vssd1 vccd1 vccd1 _2019_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1889_ _2737_/X _2931_/X vssd1 vssd1 vccd1 vccd1 _1936_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 io_i_2_in1[3] vssd1 vssd1 vccd1 vccd1 _2887_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput117 io_i_3_in1[5] vssd1 vssd1 vccd1 vccd1 _2917_/A0 sky130_fd_sc_hd__buf_1
Xinput139 io_i_6_in1[0] vssd1 vssd1 vccd1 vccd1 _2326_/A sky130_fd_sc_hd__buf_1
Xinput128 io_i_4_in1[7] vssd1 vssd1 vccd1 vccd1 _3004_/A3 sky130_fd_sc_hd__buf_1
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2930_ _2398_/Y _2318_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__mux2_1
X_2861_ _2485_/Y _2360_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2861_/X sky130_fd_sc_hd__mux2_1
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1812_ _2753_/X _2904_/X vssd1 vssd1 vccd1 vccd1 _1812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2792_ _2426_/Y _2358_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2792_/X sky130_fd_sc_hd__mux2_1
X_1743_ _2457_/B _2886_/X _1742_/X vssd1 vssd1 vccd1 vccd1 _1743_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1674_ _2795_/X _2865_/X vssd1 vssd1 vccd1 vccd1 _2267_/A sky130_fd_sc_hd__xor2_2
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2226_ _2226_/A _2226_/B vssd1 vssd1 vccd1 vccd1 _2227_/A sky130_fd_sc_hd__nand2_1
X_2157_ _2156_/X _3044_/Q _2164_/S vssd1 vssd1 vccd1 vccd1 _3044_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2088_ _2088_/A _2088_/B vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__xor2_2
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3075_/CLK _3060_/D vssd1 vssd1 vccd1 vccd1 _3060_/Q sky130_fd_sc_hd__dfxtp_1
X_2011_ _2010_/X _3073_/Q _2011_/S vssd1 vssd1 vccd1 vccd1 _3073_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2913_ _2423_/Y _2912_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__mux2_4
X_2844_ _2505_/Y _2242_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2844_/X sky130_fd_sc_hd__mux2_1
X_2775_ _2456_/Y _2774_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__mux2_1
X_1726_ _3128_/Q _2510_/A _1728_/S vssd1 vssd1 vccd1 vccd1 _3128_/D sky130_fd_sc_hd__mux2_1
X_1657_ _2017_/A vssd1 vssd1 vccd1 vccd1 _1657_/X sky130_fd_sc_hd__buf_2
X_1588_ _3169_/Q vssd1 vssd1 vccd1 vccd1 _1588_/Y sky130_fd_sc_hd__inv_2
X_3189_ _3189_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2209_ _2845_/X _3007_/X vssd1 vssd1 vccd1 vccd1 _2237_/A sky130_fd_sc_hd__and2b_2
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput207 _3106_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[3] sky130_fd_sc_hd__clkbuf_2
X_2560_ _2548_/A _3187_/Q _2631_/C vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__nand3b_1
X_2491_ _3112_/Q vssd1 vssd1 vccd1 vccd1 _2491_/Y sky130_fd_sc_hd__inv_2
X_1511_ _1511_/A vssd1 vssd1 vccd1 vccd1 _2658_/B sky130_fd_sc_hd__inv_2
Xoutput218 _3092_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput229 _3078_/Q vssd1 vssd1 vccd1 vccd1 io_o_5_out[7] sky130_fd_sc_hd__clkbuf_2
X_1442_ _2404_/A _1435_/X _1438_/X _1441_/Y vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _3138_/CLK _3112_/D vssd1 vssd1 vccd1 vccd1 _3112_/Q sky130_fd_sc_hd__dfxtp_1
X_3043_ _3075_/CLK _3043_/D vssd1 vssd1 vccd1 vccd1 _3043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2827_ _2406_/Y _2826_/X _3179_/Q vssd1 vssd1 vccd1 vccd1 _2827_/X sky130_fd_sc_hd__mux2_2
X_2758_ _2354_/Y _2422_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1709_ _2833_/X _1679_/Y _1707_/Y _1805_/S vssd1 vssd1 vccd1 vccd1 _1709_/Y sky130_fd_sc_hd__o31ai_1
X_2689_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1991_ _1657_/X _1956_/Y _1990_/Y vssd1 vssd1 vccd1 vccd1 _3078_/D sky130_fd_sc_hd__o21ai_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2612_ _2611_/X _3180_/Q _2620_/C vssd1 vssd1 vccd1 vccd1 _2612_/Y sky130_fd_sc_hd__nand3b_2
X_2543_ _2605_/C vssd1 vssd1 vccd1 vccd1 _2593_/B sky130_fd_sc_hd__clkbuf_2
X_2474_ _2872_/X vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3026_ _3074_/CLK _3026_/D vssd1 vssd1 vccd1 vccd1 _3026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _3025_/Q _2982_/X _2190_/S vssd1 vssd1 vccd1 vccd1 _3025_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1974_ _3001_/X _2959_/X vssd1 vssd1 vccd1 vccd1 _1975_/B sky130_fd_sc_hd__and2_1
X_2526_ _2526_/A vssd1 vssd1 vccd1 vccd1 _2526_/Y sky130_fd_sc_hd__inv_2
X_2457_ _2457_/A _2457_/B vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__nand2_1
X_2388_ _2938_/X vssd1 vssd1 vccd1 vccd1 _2388_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3009_ input87/X _2430_/A _2317_/A _3009_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3009_/X sky130_fd_sc_hd__mux4_2
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _1699_/B _1699_/A _1697_/A _1689_/Y vssd1 vssd1 vccd1 vccd1 _1691_/B sky130_fd_sc_hd__a31oi_4
X_2311_ _3090_/Q vssd1 vssd1 vccd1 vccd1 _2311_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2242_ _3019_/Q vssd1 vssd1 vccd1 vccd1 _2242_/Y sky130_fd_sc_hd__inv_2
X_2173_ _2819_/X _2117_/Y _2171_/Y _2192_/S vssd1 vssd1 vccd1 vccd1 _2173_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _2997_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__and2_1
X_1888_ _1882_/X _1886_/Y _1887_/Y vssd1 vssd1 vccd1 vccd1 _1936_/B sky130_fd_sc_hd__o21bai_2
X_2509_ _3129_/Q vssd1 vssd1 vccd1 vccd1 _2509_/Y sky130_fd_sc_hd__inv_2
Xinput107 io_i_2_in1[4] vssd1 vssd1 vccd1 vccd1 _2890_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput118 io_i_3_in1[6] vssd1 vssd1 vccd1 vccd1 _2920_/A0 sky130_fd_sc_hd__buf_1
Xinput129 io_i_5_ci vssd1 vssd1 vccd1 vccd1 _2375_/A sky130_fd_sc_hd__buf_1
XFILLER_71_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2860_ input96/X _3017_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__mux2_1
X_1811_ _1808_/Y _1809_/Y _1867_/A vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__a21oi_4
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ _2486_/Y _2790_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__mux2_4
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1742_ _2457_/B _2886_/X _2773_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__a211o_1
X_1673_ _1673_/A _1672_/X vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__nor2b_1
X_2225_ _2220_/B _2225_/B _2225_/C vssd1 vssd1 vccd1 vccd1 _2226_/B sky130_fd_sc_hd__nand3b_1
XFILLER_85_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2156_ _2156_/A _2156_/B vssd1 vssd1 vccd1 vccd1 _2156_/X sky130_fd_sc_hd__xor2_1
X_2087_ _2086_/Y _3058_/Q _2089_/S vssd1 vssd1 vccd1 vccd1 _3058_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ _2323_/Y _2012_/Y _1938_/Y _1787_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2989_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _2010_/A _2010_/B vssd1 vssd1 vccd1 vccd1 _2010_/X sky130_fd_sc_hd__xor2_1
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2912_ _2424_/Y _2353_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2843_ _2506_/Y _2842_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__mux2_2
X_2774_ _2392_/Y _2310_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__mux2_1
X_1725_ _3010_/X vssd1 vssd1 vccd1 vccd1 _2510_/A sky130_fd_sc_hd__inv_2
X_1656_ _2729_/X vssd1 vssd1 vccd1 vccd1 _2017_/A sky130_fd_sc_hd__buf_1
X_1587_ _1614_/A vssd1 vssd1 vccd1 vccd1 _1587_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _3189_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_2
X_2208_ _2208_/A _2208_/B _2208_/C vssd1 vssd1 vccd1 vccd1 _2244_/C sky130_fd_sc_hd__nand3_4
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2139_ _2987_/X _2805_/X vssd1 vssd1 vccd1 vccd1 _2141_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput208 _3107_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[4] sky130_fd_sc_hd__clkbuf_2
X_2490_ _2493_/A _2789_/X vssd1 vssd1 vccd1 vccd1 _2490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput219 _3093_/Q vssd1 vssd1 vccd1 vccd1 io_o_4_out[6] sky130_fd_sc_hd__clkbuf_2
X_1510_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1510_/X sky130_fd_sc_hd__buf_1
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1441_ _1451_/A _1617_/B vssd1 vssd1 vccd1 vccd1 _1441_/Y sky130_fd_sc_hd__nand2_1
X_3111_ _3138_/CLK _3111_/D vssd1 vssd1 vccd1 vccd1 _3111_/Q sky130_fd_sc_hd__dfxtp_1
X_3042_ _3074_/CLK _3042_/D vssd1 vssd1 vccd1 vccd1 _3042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2826_ _2407_/Y _2537_/A _3178_/Q vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__mux2_1
X_2757_ _2425_/Y _2756_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__mux2_1
X_1708_ _1679_/Y _1707_/Y _2833_/X vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__o21a_1
X_2688_ _2688_/A vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__clkbuf_1
X_1639_ _1650_/A _1639_/B vssd1 vssd1 vccd1 vccd1 _1639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _1987_/Y _1988_/X _2011_/S vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2611_ _2611_/A vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__buf_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2542_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__inv_4
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3075_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2473_ _3118_/Q vssd1 vssd1 vccd1 vccd1 _2473_/Y sky130_fd_sc_hd__inv_2
X_3025_ _3074_/CLK _3025_/D vssd1 vssd1 vccd1 vccd1 _3025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2809_ _2649_/Y _2808_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2809_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1973_ _3001_/X _2959_/X vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__nor2_4
X_2525_ _1754_/Y _2524_/Y _1756_/Y _1759_/A vssd1 vssd1 vccd1 vccd1 _2538_/A sky130_fd_sc_hd__a31oi_4
X_2456_ _2887_/X vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2387_ _3068_/Q vssd1 vssd1 vccd1 vccd1 _2387_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3008_ input88/X _2426_/A _2310_/A _3008_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3008_/X sky130_fd_sc_hd__mux4_2
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2310_ _2310_/A vssd1 vssd1 vccd1 vccd1 _2310_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2241_ _1666_/X _2236_/Y _2240_/Y vssd1 vssd1 vccd1 vccd1 _3020_/D sky130_fd_sc_hd__o21ai_1
X_2172_ _2117_/Y _2171_/Y _2819_/X vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _3078_/Q vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__inv_2
X_1887_ _2735_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _1887_/Y sky130_fd_sc_hd__nor2_2
X_2508_ _2508_/A _2550_/A vssd1 vssd1 vccd1 vccd1 _2508_/Y sky130_fd_sc_hd__nand2_1
Xinput108 io_i_2_in1[5] vssd1 vssd1 vccd1 vccd1 _2893_/A0 sky130_fd_sc_hd__clkbuf_1
X_2439_ _2439_/A _2751_/X vssd1 vssd1 vccd1 vccd1 _2439_/Y sky130_fd_sc_hd__nand2_1
Xinput119 io_i_3_in1[7] vssd1 vssd1 vccd1 vccd1 _2923_/A0 sky130_fd_sc_hd__buf_1
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1810_ _2751_/X _2901_/X vssd1 vssd1 vccd1 vccd1 _1867_/A sky130_fd_sc_hd__nor2_4
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _2430_/Y _2363_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2790_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1741_ _1741_/A _1741_/B vssd1 vssd1 vccd1 vccd1 _1783_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1672_ _2727_/X vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__buf_2
X_2224_ _2232_/A _2224_/B _2232_/B vssd1 vssd1 vccd1 vccd1 _2225_/B sky130_fd_sc_hd__nand3_4
X_2155_ _2158_/A _2158_/B _2111_/A vssd1 vssd1 vccd1 vccd1 _2156_/B sky130_fd_sc_hd__o21bai_1
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ _2086_/A _2086_/B vssd1 vssd1 vccd1 vccd1 _2086_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _2326_/Y _2018_/Y _1942_/Y _1794_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2988_/X sky130_fd_sc_hd__mux4_2
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _1887_/Y _1882_/X _1886_/Y vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__o21a_1
Xinput90 io_i_0_in1[5] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _2911_/A0 _3122_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2911_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2842_ _2507_/Y _2392_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2773_ _2459_/Y _2772_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__mux2_2
X_1724_ _3129_/Q _2508_/A _1724_/S vssd1 vssd1 vccd1 vccd1 _3129_/D sky130_fd_sc_hd__mux2_1
X_1655_ _1655_/A vssd1 vssd1 vccd1 vccd1 _1667_/A sky130_fd_sc_hd__clkbuf_2
X_1586_ _1611_/C _2551_/A _2552_/A vssd1 vssd1 vccd1 vccd1 _1614_/A sky130_fd_sc_hd__nand3b_2
X_2207_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2208_/C sky130_fd_sc_hd__inv_2
X_3187_ _3189_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2138_ _2147_/B vssd1 vssd1 vccd1 vccd1 _2141_/C sky130_fd_sc_hd__inv_2
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2069_ _3061_/Q vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput209 _3108_/Q vssd1 vssd1 vccd1 vccd1 io_o_3_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_57_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1440_ _1440_/A vssd1 vssd1 vccd1 vccd1 _1617_/B sky130_fd_sc_hd__inv_2
X_3110_ _3110_/CLK _3110_/D vssd1 vssd1 vccd1 vccd1 _3110_/Q sky130_fd_sc_hd__dfxtp_2
X_3041_ _3074_/CLK _3041_/D vssd1 vssd1 vccd1 vccd1 _3041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ _2374_/Y _2824_/X _3181_/Q vssd1 vssd1 vccd1 vccd1 _2825_/X sky130_fd_sc_hd__mux2_2
X_2756_ _2360_/Y _2426_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__mux2_1
X_1707_ _1707_/A vssd1 vssd1 vccd1 vccd1 _1707_/Y sky130_fd_sc_hd__inv_2
X_2687_ _2687_/A vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__clkbuf_1
X_1638_ _1638_/A vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__buf_1
XFILLER_48_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1569_ _3176_/Q _1556_/X _1557_/X _1568_/Y vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2610_ _3152_/Q _2610_/B _2627_/C vssd1 vssd1 vccd1 vccd1 _2610_/Y sky130_fd_sc_hd__nand3_2
X_2541_ _2541_/A _3200_/Q vssd1 vssd1 vccd1 vccd1 _2541_/Y sky130_fd_sc_hd__nand2_1
X_2472_ _2484_/A _2801_/X vssd1 vssd1 vccd1 vccd1 _2472_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3024_ _3201_/CLK _3024_/D vssd1 vssd1 vccd1 vccd1 _3024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2808_ _2650_/Y _2651_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__mux2_1
X_2739_ _2391_/Y _2738_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1972_ _3000_/X _2957_/X vssd1 vssd1 vccd1 vccd1 _1998_/B sky130_fd_sc_hd__xor2_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2524_ _2524_/A vssd1 vssd1 vccd1 vccd1 _2524_/Y sky130_fd_sc_hd__inv_2
X_2455_ _3099_/Q vssd1 vssd1 vccd1 vccd1 _2455_/Y sky130_fd_sc_hd__inv_2
X_2386_ _2393_/A _2743_/X vssd1 vssd1 vccd1 vccd1 _2386_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007_ input89/X _2422_/A _2303_/A _3007_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3007_/X sky130_fd_sc_hd__mux4_2
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2240_ _2238_/Y _2239_/X _2252_/S vssd1 vssd1 vccd1 vccd1 _2240_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _2171_/A vssd1 vssd1 vccd1 vccd1 _2171_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ _3079_/Q _2751_/X _1955_/S vssd1 vssd1 vccd1 vccd1 _3079_/D sky130_fd_sc_hd__mux2_1
X_1886_ _1943_/A _1884_/Y _1885_/Y vssd1 vssd1 vccd1 vccd1 _1886_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2507_ _3130_/Q vssd1 vssd1 vccd1 vccd1 _2507_/Y sky130_fd_sc_hd__inv_2
Xinput109 io_i_2_in1[6] vssd1 vssd1 vccd1 vccd1 _2896_/A0 sky130_fd_sc_hd__clkbuf_1
X_2438_ _2438_/A vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__inv_2
X_2369_ _2372_/A _2997_/X vssd1 vssd1 vccd1 vccd1 _2369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _2775_/X _2886_/X vssd1 vssd1 vccd1 vccd1 _1741_/B sky130_fd_sc_hd__and2_1
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1671_ _1673_/A _1670_/X vssd1 vssd1 vccd1 vccd1 _3141_/D sky130_fd_sc_hd__nor2b_1
XFILLER_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2223_ _2217_/C _2237_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2232_/B sky130_fd_sc_hd__a21oi_4
X_2154_ _2163_/B _2127_/Y _2129_/Y vssd1 vssd1 vccd1 vccd1 _2158_/B sky130_fd_sc_hd__a21boi_2
X_2085_ _2088_/B _2088_/A _2084_/Y vssd1 vssd1 vccd1 vccd1 _2086_/B sky130_fd_sc_hd__a21oi_2
X_2987_ _2409_/Y _2032_/Y _1956_/Y _1806_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2987_/X sky130_fd_sc_hd__mux4_2
X_1938_ _3088_/Q vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__inv_2
X_1869_ _1867_/Y _1809_/Y _1808_/Y _1862_/S vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__a31oi_1
Xinput91 io_i_0_in1[6] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
Xinput80 io_eo[6] vssd1 vssd1 vccd1 vccd1 _2666_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2910_ _2427_/Y _2909_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2841_ _2508_/Y _2840_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__mux2_2
X_2772_ _2396_/Y _2317_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__mux2_1
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1723_ _3009_/X vssd1 vssd1 vccd1 vccd1 _2508_/A sky130_fd_sc_hd__inv_2
X_1654_ _2654_/A _1642_/X _1459_/A _1653_/Y vssd1 vssd1 vccd1 vccd1 _3148_/D sky130_fd_sc_hd__o211a_1
X_1585_ _3170_/Q _1570_/A _1583_/X _1584_/Y vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__o211a_1
X_2206_ _3008_/X _2843_/X vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__and2b_1
X_3186_ _3193_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_2
X_2137_ _2986_/X _2807_/X vssd1 vssd1 vccd1 vccd1 _2147_/B sky130_fd_sc_hd__and2_1
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _1672_/X _2032_/Y _2067_/Y vssd1 vssd1 vccd1 vccd1 _3062_/D sky130_fd_sc_hd__o21ai_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3040_ _3201_/CLK _3040_/D vssd1 vssd1 vccd1 vccd1 _3040_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2824_ _2375_/Y _2536_/A _3180_/Q vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__mux2_1
X_2755_ _2429_/Y _2754_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2755_/X sky130_fd_sc_hd__mux2_4
X_1706_ _3135_/Q vssd1 vssd1 vccd1 vccd1 _1706_/Y sky130_fd_sc_hd__inv_2
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__clkbuf_1
X_1637_ _3154_/Q _1626_/X _1635_/X _1636_/Y vssd1 vssd1 vccd1 vccd1 _3154_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1568_ _1565_/X _1572_/B _1621_/B vssd1 vssd1 vccd1 vccd1 _1568_/Y sky130_fd_sc_hd__nand3b_1
X_1499_ _3198_/Q _1479_/X _1490_/X _1498_/Y vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3169_ _3201_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2540_ _2540_/A vssd1 vssd1 vccd1 vccd1 _2540_/Y sky130_fd_sc_hd__inv_2
X_2471_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2484_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3023_ _3201_/CLK _3023_/D vssd1 vssd1 vccd1 vccd1 _3023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2807_ _2652_/Y _2806_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2807_/X sky130_fd_sc_hd__mux2_1
X_2738_ _2312_/Y _2392_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2738_/X sky130_fd_sc_hd__mux2_1
X_2669_ _2669_/A vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1971_ _2010_/B _2010_/A _2008_/A _1970_/Y vssd1 vssd1 vccd1 vccd1 _1998_/A sky130_fd_sc_hd__a31o_1
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2523_ _2521_/Y _2522_/Y _2279_/A vssd1 vssd1 vccd1 vccd1 _2539_/A sky130_fd_sc_hd__a21oi_4
X_2454_ _2457_/A _2777_/X vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__nand2_1
X_2385_ _2941_/X vssd1 vssd1 vccd1 vccd1 _2385_/Y sky130_fd_sc_hd__inv_2
Xinput1 io_adr_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
X_3006_ input90/X _2418_/A _2299_/A _3006_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3006_/X sky130_fd_sc_hd__mux4_2
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_0 _2688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2170_ _3039_/Q vssd1 vssd1 vccd1 vccd1 _2170_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1954_ _3080_/Q _2753_/X _1955_/S vssd1 vssd1 vccd1 vccd1 _3080_/D sky130_fd_sc_hd__mux2_1
X_1885_ _2733_/X _2925_/X vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__nor2_4
X_2506_ _2506_/A _2506_/B vssd1 vssd1 vccd1 vccd1 _2506_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2437_ _2902_/X vssd1 vssd1 vccd1 vccd1 _2437_/Y sky130_fd_sc_hd__inv_2
X_2368_ _2368_/A vssd1 vssd1 vccd1 vccd1 _2368_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2299_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2299_/Y sky130_fd_sc_hd__inv_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput190 _3139_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[4] sky130_fd_sc_hd__clkbuf_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1670_ _2026_/A vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__buf_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2222_ _3008_/X _2202_/Y _2208_/B _2221_/Y _2208_/A vssd1 vssd1 vccd1 vccd1 _2232_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2153_ _2153_/A vssd1 vssd1 vccd1 vccd1 _2158_/A sky130_fd_sc_hd__inv_2
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2084_ _2990_/X _2969_/X vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _2414_/Y _2069_/Y _1992_/Y _1842_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2986_/X sky130_fd_sc_hd__mux4_2
X_1937_ _1936_/X _3089_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _3089_/D sky130_fd_sc_hd__mux2_1
X_1868_ _1867_/Y _1808_/Y _1809_/Y vssd1 vssd1 vccd1 vccd1 _1868_/X sky130_fd_sc_hd__a21o_1
Xinput70 io_eo[55] vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__clkbuf_1
Xinput81 io_eo[7] vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__clkbuf_2
X_1799_ _2797_/X vssd1 vssd1 vccd1 vccd1 _2478_/B sky130_fd_sc_hd__buf_1
Xinput92 io_i_0_in1[7] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2509_/Y _2396_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2840_/X sky130_fd_sc_hd__mux2_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2462_/Y _2770_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2771_/X sky130_fd_sc_hd__mux2_1
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _3130_/Q _2506_/A _1724_/S vssd1 vssd1 vccd1 vccd1 _3130_/D sky130_fd_sc_hd__mux2_1
X_1653_ _2658_/A _1653_/B vssd1 vssd1 vccd1 vccd1 _1653_/Y sky130_fd_sc_hd__nand2_1
X_1584_ _1590_/A _1584_/B _1636_/B vssd1 vssd1 vccd1 vccd1 _1584_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2205_ _3007_/X _2845_/X vssd1 vssd1 vccd1 vccd1 _2208_/B sky130_fd_sc_hd__xnor2_4
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _3201_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2113_/Y _2149_/B _2136_/C vssd1 vssd1 vccd1 vccd1 _2141_/A sky130_fd_sc_hd__nand3b_2
X_2067_ _2063_/Y _2064_/X _2089_/S vssd1 vssd1 vccd1 vccd1 _2067_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ _2320_/Y _2968_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__mux2_4
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ _2329_/Y _2822_/X _3183_/Q vssd1 vssd1 vccd1 vccd1 _2823_/X sky130_fd_sc_hd__mux2_1
X_2754_ _2365_/Y _2430_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__mux2_1
X_1705_ _1796_/S _1701_/Y _1702_/X _1704_/Y vssd1 vssd1 vccd1 vccd1 _3136_/D sky130_fd_sc_hd__o22ai_1
X_2685_ _2685_/A vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__clkbuf_1
X_1636_ _1636_/A _1636_/B vssd1 vssd1 vccd1 vccd1 _1636_/Y sky130_fd_sc_hd__nand2_1
X_1567_ _3177_/Q _1556_/X _1557_/X _1566_/Y vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__o211a_1
X_1498_ _1609_/B _1498_/B _1648_/B vssd1 vssd1 vccd1 vccd1 _1498_/Y sky130_fd_sc_hd__nand3b_1
X_3168_ _3201_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_4
X_2119_ _2981_/X _2817_/X vssd1 vssd1 vccd1 vccd1 _2119_/Y sky130_fd_sc_hd__nor2_2
X_3099_ _3123_/CLK _3099_/D vssd1 vssd1 vccd1 vccd1 _3099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2470_ _2875_/X vssd1 vssd1 vccd1 vccd1 _2470_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3022_ _3205_/CLK _3022_/D vssd1 vssd1 vccd1 vccd1 _3022_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2806_ _2653_/Y _2145_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__mux2_1
X_2737_ _2395_/Y _2736_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__mux2_2
X_2668_ _2668_/A vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__clkbuf_1
X_1619_ _1627_/A _1619_/B vssd1 vssd1 vccd1 vccd1 _1619_/Y sky130_fd_sc_hd__nand2_1
X_2599_ _3210_/Q _2610_/B _2627_/C vssd1 vssd1 vccd1 vccd1 _2599_/Y sky130_fd_sc_hd__nand3_2
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _2361_/B _2955_/X _1969_/X vssd1 vssd1 vccd1 vccd1 _1970_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2522_ _2522_/A vssd1 vssd1 vccd1 vccd1 _2522_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2453_ _2890_/X vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__inv_2
X_2384_ _3069_/Q vssd1 vssd1 vccd1 vccd1 _2384_/Y sky130_fd_sc_hd__inv_2
Xinput2 io_adr_i[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
XFILLER_28_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3005_ input91/X _2414_/A _2295_/A _3005_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3005_/X sky130_fd_sc_hd__mux4_2
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_1 _2698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3092_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1953_ _3081_/Q _2755_/X _1955_/S vssd1 vssd1 vccd1 vccd1 _3081_/D sky130_fd_sc_hd__mux2_1
X_1884_ _2827_/X vssd1 vssd1 vccd1 vccd1 _1884_/Y sky130_fd_sc_hd__inv_2
X_2505_ _3131_/Q vssd1 vssd1 vccd1 vccd1 _2505_/Y sky130_fd_sc_hd__inv_2
X_2436_ _3080_/Q vssd1 vssd1 vccd1 vccd1 _2436_/Y sky130_fd_sc_hd__inv_2
X_2367_ _3049_/Q vssd1 vssd1 vccd1 vccd1 _2367_/Y sky130_fd_sc_hd__inv_2
X_2298_ _3076_/Q vssd1 vssd1 vccd1 vccd1 _2298_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput180 _3018_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput191 _3012_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2221_ _3006_/X _2847_/X vssd1 vssd1 vccd1 vccd1 _2221_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2152_ _2184_/S _2145_/Y _2151_/X vssd1 vssd1 vccd1 vccd1 _3045_/D sky130_fd_sc_hd__o21ai_1
X_2083_ _2082_/X _3059_/Q _2089_/S vssd1 vssd1 vccd1 vccd1 _3059_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2985_ _2418_/Y _2075_/Y _2298_/Y _2346_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2985_/X sky130_fd_sc_hd__mux4_2
X_1936_ _1936_/A _1936_/B vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__xor2_1
X_1867_ _1867_/A vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__inv_2
Xinput71 io_eo[56] vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__clkbuf_1
X_1798_ _3117_/Q _2799_/X _1803_/S vssd1 vssd1 vccd1 vccd1 _3117_/D sky130_fd_sc_hd__mux2_1
Xinput82 io_eo[8] vssd1 vssd1 vccd1 vccd1 _2668_/A sky130_fd_sc_hd__clkbuf_2
Xinput60 io_eo[46] vssd1 vssd1 vccd1 vccd1 _2706_/A sky130_fd_sc_hd__clkbuf_1
Xinput93 io_i_1_ci vssd1 vssd1 vccd1 vccd1 _2496_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2419_ _2427_/A _2761_/X vssd1 vssd1 vccd1 vccd1 _2419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _2400_/Y _2323_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2770_/X sky130_fd_sc_hd__mux2_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _3008_/X vssd1 vssd1 vccd1 vccd1 _2506_/A sky130_fd_sc_hd__inv_2
X_1652_ _3148_/Q vssd1 vssd1 vccd1 vccd1 _2654_/A sky130_fd_sc_hd__clkbuf_2
X_1583_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1583_/X sky130_fd_sc_hd__clkbuf_2
X_2204_ _2251_/A _2251_/B _2203_/Y vssd1 vssd1 vccd1 vccd1 _2208_/A sky130_fd_sc_hd__o21bai_4
X_3184_ _3197_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2135_ _2147_/A vssd1 vssd1 vccd1 vccd1 _2136_/C sky130_fd_sc_hd__inv_2
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2066_ _2066_/A vssd1 vssd1 vccd1 vccd1 _2089_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ _2322_/Y _2321_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__mux2_1
X_1919_ _1920_/A _1920_/B _1920_/C vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__a21oi_1
X_2899_ _2899_/A0 _3014_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _2330_/Y _2535_/A _3182_/Q vssd1 vssd1 vccd1 vccd1 _2822_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2753_ _2433_/Y _2752_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__mux2_1
X_1704_ _1681_/Y _1676_/X _1680_/Y _1805_/S vssd1 vssd1 vccd1 vccd1 _1704_/Y sky130_fd_sc_hd__o31ai_1
X_2684_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__clkbuf_1
X_1635_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__clkbuf_2
X_1566_ _1565_/X _1572_/B _1619_/B vssd1 vssd1 vccd1 vccd1 _1566_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1497_ input7/X vssd1 vssd1 vccd1 vccd1 _1648_/B sky130_fd_sc_hd__inv_2
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _3211_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_4
X_3098_ _3139_/CLK _3098_/D vssd1 vssd1 vccd1 vccd1 _3098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _2171_/A _2116_/Y _2117_/Y vssd1 vssd1 vccd1 vccd1 _2118_/Y sky130_fd_sc_hd__a21oi_4
X_2049_ _2993_/X _2975_/X vssd1 vssd1 vccd1 vccd1 _2056_/A sky130_fd_sc_hd__nor2_4
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3021_ _3189_/CLK _3021_/D vssd1 vssd1 vccd1 vccd1 _3021_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ _2654_/Y _2804_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__mux2_2
X_2736_ _2319_/Y _2396_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__mux2_1
X_2667_ _2667_/A vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1618_ _3162_/Q _1613_/X _1583_/X _1617_/Y vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__o211a_1
X_2598_ _2598_/A vssd1 vssd1 vccd1 vccd1 _2627_/C sky130_fd_sc_hd__buf_2
X_1549_ _1532_/X _1558_/B _1645_/B vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2521_ _2521_/A _2521_/B vssd1 vssd1 vccd1 vccd1 _2521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2452_ _3100_/Q vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__inv_2
X_2383_ _2393_/A _2745_/X vssd1 vssd1 vccd1 vccd1 _2383_/Y sky130_fd_sc_hd__nand2_1
Xinput3 io_cs_i vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
X_3004_ input92/X _2409_/A _2291_/A _3004_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3004_/X sky130_fd_sc_hd__mux4_2
X_2719_ _2719_/A vssd1 vssd1 vccd1 vccd1 _2719_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_2 _2667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1952_ _3082_/Q _2427_/B _1952_/S vssd1 vssd1 vccd1 vccd1 _3082_/D sky130_fd_sc_hd__mux2_1
X_1883_ _2733_/X _2925_/X vssd1 vssd1 vccd1 vccd1 _1943_/A sky130_fd_sc_hd__nand2_2
X_2504_ _2504_/A _2506_/B vssd1 vssd1 vccd1 vccd1 _2504_/Y sky130_fd_sc_hd__nand2_1
X_2435_ _2439_/A _2753_/X vssd1 vssd1 vccd1 vccd1 _2435_/Y sky130_fd_sc_hd__nand2_1
X_2366_ _2372_/A _2998_/X vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2297_ _3037_/Q vssd1 vssd1 vccd1 vccd1 _2297_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 _2580_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput181 _3019_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[4] sky130_fd_sc_hd__clkbuf_2
Xoutput192 _3013_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2220_/A _2220_/B _2224_/B vssd1 vssd1 vccd1 vccd1 _2226_/A sky130_fd_sc_hd__nand3_1
X_2151_ _2148_/Y _2149_/Y _2164_/S vssd1 vssd1 vccd1 vccd1 _2151_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2082_ _2082_/A _2082_/B vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__xor2_1
XFILLER_53_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2984_ _2422_/Y _2307_/Y _2302_/Y _2353_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2984_/X sky130_fd_sc_hd__mux4_2
X_1935_ _1934_/Y _3090_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _3090_/D sky130_fd_sc_hd__mux2_1
X_1866_ _1659_/X _1863_/Y _1864_/X _1865_/Y vssd1 vssd1 vccd1 vccd1 _3104_/D sky130_fd_sc_hd__o22ai_1
Xinput72 io_eo[57] vssd1 vssd1 vccd1 vccd1 _2717_/A sky130_fd_sc_hd__clkbuf_1
X_1797_ _1805_/S vssd1 vssd1 vccd1 vccd1 _1803_/S sky130_fd_sc_hd__buf_2
Xinput50 io_eo[37] vssd1 vssd1 vccd1 vccd1 _2697_/A sky130_fd_sc_hd__clkbuf_2
Xinput61 io_eo[47] vssd1 vssd1 vccd1 vccd1 _2707_/A sky130_fd_sc_hd__clkbuf_1
Xinput94 io_i_1_in1[0] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
Xinput83 io_eo[9] vssd1 vssd1 vccd1 vccd1 _2669_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2418_ _2418_/A vssd1 vssd1 vccd1 vccd1 _2418_/Y sky130_fd_sc_hd__inv_2
X_2349_ _2541_/A _3194_/Q vssd1 vssd1 vccd1 vccd1 _2349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _3131_/Q _2504_/A _1724_/S vssd1 vssd1 vccd1 vccd1 _3131_/D sky130_fd_sc_hd__mux2_1
X_1651_ _3149_/Q _1642_/X _1459_/A _1650_/Y vssd1 vssd1 vccd1 vccd1 _3149_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1582_ _3171_/Q _1570_/X _1571_/X _1581_/Y vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__o211a_1
X_2203_ _3008_/X _2202_/Y _2841_/X _2508_/A vssd1 vssd1 vccd1 vccd1 _2203_/Y sky130_fd_sc_hd__o2bb2ai_1
X_3183_ _3197_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2134_ _2986_/X _2807_/X vssd1 vssd1 vccd1 vccd1 _2147_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2065_ _2727_/X vssd1 vssd1 vccd1 vccd1 _2066_/A sky130_fd_sc_hd__inv_2
X_2967_ _2324_/Y _2966_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__mux2_2
X_1918_ _1918_/A _1918_/B vssd1 vssd1 vccd1 vccd1 _1920_/C sky130_fd_sc_hd__nor2_1
X_2898_ _2445_/Y _2897_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2898_/X sky130_fd_sc_hd__mux2_2
X_1849_ _2759_/X _2913_/X vssd1 vssd1 vccd1 vccd1 _1849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _2635_/Y _2820_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__mux2_2
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2752_ _1701_/Y _2434_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _2785_/X vssd1 vssd1 vccd1 vccd1 _1805_/S sky130_fd_sc_hd__clkbuf_2
X_2683_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__clkbuf_1
X_1634_ _3155_/Q _1626_/X _1623_/X _1633_/Y vssd1 vssd1 vccd1 vccd1 _3155_/D sky130_fd_sc_hd__o211a_1
X_1565_ _1611_/C vssd1 vssd1 vccd1 vccd1 _1565_/X sky130_fd_sc_hd__buf_1
X_1496_ _3199_/Q _1479_/X _1490_/X _1495_/Y vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3166_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_4
X_3097_ _3138_/CLK _3097_/D vssd1 vssd1 vccd1 vccd1 _3097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2117_ _2980_/X _2821_/X vssd1 vssd1 vccd1 vccd1 _2117_/Y sky130_fd_sc_hd__nor2_4
X_2048_ _2992_/X _2973_/X vssd1 vssd1 vccd1 vccd1 _2082_/A sky130_fd_sc_hd__xor2_4
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_3020_ _3205_/CLK _3020_/D vssd1 vssd1 vccd1 vccd1 _3020_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2804_ _2655_/Y _2107_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2804_/X sky130_fd_sc_hd__mux2_1
X_2735_ _2399_/Y _2734_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__mux2_2
X_2666_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__clkbuf_1
X_1617_ _1627_/A _1617_/B vssd1 vssd1 vccd1 vccd1 _1617_/Y sky130_fd_sc_hd__nand2_1
X_2597_ _2596_/X _3194_/Q _2618_/C vssd1 vssd1 vccd1 vccd1 _2597_/Y sky130_fd_sc_hd__nand3b_4
X_1548_ _3184_/Q _1540_/X _1541_/X _1547_/Y vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__o211a_1
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1479_ _1522_/A vssd1 vssd1 vccd1 vccd1 _1479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3211_/CLK _3149_/D vssd1 vssd1 vccd1 vccd1 _3149_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2520_ _2225_/B _2518_/Y _2225_/C _2519_/X vssd1 vssd1 vccd1 vccd1 _2540_/A sky130_fd_sc_hd__a31oi_4
X_2451_ _2457_/A _2779_/X vssd1 vssd1 vccd1 vccd1 _2451_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2382_ _3021_/Q vssd1 vssd1 vccd1 vccd1 _2382_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 io_dat_i[0] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3003_ _2331_/Y _1881_/Y _1806_/Y _2263_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _3003_/X sky130_fd_sc_hd__mux4_2
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2718_ _2718_/A vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2649_ _2654_/A _2985_/X vssd1 vssd1 vccd1 vccd1 _2649_/Y sky130_fd_sc_hd__nand2_1
XINSDIODE3_3 _3022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1951_ _3083_/Q _2759_/X _1952_/S vssd1 vssd1 vccd1 vccd1 _3083_/D sky130_fd_sc_hd__mux2_1
X_1882_ _2735_/X _2928_/X vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__and2_1
X_2503_ _3132_/Q vssd1 vssd1 vccd1 vccd1 _2503_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2434_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2434_/Y sky130_fd_sc_hd__inv_2
X_2365_ _3137_/Q vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2296_ _2313_/A _2994_/X vssd1 vssd1 vccd1 vccd1 _2296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput160 _2554_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput171 _2586_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput182 _3020_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput193 _3014_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2150_ _2150_/A vssd1 vssd1 vccd1 vccd1 _2164_/S sky130_fd_sc_hd__buf_2
X_2081_ _1672_/X _2075_/Y _2080_/Y vssd1 vssd1 vccd1 vccd1 _3060_/D sky130_fd_sc_hd__o21ai_1
X_2983_ _2426_/Y _2314_/Y _2309_/Y _2359_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2983_/X sky130_fd_sc_hd__mux4_2
X_1934_ _1934_/A _1934_/B vssd1 vssd1 vccd1 vccd1 _1934_/Y sky130_fd_sc_hd__xnor2_1
X_1865_ _1812_/Y _1807_/X _1811_/Y _1955_/S vssd1 vssd1 vccd1 vccd1 _1865_/Y sky130_fd_sc_hd__o31ai_1
Xinput40 io_eo[28] vssd1 vssd1 vccd1 vccd1 _2688_/A sky130_fd_sc_hd__clkbuf_2
Xinput73 io_eo[58] vssd1 vssd1 vccd1 vccd1 _2718_/A sky130_fd_sc_hd__clkbuf_1
X_1796_ _3118_/Q _2801_/X _1796_/S vssd1 vssd1 vccd1 vccd1 _3118_/D sky130_fd_sc_hd__mux2_1
Xinput51 io_eo[38] vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__clkbuf_2
Xinput62 io_eo[48] vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__clkbuf_1
Xinput95 io_i_1_in1[1] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
Xinput84 io_i_0_ci vssd1 vssd1 vccd1 vccd1 _2516_/A sky130_fd_sc_hd__buf_1
XFILLER_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2417_ _2917_/X vssd1 vssd1 vccd1 vccd1 _2417_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2348_ _2348_/A _3196_/Q vssd1 vssd1 vccd1 vccd1 _2348_/Y sky130_fd_sc_hd__nand2_1
X_2279_ _2279_/A _2522_/A vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1650_ _1650_/A _1650_/B vssd1 vssd1 vccd1 vccd1 _1650_/Y sky130_fd_sc_hd__nand2_1
X_1581_ _1590_/A _1584_/B _1633_/B vssd1 vssd1 vccd1 vccd1 _1581_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2202_ _2843_/X vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__inv_2
X_3182_ _3201_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_2
X_2133_ _2133_/A _2153_/A _2156_/A vssd1 vssd1 vccd1 vccd1 _2149_/B sky130_fd_sc_hd__nand3_4
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _2532_/A _2062_/A _2059_/Y _2057_/Y vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__o211a_1
X_2966_ _2325_/Y _2090_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__mux2_1
X_1917_ _3093_/Q vssd1 vssd1 vccd1 vccd1 _1917_/Y sky130_fd_sc_hd__inv_2
X_2897_ _2446_/Y _1729_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1848_ _1848_/A vssd1 vssd1 vccd1 vccd1 _1862_/S sky130_fd_sc_hd__clkbuf_2
X_1779_ _1779_/A _1779_/B vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__xor2_1
XFILLER_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2820_ _2636_/Y _2170_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__mux2_1
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ _2437_/Y _2750_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2751_/X sky130_fd_sc_hd__mux2_2
X_1702_ _1681_/Y _1676_/X _1680_/Y vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__o21a_1
X_2682_ _2682_/A vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1633_ _1636_/A _1633_/B vssd1 vssd1 vccd1 vccd1 _1633_/Y sky130_fd_sc_hd__nand2_1
X_1564_ _3178_/Q _1556_/X _1557_/X _1563_/Y vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__o211a_1
X_1495_ _1609_/B _1498_/B _1645_/B vssd1 vssd1 vccd1 vccd1 _1495_/Y sky130_fd_sc_hd__nand3b_1
X_3165_ _3211_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_4
X_3096_ _3139_/CLK _3096_/D vssd1 vssd1 vccd1 vccd1 _3096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2116_ _2819_/X vssd1 vssd1 vccd1 vccd1 _2116_/Y sky130_fd_sc_hd__inv_2
X_2047_ _2088_/B _2088_/A _2086_/A _2046_/Y vssd1 vssd1 vccd1 vccd1 _2082_/B sky130_fd_sc_hd__a31o_2
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2949_ _2372_/Y _2948_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2949_/X sky130_fd_sc_hd__mux2_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2803_ _2335_/Y _2802_/X _3187_/Q vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__mux2_2
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ _1787_/Y _2400_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__mux2_1
X_2665_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__clkbuf_1
X_1616_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1627_/A sky130_fd_sc_hd__clkbuf_2
X_2596_ _2596_/A vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__clkbuf_2
X_1547_ _1532_/X _1558_/B _1653_/B vssd1 vssd1 vccd1 vccd1 _1547_/Y sky130_fd_sc_hd__nand3b_1
X_1478_ _2605_/C _2552_/A _1590_/A vssd1 vssd1 vccd1 vccd1 _1522_/A sky130_fd_sc_hd__nor3_4
X_3148_ _3166_/CLK _3148_/D vssd1 vssd1 vccd1 vccd1 _3148_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3079_ _3138_/CLK _3079_/D vssd1 vssd1 vccd1 vccd1 _3079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2450_ _2893_/X vssd1 vssd1 vccd1 vccd1 _2450_/Y sky130_fd_sc_hd__inv_2
X_2381_ _2944_/X vssd1 vssd1 vccd1 vccd1 _2381_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 io_dat_i[10] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3002_ _2339_/Y _1917_/Y _1842_/Y _2340_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _3002_/X sky130_fd_sc_hd__mux4_2
X_2717_ _2717_/A vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__clkbuf_2
X_2648_ _3043_/Q vssd1 vssd1 vccd1 vccd1 _2648_/Y sky130_fd_sc_hd__inv_2
X_2579_ _2600_/A _2600_/B _3158_/Q vssd1 vssd1 vccd1 vccd1 _2579_/Y sky130_fd_sc_hd__nand3_2
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _3084_/Q _2761_/X _1952_/S vssd1 vssd1 vccd1 vccd1 _3084_/D sky130_fd_sc_hd__mux2_1
X_1881_ _3094_/Q vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__inv_2
X_2502_ _2502_/A _2506_/B vssd1 vssd1 vccd1 vccd1 _2502_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2433_ _2905_/X vssd1 vssd1 vccd1 vccd1 _2433_/Y sky130_fd_sc_hd__inv_2
X_2364_ _3105_/Q vssd1 vssd1 vccd1 vccd1 _2364_/Y sky130_fd_sc_hd__inv_2
X_2295_ _2295_/A vssd1 vssd1 vccd1 vccd1 _2295_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput161 _2613_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput172 _2590_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput194 _2538_/Y vssd1 vssd1 vccd1 vccd1 io_o_2_co sky130_fd_sc_hd__clkbuf_2
Xoutput183 _3021_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2080_/A _2177_/S vssd1 vssd1 vccd1 vccd1 _2080_/Y sky130_fd_sc_hd__nand2_1
X_2982_ _2430_/Y _2321_/Y _2316_/Y _2364_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2982_/X sky130_fd_sc_hd__mux4_2
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1933_ _2737_/X _2931_/X _1932_/Y vssd1 vssd1 vccd1 vccd1 _1934_/B sky130_fd_sc_hd__o21a_1
X_1864_ _1812_/Y _1807_/X _1811_/Y vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__o21a_1
Xinput30 io_eo[19] vssd1 vssd1 vccd1 vccd1 _2679_/A sky130_fd_sc_hd__clkbuf_2
Xinput63 io_eo[49] vssd1 vssd1 vccd1 vccd1 _2709_/A sky130_fd_sc_hd__clkbuf_1
X_1795_ _1792_/X _1793_/Y _1661_/X _1794_/Y vssd1 vssd1 vccd1 vccd1 _3119_/D sky130_fd_sc_hd__o2bb2ai_1
Xinput41 io_eo[29] vssd1 vssd1 vccd1 vccd1 _2689_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 io_eo[39] vssd1 vssd1 vccd1 vccd1 _2699_/A sky130_fd_sc_hd__clkbuf_2
Xinput74 io_eo[59] vssd1 vssd1 vccd1 vccd1 _2719_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3074_/CLK
+ sky130_fd_sc_hd__clkbuf_1
Xinput96 io_i_1_in1[2] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
Xinput85 io_i_0_in1[0] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
X_2416_ _3085_/Q vssd1 vssd1 vccd1 vccd1 _2416_/Y sky130_fd_sc_hd__inv_2
X_2347_ _3012_/Q vssd1 vssd1 vccd1 vccd1 _2347_/Y sky130_fd_sc_hd__inv_2
X_2278_ _2801_/X _2874_/X vssd1 vssd1 vccd1 vccd1 _2522_/A sky130_fd_sc_hd__and2_1
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _3172_/Q _1570_/X _1571_/X _1579_/Y vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__o211a_1
X_2201_ _2253_/B _2253_/C _2200_/X vssd1 vssd1 vccd1 vccd1 _2251_/B sky130_fd_sc_hd__a21oi_4
X_3181_ _3197_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2132_ _2132_/A _2132_/B vssd1 vssd1 vccd1 vccd1 _2156_/A sky130_fd_sc_hd__nor2_4
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2063_ _2057_/Y _2059_/Y _2062_/Y vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2965_ _2327_/Y _2964_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__mux2_2
X_2896_ _2896_/A0 _3013_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2896_/X sky130_fd_sc_hd__mux2_1
X_1916_ _1670_/X _1881_/Y _1915_/Y vssd1 vssd1 vccd1 vccd1 _3094_/D sky130_fd_sc_hd__o21ai_1
X_1847_ _1659_/X _1842_/Y _1846_/Y vssd1 vssd1 vccd1 vccd1 _3109_/D sky130_fd_sc_hd__o21ai_1
XFILLER_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1778_ _1661_/X _1772_/Y _1777_/Y vssd1 vssd1 vccd1 vccd1 _3124_/D sky130_fd_sc_hd__o21ai_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _1706_/Y _2438_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__mux2_1
X_1701_ _3136_/Q vssd1 vssd1 vccd1 vccd1 _1701_/Y sky130_fd_sc_hd__inv_2
X_2681_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__clkbuf_1
X_1632_ _3156_/Q _1626_/X _1623_/X _1631_/Y vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__o211a_1
X_1563_ _1551_/X _1572_/B _1617_/B vssd1 vssd1 vccd1 vccd1 _1563_/Y sky130_fd_sc_hd__nand3b_1
X_1494_ input8/X vssd1 vssd1 vccd1 vccd1 _1645_/B sky130_fd_sc_hd__inv_2
X_3164_ _3197_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_4
X_3095_ _3123_/CLK _3095_/D vssd1 vssd1 vccd1 vccd1 _3095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2115_ _2980_/X _2821_/X vssd1 vssd1 vccd1 vccd1 _2171_/A sky130_fd_sc_hd__nand2_2
X_2046_ _2313_/B _2971_/X _2045_/X vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _2373_/Y _2018_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__mux2_1
X_2879_ _2464_/Y _1787_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2802_ _2802_/A0 _3142_/Q _3186_/Q vssd1 vssd1 vccd1 vccd1 _2802_/X sky130_fd_sc_hd__mux2_1
X_2733_ _2403_/Y _2732_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__mux2_2
X_2664_ _2664_/A vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__clkbuf_1
X_1615_ _3163_/Q _1613_/X _1583_/X _1614_/X vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__o211a_1
X_2595_ _3177_/Q _1544_/B _2591_/Y _2594_/Y vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__a211o_1
XFILLER_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1546_ _2542_/A vssd1 vssd1 vccd1 vccd1 _1558_/B sky130_fd_sc_hd__buf_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1477_ _1611_/C vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__buf_2
XFILLER_86_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3147_ _3201_/CLK _3147_/D vssd1 vssd1 vccd1 vccd1 _3147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ _3166_/CLK _3078_/D vssd1 vssd1 vccd1 vccd1 _3078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2029_ _3065_/Q _2737_/X _2031_/S vssd1 vssd1 vccd1 vccd1 _3065_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2380_ _3070_/Q vssd1 vssd1 vccd1 vccd1 _2380_/Y sky130_fd_sc_hd__inv_2
Xinput6 io_dat_i[11] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
X_3001_ _2345_/Y _1923_/Y _2346_/Y _2347_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _3001_/X sky130_fd_sc_hd__mux4_2
XFILLER_24_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2716_ _2716_/A vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__clkbuf_2
X_2647_ _3027_/Q vssd1 vssd1 vccd1 vccd1 _2647_/Y sky130_fd_sc_hd__inv_2
Xoutput310 _2667_/X vssd1 vssd1 vccd1 vccd1 io_wo[7] sky130_fd_sc_hd__clkbuf_2
X_2578_ _3206_/Q _2610_/B _2626_/C vssd1 vssd1 vccd1 vccd1 _2578_/Y sky130_fd_sc_hd__nand3_2
X_1529_ _3189_/Q _1522_/X _1525_/X _1528_/Y vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _3095_/Q _2769_/X _1880_/S vssd1 vssd1 vccd1 vccd1 _3095_/D sky130_fd_sc_hd__mux2_1
XFILLER_41_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2501_ _3133_/Q vssd1 vssd1 vccd1 vccd1 _2501_/Y sky130_fd_sc_hd__inv_2
X_2432_ _3081_/Q vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2363_ _2363_/A vssd1 vssd1 vccd1 vccd1 _2363_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2294_ _3038_/Q vssd1 vssd1 vccd1 vccd1 _2294_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput162 _2617_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput173 _2595_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput195 _3119_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput184 _3022_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2981_ _2434_/Y _2090_/Y _2012_/Y _1863_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2981_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1932_ _1936_/B _1936_/A vssd1 vssd1 vccd1 vccd1 _1932_/Y sky130_fd_sc_hd__nand2_1
X_1863_ _3104_/Q vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__inv_2
Xinput20 io_eo[0] vssd1 vssd1 vccd1 vccd1 _2660_/A sky130_fd_sc_hd__clkbuf_2
Xinput31 io_eo[1] vssd1 vssd1 vccd1 vccd1 _2661_/A sky130_fd_sc_hd__clkbuf_2
X_1794_ _3119_/Q vssd1 vssd1 vccd1 vccd1 _1794_/Y sky130_fd_sc_hd__inv_2
Xinput64 io_eo[4] vssd1 vssd1 vccd1 vccd1 _2664_/A sky130_fd_sc_hd__clkbuf_2
Xinput42 io_eo[2] vssd1 vssd1 vccd1 vccd1 _2662_/A sky130_fd_sc_hd__clkbuf_2
Xinput53 io_eo[3] vssd1 vssd1 vccd1 vccd1 _2663_/A sky130_fd_sc_hd__clkbuf_2
Xinput97 io_i_1_in1[3] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
Xinput86 io_i_0_in1[1] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput75 io_eo[5] vssd1 vssd1 vccd1 vccd1 _2665_/A sky130_fd_sc_hd__clkbuf_2
X_2415_ _2427_/A _2763_/X vssd1 vssd1 vccd1 vccd1 _2415_/Y sky130_fd_sc_hd__nand2_1
X_2346_ _3108_/Q vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__inv_2
X_2277_ _2801_/X _2874_/X vssd1 vssd1 vccd1 vccd1 _2279_/A sky130_fd_sc_hd__nor2_2
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2200_ _2839_/X _3010_/X vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__and2b_1
X_3180_ _3197_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2131_ _2984_/X _2811_/X vssd1 vssd1 vccd1 vccd1 _2153_/A sky130_fd_sc_hd__xor2_4
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2062_ _2062_/A _2532_/A vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _2328_/Y _2097_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__mux2_1
X_1915_ _1912_/Y _1913_/X _1937_/S vssd1 vssd1 vccd1 vccd1 _1915_/Y sky130_fd_sc_hd__o21bai_1
X_2895_ _2448_/Y _2894_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2895_/X sky130_fd_sc_hd__mux2_1
X_1846_ _1844_/Y _1845_/X _1848_/A vssd1 vssd1 vccd1 vccd1 _1846_/Y sky130_fd_sc_hd__o21bai_1
X_1777_ _1777_/A _1874_/S vssd1 vssd1 vccd1 vccd1 _1777_/Y sky130_fd_sc_hd__nand2_1
X_2329_ _3182_/Q vssd1 vssd1 vccd1 vccd1 _2329_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1700_ _1699_/X _3137_/Q _2290_/S vssd1 vssd1 vccd1 vccd1 _3137_/D sky130_fd_sc_hd__mux2_1
X_2680_ _2680_/A vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__clkbuf_1
X_1631_ _1636_/A _1631_/B vssd1 vssd1 vccd1 vccd1 _1631_/Y sky130_fd_sc_hd__nand2_1
X_1562_ _3179_/Q _1556_/X _1557_/X _1561_/Y vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__o211a_1
X_1493_ _3200_/Q _1479_/X _1490_/X _1492_/Y vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__o211a_1
X_3163_ _3193_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_4
X_2114_ _2981_/X _2817_/X vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__and2_1
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3094_ _3211_/CLK _3094_/D vssd1 vssd1 vccd1 vccd1 _3094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2045_ _2313_/B _2971_/X _2990_/X _2969_/X vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__a211o_1
X_2947_ _3004_/A3 _3110_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__mux2_1
X_2878_ _2878_/A0 _3135_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__mux2_2
X_1829_ _2761_/X _2916_/X _2759_/X _2913_/X vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__a211oi_4
XFILLER_89_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2801_ _2470_/Y _2800_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2801_/X sky130_fd_sc_hd__mux2_2
X_2732_ _1794_/Y _2261_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _2663_/A vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__clkbuf_1
X_1614_ _1614_/A _2658_/B vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__or2b_1
X_2594_ _2594_/A _2594_/B vssd1 vssd1 vccd1 vccd1 _2594_/Y sky130_fd_sc_hd__nand2_1
X_1545_ _3185_/Q _1540_/X _1541_/X _1544_/Y vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1476_ _1500_/A vssd1 vssd1 vccd1 vccd1 _1611_/C sky130_fd_sc_hd__clkbuf_2
X_3146_ _3197_/CLK _3146_/D vssd1 vssd1 vccd1 vccd1 _3146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _3092_/CLK _3077_/D vssd1 vssd1 vccd1 vccd1 _3077_/Q sky130_fd_sc_hd__dfxtp_1
X_2028_ _3066_/Q _2393_/B _2031_/S vssd1 vssd1 vccd1 vccd1 _3066_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 io_dat_i[12] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
X_3000_ _2352_/Y _2304_/Y _2353_/Y _2354_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _3000_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _2715_/A vssd1 vssd1 vccd1 vccd1 _2715_/X sky130_fd_sc_hd__clkbuf_2
Xoutput300 _2716_/X vssd1 vssd1 vccd1 vccd1 io_wo[56] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2646_ _2646_/A _2984_/X vssd1 vssd1 vccd1 vccd1 _2646_/Y sky130_fd_sc_hd__nand2_1
Xoutput311 _2668_/X vssd1 vssd1 vccd1 vccd1 io_wo[8] sky130_fd_sc_hd__clkbuf_2
X_2577_ _2593_/B _3190_/Q _2618_/C vssd1 vssd1 vccd1 vccd1 _2577_/Y sky130_fd_sc_hd__nand3b_4
X_1528_ _1518_/X _1530_/B _1629_/B vssd1 vssd1 vccd1 vccd1 _1528_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_19_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1459_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1459_/X sky130_fd_sc_hd__buf_2
XFILLER_19_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3129_ _3139_/CLK _3129_/D vssd1 vssd1 vccd1 vccd1 _3129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2500_ _2500_/A _2506_/B vssd1 vssd1 vccd1 vccd1 _2500_/Y sky130_fd_sc_hd__nand2_1
X_2431_ _2439_/A _2755_/X vssd1 vssd1 vccd1 vccd1 _2431_/Y sky130_fd_sc_hd__nand2_1
X_2362_ _3050_/Q vssd1 vssd1 vccd1 vccd1 _2362_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2293_ _2313_/A _2995_/X vssd1 vssd1 vccd1 vccd1 _2293_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2629_ _1595_/Y _2608_/X _2626_/Y _2627_/Y _2628_/Y vssd1 vssd1 vccd1 vccd1 _2629_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput163 _2621_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput174 _2601_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput185 _2539_/Y vssd1 vssd1 vccd1 vccd1 io_o_1_co sky130_fd_sc_hd__clkbuf_2
Xoutput196 _3120_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _2438_/Y _2097_/Y _2018_/Y _1870_/Y _3168_/Q _3169_/Q vssd1 vssd1 vccd1 vccd1
+ _2980_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1931_ _1930_/X _3091_/Q _1937_/S vssd1 vssd1 vccd1 vccd1 _3091_/D sky130_fd_sc_hd__mux2_1
X_1862_ _1861_/X _3105_/Q _1862_/S vssd1 vssd1 vccd1 vccd1 _3105_/D sky130_fd_sc_hd__mux2_1
Xinput10 io_dat_i[15] vssd1 vssd1 vccd1 vccd1 _1593_/A sky130_fd_sc_hd__buf_2
Xinput21 io_eo[10] vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__clkbuf_2
X_1793_ _1791_/Y _1732_/Y _1731_/Y _1786_/S vssd1 vssd1 vccd1 vccd1 _1793_/Y sky130_fd_sc_hd__a31oi_1
Xinput32 io_eo[20] vssd1 vssd1 vccd1 vccd1 _2680_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 io_eo[30] vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__clkbuf_2
Xinput54 io_eo[40] vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__clkbuf_2
Xinput76 io_eo[60] vssd1 vssd1 vccd1 vccd1 _2720_/A sky130_fd_sc_hd__clkbuf_1
Xinput87 io_i_0_in1[2] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput98 io_i_1_in1[4] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
Xinput65 io_eo[50] vssd1 vssd1 vccd1 vccd1 _2710_/A sky130_fd_sc_hd__clkbuf_1
X_2414_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2414_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2345_ _2345_/A vssd1 vssd1 vccd1 vccd1 _2345_/Y sky130_fd_sc_hd__inv_2
X_2276_ _2284_/A vssd1 vssd1 vccd1 vccd1 _2521_/B sky130_fd_sc_hd__inv_2
XFILLER_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2130_ _2163_/B _2127_/Y _2129_/Y vssd1 vssd1 vccd1 vccd1 _2133_/A sky130_fd_sc_hd__a21bo_1
XFILLER_19_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _2995_/X _2979_/X vssd1 vssd1 vccd1 vccd1 _2532_/A sky130_fd_sc_hd__and2_1
XFILLER_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2963_ _2337_/Y _2962_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__mux2_2
X_1914_ _2731_/X vssd1 vssd1 vccd1 vccd1 _1937_/S sky130_fd_sc_hd__inv_2
X_2894_ _2449_/Y _1766_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__mux2_1
X_1845_ _1845_/A _1845_/B _1845_/C vssd1 vssd1 vccd1 vccd1 _1845_/X sky130_fd_sc_hd__and3_1
X_1776_ _2767_/X vssd1 vssd1 vccd1 vccd1 _1874_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2328_ _3031_/Q vssd1 vssd1 vccd1 vccd1 _2328_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2259_ _2257_/Y _2196_/Y _2258_/Y vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _3157_/Q _1626_/X _1623_/X _1629_/Y vssd1 vssd1 vccd1 vccd1 _3157_/D sky130_fd_sc_hd__o211a_1
X_1561_ _1551_/X _1572_/B _2658_/B vssd1 vssd1 vccd1 vccd1 _1561_/Y sky130_fd_sc_hd__nand3b_1
X_1492_ _1609_/B _1498_/B _1653_/B vssd1 vssd1 vccd1 vccd1 _1492_/Y sky130_fd_sc_hd__nand3b_1
X_3162_ _3193_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_4
X_2113_ _2132_/B _2111_/Y _2132_/A vssd1 vssd1 vccd1 vccd1 _2113_/Y sky130_fd_sc_hd__o21bai_1
X_3093_ _3211_/CLK _3093_/D vssd1 vssd1 vccd1 vccd1 _3093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2044_ _2044_/A _2044_/B vssd1 vssd1 vccd1 vccd1 _2086_/A sky130_fd_sc_hd__nor2_2
XFILLER_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2946_ _2379_/Y _2945_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__mux2_2
XFILLER_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2877_ _2466_/Y _2876_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__mux2_2
X_1828_ _1843_/A vssd1 vssd1 vccd1 vccd1 _1831_/B sky130_fd_sc_hd__inv_2
X_1759_ _1759_/A _2524_/A vssd1 vssd1 vccd1 vccd1 _1759_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ _2409_/Y _2331_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2800_/X sky130_fd_sc_hd__mux2_1
X_2731_ _2349_/Y _2730_/X _3195_/Q vssd1 vssd1 vccd1 vccd1 _2731_/X sky130_fd_sc_hd__mux2_2
XFILLER_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2662_ _2662_/A vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1613_ _1636_/A vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__clkbuf_2
X_2593_ _3209_/Q _2593_/B _2593_/C vssd1 vssd1 vccd1 vccd1 _2594_/B sky130_fd_sc_hd__nand3_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_1544_ _1532_/X _1544_/B _1650_/B vssd1 vssd1 vccd1 vccd1 _1544_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1475_ input2/X vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__inv_2
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3145_ _3193_/CLK _3145_/D vssd1 vssd1 vccd1 vccd1 _3145_/Q sky130_fd_sc_hd__dfxtp_1
X_3076_ _3092_/CLK _3076_/D vssd1 vssd1 vccd1 vccd1 _3076_/Q sky130_fd_sc_hd__dfxtp_1
X_2027_ _3067_/Q _2741_/X _2031_/S vssd1 vssd1 vccd1 vccd1 _3067_/D sky130_fd_sc_hd__mux2_1
X_2929_ _3010_/A3 _3104_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 io_dat_i[13] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_76_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _2714_/A vssd1 vssd1 vccd1 vccd1 _2714_/X sky130_fd_sc_hd__clkbuf_2
Xoutput301 _2717_/X vssd1 vssd1 vccd1 vccd1 io_wo[57] sky130_fd_sc_hd__clkbuf_2
X_2645_ _3042_/Q vssd1 vssd1 vccd1 vccd1 _2645_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput312 _2669_/X vssd1 vssd1 vccd1 vccd1 io_wo[9] sky130_fd_sc_hd__clkbuf_2
X_2576_ _2603_/C vssd1 vssd1 vccd1 vccd1 _2618_/C sky130_fd_sc_hd__buf_4
X_1527_ _3190_/Q _1522_/X _1525_/X _1526_/Y vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1458_ _2658_/A vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3128_ _3139_/CLK _3128_/D vssd1 vssd1 vccd1 vccd1 _3128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3059_ _3075_/CLK _3059_/D vssd1 vssd1 vccd1 vccd1 _3059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2430_/Y sky130_fd_sc_hd__inv_2
X_2361_ _2361_/A _2361_/B vssd1 vssd1 vccd1 vccd1 _2361_/Y sky130_fd_sc_hd__nand2_1
X_2292_ _2327_/A vssd1 vssd1 vccd1 vccd1 _2313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2628_ _2611_/X _3184_/Q _2630_/C vssd1 vssd1 vccd1 vccd1 _2628_/Y sky130_fd_sc_hd__nand3b_2
Xoutput164 _2625_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput175 _2607_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput186 _3135_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[0] sky130_fd_sc_hd__clkbuf_2
X_2559_ _2598_/A vssd1 vssd1 vccd1 vccd1 _2631_/C sky130_fd_sc_hd__buf_2
Xoutput197 _3121_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1930_ _1930_/A _1930_/B vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__xor2_1
X_1861_ _1861_/A _1861_/B vssd1 vssd1 vccd1 vccd1 _1861_/X sky130_fd_sc_hd__xor2_1
Xinput11 io_dat_i[1] vssd1 vssd1 vccd1 vccd1 _1467_/A sky130_fd_sc_hd__clkbuf_1
Xinput22 io_eo[11] vssd1 vssd1 vccd1 vccd1 _2671_/A sky130_fd_sc_hd__clkbuf_2
X_1792_ _1791_/Y _1731_/Y _1732_/Y vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__a21o_1
Xinput33 io_eo[21] vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__clkbuf_2
Xinput44 io_eo[31] vssd1 vssd1 vccd1 vccd1 _2691_/A sky130_fd_sc_hd__clkbuf_2
Xinput55 io_eo[41] vssd1 vssd1 vccd1 vccd1 _2701_/A sky130_fd_sc_hd__clkbuf_2
Xinput77 io_eo[61] vssd1 vssd1 vccd1 vccd1 _2721_/A sky130_fd_sc_hd__clkbuf_1
Xinput66 io_eo[51] vssd1 vssd1 vccd1 vccd1 _2711_/A sky130_fd_sc_hd__clkbuf_1
Xinput88 io_i_0_in1[3] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput99 io_i_1_in1[5] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
X_2413_ _2920_/X vssd1 vssd1 vccd1 vccd1 _2413_/Y sky130_fd_sc_hd__inv_2
X_2344_ _3053_/Q vssd1 vssd1 vccd1 vccd1 _2344_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2275_ _2799_/X _2871_/X vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _2995_/X _2979_/X vssd1 vssd1 vccd1 vccd1 _2062_/A sky130_fd_sc_hd__nor2_4
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2962_ _2338_/Y _1956_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__mux2_1
X_1913_ _2528_/A _1911_/A _1908_/Y _1906_/Y vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__o211a_1
X_2893_ _2893_/A0 _3012_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__mux2_1
X_1844_ _1845_/A _1845_/B _1845_/C vssd1 vssd1 vccd1 vccd1 _1844_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1775_ _1775_/A _1775_/B vssd1 vssd1 vccd1 vccd1 _1777_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2327_ _2327_/A _2988_/X vssd1 vssd1 vccd1 vccd1 _2327_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2258_ _2835_/X vssd1 vssd1 vccd1 vccd1 _2258_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2189_ _3026_/Q _2983_/X _2190_/S vssd1 vssd1 vccd1 vccd1 _3026_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3110_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ _2542_/A vssd1 vssd1 vccd1 vccd1 _1572_/B sky130_fd_sc_hd__buf_1
X_1491_ input9/X vssd1 vssd1 vccd1 vccd1 _1653_/B sky130_fd_sc_hd__inv_2
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3161_ _3193_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_4
X_2112_ _2985_/X _2809_/X vssd1 vssd1 vccd1 vccd1 _2132_/A sky130_fd_sc_hd__nor2_2
X_3092_ _3092_/CLK _3092_/D vssd1 vssd1 vccd1 vccd1 _3092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2043_ _2991_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _2044_/B sky130_fd_sc_hd__and2_1
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2945_ _2380_/Y _1881_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__mux2_1
X_2876_ _2467_/Y _1794_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2876_/X sky130_fd_sc_hd__mux2_1
X_1827_ _2763_/X _2919_/X vssd1 vssd1 vccd1 vccd1 _1843_/A sky130_fd_sc_hd__nor2_1
X_1758_ _2783_/X _2898_/X vssd1 vssd1 vccd1 vccd1 _2524_/A sky130_fd_sc_hd__and2_1
X_1689_ _2484_/B _2862_/X _1688_/X vssd1 vssd1 vccd1 vccd1 _1689_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2730_ _2749_/X _3146_/Q _3194_/Q vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__mux2_1
X_2661_ _2661_/A vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__clkbuf_1
X_1612_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1636_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2592_ _2548_/A _3193_/Q _2593_/C vssd1 vssd1 vccd1 vccd1 _2594_/A sky130_fd_sc_hd__nand3b_1
X_1543_ _2542_/A vssd1 vssd1 vccd1 vccd1 _1544_/B sky130_fd_sc_hd__clkbuf_2
X_1474_ input1/X vssd1 vssd1 vccd1 vccd1 _2605_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3189_/CLK _3144_/D vssd1 vssd1 vccd1 vccd1 _3144_/Q sky130_fd_sc_hd__dfxtp_1
X_3075_ _3075_/CLK _3075_/D vssd1 vssd1 vccd1 vccd1 _3075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2026_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2031_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _2401_/Y _2927_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2859_ _2487_/Y _2858_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__mux2_2
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 io_dat_i[14] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _2713_/A vssd1 vssd1 vccd1 vccd1 _2713_/X sky130_fd_sc_hd__clkbuf_2
X_2644_ _3026_/Q vssd1 vssd1 vccd1 vccd1 _2644_/Y sky130_fd_sc_hd__inv_2
Xoutput302 _2718_/X vssd1 vssd1 vccd1 vccd1 io_wo[58] sky130_fd_sc_hd__clkbuf_2
X_2575_ _3173_/Q _1544_/B _2571_/Y _2574_/Y vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__a211o_1
X_1526_ _1518_/X _1530_/B _1627_/B vssd1 vssd1 vccd1 vccd1 _1526_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_19_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1457_ _2466_/A _1435_/X _1438_/X _1456_/Y vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3127_ _3139_/CLK _3127_/D vssd1 vssd1 vccd1 vccd1 _3127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3058_ _3075_/CLK _3058_/D vssd1 vssd1 vccd1 vccd1 _3058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _2008_/Y _3074_/Q _2011_/S vssd1 vssd1 vccd1 vccd1 _3074_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2360_ _3138_/Q vssd1 vssd1 vccd1 vccd1 _2360_/Y sky130_fd_sc_hd__inv_2
X_2291_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2291_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2627_ _3148_/Q _2627_/B _2627_/C vssd1 vssd1 vccd1 vccd1 _2627_/Y sky130_fd_sc_hd__nand3_2
Xoutput165 _2629_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput176 _2540_/Y vssd1 vssd1 vccd1 vccd1 io_o_0_co sky130_fd_sc_hd__clkbuf_2
X_2558_ _2632_/B _2616_/C _3155_/Q vssd1 vssd1 vccd1 vccd1 _2558_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1509_ _3196_/Q _1506_/X _1490_/X _1508_/Y vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__o211a_1
X_2489_ _2857_/X vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__inv_2
Xoutput187 _3136_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput198 _3122_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _1859_/Y _3106_/Q _1862_/S vssd1 vssd1 vccd1 vccd1 _3106_/D sky130_fd_sc_hd__mux2_1
Xinput12 io_dat_i[2] vssd1 vssd1 vccd1 vccd1 _1464_/A sky130_fd_sc_hd__buf_1
X_1791_ _1791_/A vssd1 vssd1 vccd1 vccd1 _1791_/Y sky130_fd_sc_hd__inv_2
Xinput23 io_eo[12] vssd1 vssd1 vccd1 vccd1 _2672_/A sky130_fd_sc_hd__clkbuf_2
Xinput34 io_eo[22] vssd1 vssd1 vccd1 vccd1 _2682_/A sky130_fd_sc_hd__clkbuf_2
Xinput45 io_eo[32] vssd1 vssd1 vccd1 vccd1 _2692_/A sky130_fd_sc_hd__clkbuf_2
Xinput78 io_eo[62] vssd1 vssd1 vccd1 vccd1 _2722_/A sky130_fd_sc_hd__clkbuf_1
Xinput67 io_eo[52] vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__clkbuf_1
Xinput89 io_i_0_in1[4] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput56 io_eo[42] vssd1 vssd1 vccd1 vccd1 _2702_/A sky130_fd_sc_hd__clkbuf_2
X_2412_ _3086_/Q vssd1 vssd1 vccd1 vccd1 _2412_/Y sky130_fd_sc_hd__inv_2
X_2343_ _2361_/A _3002_/X vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__nand2_1
X_2274_ _2285_/B _2274_/B vssd1 vssd1 vccd1 vccd1 _2521_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1989_ _2729_/X vssd1 vssd1 vccd1 vccd1 _2011_/S sky130_fd_sc_hd__inv_2
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2961_ _2343_/Y _2960_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__mux2_1
X_1912_ _1906_/Y _1908_/Y _1911_/Y vssd1 vssd1 vccd1 vccd1 _1912_/Y sky130_fd_sc_hd__a21boi_1
X_2892_ _2451_/Y _2891_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__mux2_2
X_1843_ _1843_/A _1843_/B vssd1 vssd1 vccd1 vccd1 _1845_/C sky130_fd_sc_hd__nor2_1
X_1774_ _1779_/B _1779_/A _1773_/Y vssd1 vssd1 vccd1 vccd1 _1775_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2326_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2326_/Y sky130_fd_sc_hd__inv_2
X_2257_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2188_ _3027_/Q _2984_/X _2190_/S vssd1 vssd1 vccd1 vccd1 _3027_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1490_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__buf_1
X_3160_ _3193_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_4
X_2111_ _2111_/A vssd1 vssd1 vccd1 vccd1 _2111_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3091_ _3092_/CLK _3091_/D vssd1 vssd1 vccd1 vccd1 _3091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2042_ _2313_/B _2971_/X vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2944_ _3005_/A3 _3109_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2944_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2875_ _2875_/A0 _3022_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__mux2_1
X_1826_ _1855_/B _1855_/A _1851_/A vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__nand3_4
X_1757_ _2783_/X _2898_/X vssd1 vssd1 vccd1 vccd1 _1759_/A sky130_fd_sc_hd__nor2_4
X_1688_ _2484_/B _2862_/X _2791_/X _2859_/X vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__a211o_1
X_2309_ _3074_/Q vssd1 vssd1 vccd1 vccd1 _2309_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2660_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1611_ input1/X input2/X _1611_/C vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__nor3_4
X_2591_ _2620_/C _2616_/C _3161_/Q vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1542_ _2611_/A _2596_/A vssd1 vssd1 vccd1 vccd1 _2542_/A sky130_fd_sc_hd__nor2b_4
X_1473_ _2550_/A _1458_/X _1459_/X _1472_/Y vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__o211a_1
X_3143_ _3189_/CLK _3143_/D vssd1 vssd1 vccd1 vccd1 _3143_/Q sky130_fd_sc_hd__dfxtp_1
X_3074_ _3074_/CLK _3074_/D vssd1 vssd1 vccd1 vccd1 _3074_/Q sky130_fd_sc_hd__dfxtp_1
X_2025_ _3068_/Q _2743_/X _2025_/S vssd1 vssd1 vccd1 vccd1 _3068_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ _2402_/Y _1938_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2927_/X sky130_fd_sc_hd__mux2_1
X_2858_ _2488_/Y _2365_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__mux2_1
X_2789_ _2489_/Y _2788_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__mux2_2
X_1809_ _2829_/X vssd1 vssd1 vccd1 vccd1 _1809_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2643_ _2646_/A _2983_/X vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__nand2_1
Xoutput303 _2719_/X vssd1 vssd1 vccd1 vccd1 io_wo[59] sky130_fd_sc_hd__clkbuf_2
X_2574_ _2574_/A _2574_/B vssd1 vssd1 vccd1 vccd1 _2574_/Y sky130_fd_sc_hd__nand2_1
X_1525_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1525_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1456_ _1472_/A _1627_/B vssd1 vssd1 vccd1 vccd1 _1456_/Y sky130_fd_sc_hd__nand2_1
X_3126_ _3209_/CLK _3126_/D vssd1 vssd1 vccd1 vccd1 _3126_/Q sky130_fd_sc_hd__dfxtp_2
X_3057_ _3075_/CLK _3057_/D vssd1 vssd1 vccd1 vccd1 _3057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2008_ _2008_/A _2008_/B vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_50_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2290_ _2289_/X _3012_/Q _2290_/S vssd1 vssd1 vccd1 vccd1 _3012_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2626_ _2596_/X _3200_/Q _2626_/C vssd1 vssd1 vccd1 vccd1 _2626_/Y sky130_fd_sc_hd__nand3b_4
Xoutput166 _2633_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput177 _3015_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[0] sky130_fd_sc_hd__clkbuf_2
X_2557_ _2603_/C vssd1 vssd1 vccd1 vccd1 _2616_/C sky130_fd_sc_hd__clkbuf_4
Xoutput188 _3137_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[2] sky130_fd_sc_hd__clkbuf_2
X_2488_ _3113_/Q vssd1 vssd1 vccd1 vccd1 _2488_/Y sky130_fd_sc_hd__inv_2
Xoutput199 _3123_/Q vssd1 vssd1 vccd1 vccd1 io_o_2_out[4] sky130_fd_sc_hd__clkbuf_2
X_1508_ _1501_/X _1516_/B _1643_/B vssd1 vssd1 vccd1 vccd1 _1508_/Y sky130_fd_sc_hd__nand3b_1
X_1439_ _1638_/A vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__buf_1
X_3109_ _3110_/CLK _3109_/D vssd1 vssd1 vccd1 vccd1 _3109_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 io_dat_i[3] vssd1 vssd1 vccd1 vccd1 _1460_/A sky130_fd_sc_hd__buf_1
X_1790_ _1874_/S _1787_/Y _1788_/X _1789_/Y vssd1 vssd1 vccd1 vccd1 _3120_/D sky130_fd_sc_hd__o22ai_1
Xinput24 io_eo[13] vssd1 vssd1 vccd1 vccd1 _2673_/A sky130_fd_sc_hd__clkbuf_2
Xinput35 io_eo[23] vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__clkbuf_2
Xinput46 io_eo[33] vssd1 vssd1 vccd1 vccd1 _2693_/A sky130_fd_sc_hd__clkbuf_2
Xinput79 io_eo[63] vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__clkbuf_1
Xinput68 io_eo[53] vssd1 vssd1 vccd1 vccd1 _2713_/A sky130_fd_sc_hd__clkbuf_1
Xinput57 io_eo[43] vssd1 vssd1 vccd1 vccd1 _2703_/A sky130_fd_sc_hd__clkbuf_2
X_2411_ _2427_/A _2765_/X vssd1 vssd1 vccd1 vccd1 _2411_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2342_ _2348_/A _3190_/Q vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__nand2_1
X_2273_ _2284_/B vssd1 vssd1 vccd1 vccd1 _2274_/B sky130_fd_sc_hd__inv_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1988_ _2530_/A _1986_/A _1983_/Y _1981_/Y vssd1 vssd1 vccd1 vccd1 _1988_/X sky130_fd_sc_hd__o211a_1
X_2609_ _2596_/X _3196_/Q _2618_/C vssd1 vssd1 vccd1 vccd1 _2609_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _2344_/Y _1992_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__mux2_1
X_2891_ _2452_/Y _1772_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2891_/X sky130_fd_sc_hd__mux2_1
X_1911_ _1911_/A _2528_/A vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1842_ _3109_/Q vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__inv_2
X_1773_ _2777_/X _2889_/X vssd1 vssd1 vccd1 vccd1 _1773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2325_ _3032_/Q vssd1 vssd1 vccd1 vccd1 _2325_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2256_ _2253_/Y _2254_/Y _2244_/B _2255_/X vssd1 vssd1 vccd1 vccd1 _3016_/D sky130_fd_sc_hd__a31o_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2187_ _3028_/Q _2985_/X _2190_/S vssd1 vssd1 vccd1 vccd1 _3028_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2110_ _2984_/X _2811_/X vssd1 vssd1 vccd1 vccd1 _2111_/A sky130_fd_sc_hd__nor2_1
X_3090_ _3110_/CLK _3090_/D vssd1 vssd1 vccd1 vccd1 _3090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2041_ _2991_/X vssd1 vssd1 vccd1 vccd1 _2313_/B sky130_fd_sc_hd__buf_1
XFILLER_81_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2943_ _2383_/Y _2942_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2943_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2874_ _2472_/Y _2873_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__mux2_1
X_1825_ _1830_/A _1825_/B vssd1 vssd1 vccd1 vccd1 _1851_/A sky130_fd_sc_hd__nor2_4
X_1756_ _1767_/B vssd1 vssd1 vccd1 vccd1 _1756_/Y sky130_fd_sc_hd__inv_2
X_1687_ _1687_/A _1687_/B vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__nor2_4
X_2308_ _3035_/Q vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2239_ _2504_/A _2845_/X _2221_/Y _2244_/C vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__o211a_1
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1610_ _1614_/A _1608_/Y _1655_/A _1609_/Y vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__a211oi_1
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2441_/Y _2542_/Y _2587_/Y _2588_/Y _2589_/Y vssd1 vssd1 vccd1 vccd1 _2590_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_1541_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1472_ _1472_/A _1636_/B vssd1 vssd1 vccd1 vccd1 _1472_/Y sky130_fd_sc_hd__nand2_1
X_3211_ _3211_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3142_ _3189_/CLK _3142_/D vssd1 vssd1 vccd1 vccd1 _3142_/Q sky130_fd_sc_hd__dfxtp_1
X_3073_ _3074_/CLK _3073_/D vssd1 vssd1 vccd1 vccd1 _3073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2024_ _3069_/Q _2745_/X _2025_/S vssd1 vssd1 vccd1 vccd1 _3069_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2926_ _3011_/A3 _3103_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2926_/X sky130_fd_sc_hd__mux2_2
X_2857_ input95/X _3016_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__mux2_1
X_1808_ _2751_/X _2901_/X vssd1 vssd1 vccd1 vccd1 _1808_/Y sky130_fd_sc_hd__nand2_2
X_2788_ _2434_/Y _2368_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__mux2_1
X_1739_ _2457_/B _2886_/X vssd1 vssd1 vccd1 vccd1 _1741_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2711_ _2711_/A vssd1 vssd1 vccd1 vccd1 _2711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _3041_/Q vssd1 vssd1 vccd1 vccd1 _2642_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput304 _2665_/X vssd1 vssd1 vccd1 vccd1 io_wo[5] sky130_fd_sc_hd__clkbuf_2
X_2573_ _3205_/Q _2627_/B _2593_/C vssd1 vssd1 vccd1 vccd1 _2574_/B sky130_fd_sc_hd__nand3_1
X_1524_ _3191_/Q _1522_/X _1510_/X _1523_/Y vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__o211a_1
X_1455_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1627_/B sky130_fd_sc_hd__inv_2
X_3125_ _3209_/CLK _3125_/D vssd1 vssd1 vccd1 vccd1 _3125_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _3074_/CLK _3056_/D vssd1 vssd1 vccd1 vccd1 _3056_/Q sky130_fd_sc_hd__dfxtp_1
X_2007_ _2998_/X _2953_/X _2006_/Y vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__o21a_1
X_2909_ _2428_/Y _2359_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2625_ _1598_/Y _2608_/X _2622_/Y _2623_/Y _2624_/Y vssd1 vssd1 vccd1 vccd1 _2625_/Y
+ sky130_fd_sc_hd__o2111ai_4
Xoutput167 _2565_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[1] sky130_fd_sc_hd__clkbuf_2
X_2556_ _2603_/B vssd1 vssd1 vccd1 vccd1 _2632_/B sky130_fd_sc_hd__clkbuf_4
X_2487_ _2493_/A _2791_/X vssd1 vssd1 vccd1 vccd1 _2487_/Y sky130_fd_sc_hd__nand2_1
Xoutput178 _3016_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput189 _3138_/Q vssd1 vssd1 vccd1 vccd1 io_o_1_out[3] sky130_fd_sc_hd__clkbuf_2
X_1507_ input5/X vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__inv_2
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1438_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__buf_1
X_3108_ _3122_/CLK _3108_/D vssd1 vssd1 vccd1 vccd1 _3108_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3039_ _3201_/CLK _3039_/D vssd1 vssd1 vccd1 vccd1 _3039_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_dat_i[4] vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 io_eo[14] vssd1 vssd1 vccd1 vccd1 _2674_/A sky130_fd_sc_hd__clkbuf_2
Xinput36 io_eo[24] vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 io_eo[54] vssd1 vssd1 vccd1 vccd1 _2714_/A sky130_fd_sc_hd__clkbuf_1
Xinput47 io_eo[34] vssd1 vssd1 vccd1 vccd1 _2694_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 io_eo[44] vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__clkbuf_1
X_2410_ _2439_/A vssd1 vssd1 vccd1 vccd1 _2427_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2341_ _2348_/A _3192_/Q vssd1 vssd1 vccd1 vccd1 _2341_/Y sky130_fd_sc_hd__nand2_1
X_2272_ _2799_/X _2871_/X vssd1 vssd1 vccd1 vccd1 _2284_/B sky130_fd_sc_hd__and2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _1981_/Y _1983_/Y _1986_/Y vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__a21boi_1
X_2608_ _2608_/A vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__buf_4
X_2539_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2539_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _2890_/A0 _3139_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1910_ _2747_/X _2946_/X vssd1 vssd1 vccd1 vccd1 _2528_/A sky130_fd_sc_hd__and2_1
XFILLER_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1841_ _1659_/X _1806_/Y _1840_/Y vssd1 vssd1 vccd1 vccd1 _3110_/D sky130_fd_sc_hd__o21ai_1
X_1772_ _3124_/Q vssd1 vssd1 vccd1 vccd1 _1772_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2324_ _2327_/A _2989_/X vssd1 vssd1 vccd1 vccd1 _2324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2255_ _1728_/S _3016_/Q vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__and2b_1
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2186_ _3029_/Q _2986_/X _2190_/S vssd1 vssd1 vccd1 vccd1 _3029_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2990_/X _2969_/X vssd1 vssd1 vccd1 vccd1 _2088_/A sky130_fd_sc_hd__xor2_4
XFILLER_62_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _2384_/Y _1917_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2873_ _2473_/Y _2263_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__mux2_1
X_1824_ _2761_/X _2916_/X vssd1 vssd1 vccd1 vccd1 _1825_/B sky130_fd_sc_hd__and2_1
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1755_ _2781_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _1767_/B sky130_fd_sc_hd__and2_1
X_1686_ _2793_/X _2862_/X vssd1 vssd1 vccd1 vccd1 _1687_/B sky130_fd_sc_hd__and2_1
X_2307_ _3059_/Q vssd1 vssd1 vccd1 vccd1 _2307_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2238_ _2244_/C _2237_/Y _2221_/Y vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__a21oi_1
X_2169_ _2184_/S _2165_/Y _2166_/X _2168_/Y vssd1 vssd1 vccd1 vccd1 _3040_/D sky130_fd_sc_hd__o22ai_1
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1540_/X sky130_fd_sc_hd__clkbuf_2
X_1471_ input4/X vssd1 vssd1 vccd1 vccd1 _1636_/B sky130_fd_sc_hd__inv_2
X_3210_ _3211_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3141_ _3197_/CLK _3141_/D vssd1 vssd1 vccd1 vccd1 _3141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3072_ _3074_/CLK _3072_/D vssd1 vssd1 vccd1 vccd1 _3072_/Q sky130_fd_sc_hd__dfxtp_1
X_2023_ _3070_/Q _2747_/X _2025_/S vssd1 vssd1 vccd1 vccd1 _3070_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2925_ _2404_/Y _2924_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2925_/X sky130_fd_sc_hd__mux2_2
X_2856_ _2490_/Y _2855_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__mux2_1
X_1807_ _2753_/X _2904_/X vssd1 vssd1 vccd1 vccd1 _1807_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3123_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_2787_ _2492_/Y _2786_/X _3157_/Q vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__mux2_2
X_1738_ _2775_/X vssd1 vssd1 vccd1 vccd1 _2457_/B sky130_fd_sc_hd__buf_1
X_1669_ _2731_/X vssd1 vssd1 vccd1 vccd1 _2026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _2710_/A vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__clkbuf_2
X_2641_ _3025_/Q vssd1 vssd1 vccd1 vccd1 _2641_/Y sky130_fd_sc_hd__inv_2
Xoutput305 _2720_/X vssd1 vssd1 vccd1 vccd1 io_wo[60] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2572_ _2548_/A _3189_/Q _2631_/C vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__nand3b_1
X_1523_ _1518_/X _1530_/B _1624_/B vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__nand3b_1
X_1454_ _1638_/A vssd1 vssd1 vccd1 vccd1 _1472_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3124_ _3209_/CLK _3124_/D vssd1 vssd1 vccd1 vccd1 _3124_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3055_ _3075_/CLK _3055_/D vssd1 vssd1 vccd1 vccd1 _3055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2006_ _2010_/B _2010_/A vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2908_ _2908_/A0 _3121_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__mux2_1
X_2839_ _2510_/Y _2838_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2624_ _3151_/Q _2632_/B _2632_/C vssd1 vssd1 vccd1 vccd1 _2624_/Y sky130_fd_sc_hd__nand3_2
Xoutput168 _2570_/Y vssd1 vssd1 vccd1 vccd1 io_dat_o[2] sky130_fd_sc_hd__clkbuf_2
X_2555_ _2596_/A vssd1 vssd1 vccd1 vccd1 _2603_/B sky130_fd_sc_hd__buf_1
X_2486_ _2860_/X vssd1 vssd1 vccd1 vccd1 _2486_/Y sky130_fd_sc_hd__inv_2
Xoutput179 _3017_/Q vssd1 vssd1 vccd1 vccd1 io_o_0_out[2] sky130_fd_sc_hd__clkbuf_2
X_1506_ _1522_/A vssd1 vssd1 vccd1 vccd1 _1506_/X sky130_fd_sc_hd__clkbuf_2
X_1437_ _1488_/A vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__buf_1
XFILLER_87_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _3122_/CLK _3107_/D vssd1 vssd1 vccd1 vccd1 _3107_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _3166_/CLK _3038_/D vssd1 vssd1 vccd1 vccd1 _3038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 io_dat_i[5] vssd1 vssd1 vccd1 vccd1 _1450_/A sky130_fd_sc_hd__buf_1
Xinput26 io_eo[15] vssd1 vssd1 vccd1 vccd1 _2675_/A sky130_fd_sc_hd__clkbuf_2
Xinput37 io_eo[25] vssd1 vssd1 vccd1 vccd1 _2685_/A sky130_fd_sc_hd__clkbuf_2
Xinput48 io_eo[35] vssd1 vssd1 vccd1 vccd1 _2695_/A sky130_fd_sc_hd__clkbuf_2
Xinput59 io_eo[45] vssd1 vssd1 vccd1 vccd1 _2705_/A sky130_fd_sc_hd__clkbuf_1
X_2340_ _3013_/Q vssd1 vssd1 vccd1 vccd1 _2340_/Y sky130_fd_sc_hd__inv_2
X_2271_ _2268_/Y _1691_/B _2270_/Y vssd1 vssd1 vccd1 vccd1 _2285_/B sky130_fd_sc_hd__o21bai_2
XFILLER_69_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _1986_/A _2530_/A vssd1 vssd1 vccd1 vccd1 _1986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2607_ _1498_/B _3195_/Q _2602_/Y _2604_/Y _2606_/Y vssd1 vssd1 vccd1 vccd1 _2607_/X
+ sky130_fd_sc_hd__a2111o_1
X_2538_ _2538_/A vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__inv_2
X_2469_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2469_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1840_ _1837_/Y _1838_/X _1848_/A vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__o21bai_1
X_1771_ _1661_/X _1766_/Y _1770_/Y vssd1 vssd1 vccd1 vccd1 _3125_/D sky130_fd_sc_hd__o21ai_1
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2323_ _2323_/A vssd1 vssd1 vccd1 vccd1 _2323_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2254_ _2835_/X _2257_/A _2200_/X _2199_/A _2196_/Y vssd1 vssd1 vccd1 vccd1 _2254_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ _2192_/S vssd1 vssd1 vccd1 vccd1 _2190_/S sky130_fd_sc_hd__buf_2
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1969_ _2361_/B _2955_/X _2998_/X _2953_/X vssd1 vssd1 vccd1 vccd1 _1969_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2941_ _3006_/A3 _3108_/Q _3162_/Q vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__mux2_1
X_2872_ _2872_/A0 _3021_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _2761_/X _2916_/X vssd1 vssd1 vccd1 vccd1 _1830_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1754_ _1769_/A _1754_/B _1769_/B vssd1 vssd1 vccd1 vccd1 _1754_/Y sky130_fd_sc_hd__nand3_4
X_1685_ _2484_/B _2862_/X vssd1 vssd1 vccd1 vccd1 _1687_/A sky130_fd_sc_hd__nor2_2
X_2306_ _2313_/A _2992_/X vssd1 vssd1 vccd1 vccd1 _2306_/Y sky130_fd_sc_hd__nand2_1
X_2237_ _2237_/A vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _2119_/Y _2114_/X _2118_/Y _2192_/S vssd1 vssd1 vccd1 vccd1 _2168_/Y sky130_fd_sc_hd__o31ai_1
X_2099_ _3054_/Q _3003_/X _2102_/S vssd1 vssd1 vccd1 vccd1 _3054_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _3202_/Q vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__buf_2
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3140_ _3201_/CLK _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/Q sky130_fd_sc_hd__dfxtp_1
X_3071_ _3092_/CLK _3071_/D vssd1 vssd1 vccd1 vccd1 _3071_/Q sky130_fd_sc_hd__dfxtp_1
X_2022_ _2102_/S _2018_/Y _2020_/X _2021_/Y vssd1 vssd1 vccd1 vccd1 _3071_/D sky130_fd_sc_hd__o22ai_1
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2924_ _2405_/Y _1942_/Y _3210_/Q vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__mux2_1
X_2855_ _2491_/Y _1701_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__mux2_1
X_1806_ _3110_/Q vssd1 vssd1 vccd1 vccd1 _1806_/Y sky130_fd_sc_hd__inv_2
X_2786_ _2438_/Y _2371_/Y _3156_/Q vssd1 vssd1 vccd1 vccd1 _2786_/X sky130_fd_sc_hd__mux2_1
X_1737_ _2773_/X _2883_/X vssd1 vssd1 vccd1 vccd1 _1785_/A sky130_fd_sc_hd__xor2_2
X_1668_ _1673_/A _2802_/A0 vssd1 vssd1 vccd1 vccd1 _3142_/D sky130_fd_sc_hd__nor2b_1
X_1599_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1655_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ _2646_/A _2982_/X vssd1 vssd1 vccd1 vccd1 _2640_/Y sky130_fd_sc_hd__nand2_1
Xoutput306 _2721_/X vssd1 vssd1 vccd1 vccd1 io_wo[61] sky130_fd_sc_hd__clkbuf_2
X_2571_ _2632_/B _2616_/C _3157_/Q vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__nor3b_2
X_1522_ _1522_/A vssd1 vssd1 vccd1 vccd1 _1522_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1453_ _3206_/Q vssd1 vssd1 vccd1 vccd1 _2466_/A sky130_fd_sc_hd__clkbuf_2
X_3123_ _3123_/CLK _3123_/D vssd1 vssd1 vccd1 vccd1 _3123_/Q sky130_fd_sc_hd__dfxtp_2
X_3054_ _3211_/CLK _3054_/D vssd1 vssd1 vccd1 vccd1 _3054_/Q sky130_fd_sc_hd__dfxtp_1
X_2005_ _2003_/X _1998_/Y _1657_/X _2004_/X vssd1 vssd1 vccd1 vccd1 _3075_/D sky130_fd_sc_hd__a31o_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2907_ _2431_/Y _2906_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__mux2_2
X_2838_ _2511_/Y _2400_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__mux2_1
X_2769_ _2465_/Y _2768_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ _2603_/B _3199_/Q _2631_/C vssd1 vssd1 vccd1 vccd1 _2623_/Y sky130_fd_sc_hd__nand3b_2
X_2554_ _2514_/Y _2542_/Y _2546_/Y _2550_/Y _2553_/Y vssd1 vssd1 vccd1 vccd1 _2554_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_1505_ _3197_/Q _1479_/X _1490_/X _1504_/Y vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__o211a_1
Xoutput169 _2575_/X vssd1 vssd1 vccd1 vccd1 io_dat_o[3] sky130_fd_sc_hd__clkbuf_2
X_2485_ _3114_/Q vssd1 vssd1 vccd1 vccd1 _2485_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1436_ _1599_/A vssd1 vssd1 vccd1 vccd1 _1488_/A sky130_fd_sc_hd__inv_2
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3106_ _3122_/CLK _3106_/D vssd1 vssd1 vccd1 vccd1 _3106_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3037_ _3166_/CLK _3037_/D vssd1 vssd1 vccd1 vccd1 _3037_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput16 io_dat_i[6] vssd1 vssd1 vccd1 vccd1 _1447_/A sky130_fd_sc_hd__buf_1
Xinput27 io_eo[16] vssd1 vssd1 vccd1 vccd1 _2676_/A sky130_fd_sc_hd__clkbuf_2
Xinput38 io_eo[26] vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__clkbuf_2
Xinput49 io_eo[36] vssd1 vssd1 vccd1 vccd1 _2696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2270_ _2478_/B _2868_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _2270_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1985_ _3003_/X _2963_/X vssd1 vssd1 vccd1 vccd1 _2530_/A sky130_fd_sc_hd__and2_1
X_2606_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2606_/Y sky130_fd_sc_hd__inv_2
X_2537_ _2537_/A vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__inv_2
X_2468_ _3174_/Q vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2399_ _2929_/X vssd1 vssd1 vccd1 vccd1 _2399_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1770_ _1768_/Y _1769_/X _1763_/A vssd1 vssd1 vccd1 vccd1 _1770_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2322_ _3033_/Q vssd1 vssd1 vccd1 vccd1 _2322_/Y sky130_fd_sc_hd__inv_2
X_2253_ _2200_/X _2253_/B _2253_/C vssd1 vssd1 vccd1 vccd1 _2253_/Y sky130_fd_sc_hd__nand3b_1
X_2184_ _3030_/Q _2987_/X _2184_/S vssd1 vssd1 vccd1 vccd1 _3030_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1968_ _1968_/A _1968_/B vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__nor2_2
X_1899_ _2743_/X _2940_/X vssd1 vssd1 vccd1 vccd1 _1900_/B sky130_fd_sc_hd__and2_1
XFILLER_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _2386_/Y _2939_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _2940_/X sky130_fd_sc_hd__mux2_2
X_2871_ _2475_/Y _2870_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2871_/X sky130_fd_sc_hd__mux2_1
X_1822_ _2759_/X _2913_/X vssd1 vssd1 vccd1 vccd1 _1855_/A sky130_fd_sc_hd__xor2_4
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1753_ _1753_/A _1753_/B vssd1 vssd1 vccd1 vccd1 _1769_/B sky130_fd_sc_hd__nor2_4
X_1684_ _2793_/X vssd1 vssd1 vccd1 vccd1 _2484_/B sky130_fd_sc_hd__clkbuf_2
X_2305_ _3123_/Q vssd1 vssd1 vccd1 vccd1 _2305_/Y sky130_fd_sc_hd__inv_2
X_2236_ _3020_/Q vssd1 vssd1 vccd1 vccd1 _2236_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2167_ _2725_/X vssd1 vssd1 vccd1 vccd1 _2192_/S sky130_fd_sc_hd__clkbuf_2
X_2098_ _2095_/X _2096_/Y _1672_/X _2097_/Y vssd1 vssd1 vccd1 vccd1 _3055_/D sky130_fd_sc_hd__o2bb2ai_1
XFILLER_21_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _3209_/CLK _3070_/D vssd1 vssd1 vccd1 vccd1 _3070_/Q sky130_fd_sc_hd__dfxtp_1
X_2021_ _2825_/X _1960_/Y _2019_/Y _2017_/A vssd1 vssd1 vccd1 vccd1 _2021_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2923_ _2923_/A0 _3126_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2923_/X sky130_fd_sc_hd__mux2_1
X_2854_ input94/X _3015_/Q _3156_/Q vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__mux2_1
X_1805_ _3111_/Q _2787_/X _1805_/S vssd1 vssd1 vccd1 vccd1 _3111_/D sky130_fd_sc_hd__mux2_1
X_2785_ _2334_/Y _2784_/X _3189_/Q vssd1 vssd1 vccd1 vccd1 _2785_/X sky130_fd_sc_hd__mux2_4
X_1736_ _1730_/X _1734_/Y _1735_/Y vssd1 vssd1 vccd1 vccd1 _1785_/B sky130_fd_sc_hd__o21bai_2
X_1667_ _1667_/A _1666_/X vssd1 vssd1 vccd1 vccd1 _3143_/D sky130_fd_sc_hd__nor2b_1
X_1598_ _3167_/Q vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3199_ _3201_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2219_ _2849_/X _3005_/X vssd1 vssd1 vccd1 vccd1 _2224_/B sky130_fd_sc_hd__or2b_2
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput307 _2722_/X vssd1 vssd1 vccd1 vccd1 io_wo[62] sky130_fd_sc_hd__clkbuf_2
X_2570_ _2495_/Y _2542_/Y _2566_/Y _2568_/Y _2569_/Y vssd1 vssd1 vccd1 vccd1 _2570_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_1521_ _3192_/Q _1506_/X _1510_/X _1520_/Y vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__o211a_1
X_1452_ _3207_/Q _1435_/X _1438_/X _1451_/Y vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__o211a_1
X_3122_ _3122_/CLK _3122_/D vssd1 vssd1 vccd1 vccd1 _3122_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3053_ _3092_/CLK _3053_/D vssd1 vssd1 vccd1 vccd1 _3053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _2017_/A _3075_/Q vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__and2b_1
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2906_ _2432_/Y _2364_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2906_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2837_ _2512_/Y _2836_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__mux2_1
X_2768_ _2261_/Y _2326_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2768_/X sky130_fd_sc_hd__mux2_1
X_1719_ _3007_/X vssd1 vssd1 vccd1 vccd1 _2504_/A sky130_fd_sc_hd__inv_2
X_2699_ _2699_/A vssd1 vssd1 vccd1 vccd1 _2699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2622_ _2611_/X _3183_/Q _2630_/C vssd1 vssd1 vccd1 vccd1 _2622_/Y sky130_fd_sc_hd__nand3b_2
X_2553_ _2600_/A _2600_/B _3154_/Q vssd1 vssd1 vccd1 vccd1 _2553_/Y sky130_fd_sc_hd__nand3_2
X_1504_ _1501_/X _1516_/B _1639_/B vssd1 vssd1 vccd1 vccd1 _1504_/Y sky130_fd_sc_hd__nand3b_1
X_2484_ _2484_/A _2484_/B vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__nand2_1
X_1435_ _2658_/A vssd1 vssd1 vccd1 vccd1 _1435_/X sky130_fd_sc_hd__clkbuf_2
X_3105_ _3122_/CLK _3105_/D vssd1 vssd1 vccd1 vccd1 _3105_/Q sky130_fd_sc_hd__dfxtp_2
X_3036_ _3075_/CLK _3036_/D vssd1 vssd1 vccd1 vccd1 _3036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput17 io_dat_i[7] vssd1 vssd1 vccd1 vccd1 _1443_/A sky130_fd_sc_hd__buf_1
Xinput28 io_eo[17] vssd1 vssd1 vccd1 vccd1 _2677_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput39 io_eo[27] vssd1 vssd1 vccd1 vccd1 _2687_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1984_ _3003_/X _2963_/X vssd1 vssd1 vccd1 vccd1 _1986_/A sky130_fd_sc_hd__nor2_4
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2605_ _2611_/A _3179_/Q _2605_/C vssd1 vssd1 vccd1 vccd1 _2606_/A sky130_fd_sc_hd__nand3b_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_2536_ _2536_/A vssd1 vssd1 vccd1 vccd1 _2536_/Y sky130_fd_sc_hd__inv_2
X_2467_ _3095_/Q vssd1 vssd1 vccd1 vccd1 _2467_/Y sky130_fd_sc_hd__inv_2
X_2398_ _3065_/Q vssd1 vssd1 vccd1 vccd1 _2398_/Y sky130_fd_sc_hd__inv_2
X_3019_ _3205_/CLK _3019_/D vssd1 vssd1 vccd1 vccd1 _3019_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2321_ _3057_/Q vssd1 vssd1 vccd1 vccd1 _2321_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2252_ _2251_/X _3017_/Q _2252_/S vssd1 vssd1 vccd1 vccd1 _3017_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _3031_/Q _2988_/X _2183_/S vssd1 vssd1 vccd1 vccd1 _3031_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1967_ _2999_/X _2955_/X vssd1 vssd1 vccd1 vccd1 _1968_/B sky130_fd_sc_hd__and2_1
X_1898_ _2743_/X _2940_/X vssd1 vssd1 vccd1 vccd1 _1905_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2519_ _2851_/X _3004_/X vssd1 vssd1 vccd1 vccd1 _2519_/X sky130_fd_sc_hd__and2b_1
XFILLER_75_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _2476_/Y _2340_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1821_ _1861_/B _1861_/A _1859_/A _1820_/Y vssd1 vssd1 vccd1 vccd1 _1855_/B sky130_fd_sc_hd__a31o_2
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1752_ _2779_/X _2892_/X _2777_/X _2889_/X vssd1 vssd1 vccd1 vccd1 _1753_/B sky130_fd_sc_hd__a211oi_4
X_1683_ _2791_/X _2859_/X vssd1 vssd1 vccd1 vccd1 _1699_/A sky130_fd_sc_hd__xor2_4
X_2304_ _3091_/Q vssd1 vssd1 vccd1 vccd1 _2304_/Y sky130_fd_sc_hd__inv_2
X_2235_ _2233_/Y _1666_/X _2234_/Y vssd1 vssd1 vccd1 vccd1 _3021_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2166_ _2119_/Y _2114_/X _2118_/Y vssd1 vssd1 vccd1 vccd1 _2166_/X sky130_fd_sc_hd__o21a_1
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2097_ _3055_/Q vssd1 vssd1 vccd1 vccd1 _2097_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2999_ _2358_/Y _2311_/Y _2359_/Y _2360_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _2999_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2020_ _1960_/Y _2019_/Y _2825_/X vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ _2411_/Y _2921_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2922_/X sky130_fd_sc_hd__mux2_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2853_ _2493_/Y _2852_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _2853_/X sky130_fd_sc_hd__mux2_2
X_2784_ _2803_/X _3143_/Q _3188_/Q vssd1 vssd1 vccd1 vccd1 _2784_/X sky130_fd_sc_hd__mux2_1
X_1804_ _3112_/Q _2789_/X _1805_/S vssd1 vssd1 vccd1 vccd1 _3112_/D sky130_fd_sc_hd__mux2_1
X_1735_ _2771_/X _2880_/X vssd1 vssd1 vccd1 vccd1 _1735_/Y sky130_fd_sc_hd__nor2_1
X_1666_ _1728_/S vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__clkbuf_2
X_1597_ _1587_/X _1595_/Y _1673_/A _1596_/Y vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__a211oi_1
X_3198_ _3201_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_2
X_2218_ _3004_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _2220_/B sky130_fd_sc_hd__xnor2_1
X_2149_ _2113_/Y _2149_/B _2149_/C vssd1 vssd1 vccd1 vccd1 _2149_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_41_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput308 _2723_/X vssd1 vssd1 vccd1 vccd1 io_wo[63] sky130_fd_sc_hd__clkbuf_2
X_1520_ _1518_/X _1530_/B _1621_/B vssd1 vssd1 vccd1 vccd1 _1520_/Y sky130_fd_sc_hd__nand3b_1
X_1451_ _1451_/A _1624_/B vssd1 vssd1 vccd1 vccd1 _1451_/Y sky130_fd_sc_hd__nand2_1
X_3121_ _3122_/CLK _3121_/D vssd1 vssd1 vccd1 vccd1 _3121_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _3092_/CLK _3052_/D vssd1 vssd1 vccd1 vccd1 _3052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _2010_/B _2010_/A _2008_/A _1998_/B _1970_/Y vssd1 vssd1 vccd1 vccd1 _2003_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_23_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2905_ _2905_/A0 _3120_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2836_ _2513_/Y _2261_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__mux2_1
X_2767_ _2342_/Y _2766_/X _3191_/Q vssd1 vssd1 vccd1 vccd1 _2767_/X sky130_fd_sc_hd__mux2_4
X_1718_ _3132_/Q _2502_/A _1724_/S vssd1 vssd1 vccd1 vccd1 _3132_/D sky130_fd_sc_hd__mux2_1
X_2698_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__clkbuf_1
X_1649_ _2327_/A _1642_/X _1635_/X _1648_/Y vssd1 vssd1 vccd1 vccd1 _3150_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3139_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2621_ _1602_/Y _2608_/X _2618_/Y _2619_/Y _2620_/Y vssd1 vssd1 vccd1 vccd1 _2621_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2552_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2600_/B sky130_fd_sc_hd__buf_2
X_1503_ input6/X vssd1 vssd1 vccd1 vccd1 _1639_/B sky130_fd_sc_hd__inv_2
X_2483_ _2863_/X vssd1 vssd1 vccd1 vccd1 _2483_/Y sky130_fd_sc_hd__inv_2
X_1434_ _1638_/A vssd1 vssd1 vccd1 vccd1 _2658_/A sky130_fd_sc_hd__buf_1
X_3104_ _3122_/CLK _3104_/D vssd1 vssd1 vccd1 vccd1 _3104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _3075_/CLK _3035_/D vssd1 vssd1 vccd1 vccd1 _3035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ _2637_/Y _2818_/X _3185_/Q vssd1 vssd1 vccd1 vccd1 _2819_/X sky130_fd_sc_hd__mux2_2
XFILLER_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 io_dat_i[8] vssd1 vssd1 vccd1 vccd1 _1440_/A sky130_fd_sc_hd__buf_1
Xinput29 io_eo[18] vssd1 vssd1 vccd1 vccd1 _2678_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1983_ _1993_/B vssd1 vssd1 vccd1 vccd1 _1983_/Y sky130_fd_sc_hd__inv_2
X_2604_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2604_/Y sky130_fd_sc_hd__inv_2
X_2535_ _2535_/A vssd1 vssd1 vccd1 vccd1 _2535_/Y sky130_fd_sc_hd__inv_2
X_2466_ _2466_/A _2769_/X vssd1 vssd1 vccd1 vccd1 _2466_/Y sky130_fd_sc_hd__nand2_1
X_2397_ _2404_/A _2737_/X vssd1 vssd1 vccd1 vccd1 _2397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018_ _3138_/CLK _3018_/D vssd1 vssd1 vccd1 vccd1 _3018_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2320_ _2327_/A _2990_/X vssd1 vssd1 vccd1 vccd1 _2320_/Y sky130_fd_sc_hd__nand2_1
X_2251_ _2251_/A _2251_/B vssd1 vssd1 vccd1 vccd1 _2251_/X sky130_fd_sc_hd__xor2_1
XFILLER_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2182_ _3032_/Q _2989_/X _2183_/S vssd1 vssd1 vccd1 vccd1 _3032_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1966_ _2361_/B _2955_/X vssd1 vssd1 vccd1 vccd1 _1968_/A sky130_fd_sc_hd__nor2_1
X_1897_ _2741_/X _2937_/X vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__xor2_4
X_2518_ _2518_/A vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__inv_2
X_2449_ _3101_/Q vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1820_ _2427_/B _2910_/X _1819_/X vssd1 vssd1 vccd1 vccd1 _1820_/Y sky130_fd_sc_hd__o21ai_1
X_1751_ _1767_/A vssd1 vssd1 vccd1 vccd1 _1754_/B sky130_fd_sc_hd__inv_2
X_1682_ _1676_/X _1680_/Y _1681_/Y vssd1 vssd1 vccd1 vccd1 _1699_/B sky130_fd_sc_hd__o21bai_4
X_2303_ _2303_/A vssd1 vssd1 vccd1 vccd1 _2303_/Y sky130_fd_sc_hd__inv_2
X_2234_ _2244_/B _3021_/Q vssd1 vssd1 vccd1 vccd1 _2234_/Y sky130_fd_sc_hd__nor2_1
X_2165_ _3040_/Q vssd1 vssd1 vccd1 vccd1 _2165_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2096_ _2094_/Y _2035_/Y _2034_/Y _2089_/S vssd1 vssd1 vccd1 vccd1 _2096_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2998_ _2363_/Y _2318_/Y _2364_/Y _2365_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _2998_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3201_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_1949_ _3085_/Q _2763_/X _1952_/S vssd1 vssd1 vccd1 vccd1 _3085_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _2412_/Y _1806_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2921_/X sky130_fd_sc_hd__mux2_1
X_2852_ _2494_/Y _1706_/Y _3204_/Q vssd1 vssd1 vccd1 vccd1 _2852_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1803_ _3113_/Q _2791_/X _1803_/S vssd1 vssd1 vccd1 vccd1 _3113_/D sky130_fd_sc_hd__mux2_1
X_2783_ _2443_/Y _2782_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2783_/X sky130_fd_sc_hd__mux2_2
X_1734_ _1731_/Y _1732_/Y _1791_/A vssd1 vssd1 vccd1 vccd1 _1734_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1665_ _2803_/X vssd1 vssd1 vccd1 vccd1 _1728_/S sky130_fd_sc_hd__clkbuf_2
X_1596_ input9/X _1606_/B _1603_/C vssd1 vssd1 vccd1 vccd1 _1596_/Y sky130_fd_sc_hd__nor3_2
X_2217_ _2217_/A _2225_/C _2217_/C vssd1 vssd1 vccd1 vccd1 _2220_/A sky130_fd_sc_hd__nand3_1
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3197_ _3197_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _2113_/Y _2146_/Y _2149_/C vssd1 vssd1 vccd1 vccd1 _2148_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _2727_/X vssd1 vssd1 vccd1 vccd1 _2177_/S sky130_fd_sc_hd__buf_2
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput309 _2666_/X vssd1 vssd1 vccd1 vccd1 io_wo[6] sky130_fd_sc_hd__clkbuf_2
X_1450_ _1450_/A vssd1 vssd1 vccd1 vccd1 _1624_/B sky130_fd_sc_hd__inv_2
X_3120_ _3123_/CLK _3120_/D vssd1 vssd1 vccd1 vccd1 _3120_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3092_/CLK _3051_/D vssd1 vssd1 vccd1 vccd1 _3051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _2011_/S _2000_/X _2001_/X vssd1 vssd1 vccd1 vccd1 _3076_/D sky130_fd_sc_hd__o21bai_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2904_ _2435_/Y _2903_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__mux2_1
X_2835_ _2514_/Y _2834_/X _3171_/Q vssd1 vssd1 vccd1 vccd1 _2835_/X sky130_fd_sc_hd__mux2_2
X_2766_ _2785_/X _3144_/Q _3190_/Q vssd1 vssd1 vccd1 vccd1 _2766_/X sky130_fd_sc_hd__mux2_1
X_1717_ _3006_/X vssd1 vssd1 vccd1 vccd1 _2502_/A sky130_fd_sc_hd__inv_2
X_2697_ _2697_/A vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__clkbuf_1
X_1648_ _1650_/A _1648_/B vssd1 vssd1 vccd1 vccd1 _1648_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1579_ _1590_/A _1584_/B _1631_/B vssd1 vssd1 vccd1 vccd1 _1579_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _2611_/X _3182_/Q _2620_/C vssd1 vssd1 vccd1 vccd1 _2620_/Y sky130_fd_sc_hd__nand3b_2
X_2551_ _2551_/A vssd1 vssd1 vccd1 vccd1 _2600_/A sky130_fd_sc_hd__buf_2
X_2482_ _3115_/Q vssd1 vssd1 vccd1 vccd1 _2482_/Y sky130_fd_sc_hd__inv_2
X_1502_ _1535_/B vssd1 vssd1 vccd1 vccd1 _1516_/B sky130_fd_sc_hd__buf_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1433_ _1433_/A _1500_/A vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__nor2_2
X_3103_ _3122_/CLK _3103_/D vssd1 vssd1 vccd1 vccd1 _3103_/Q sky130_fd_sc_hd__dfxtp_1
X_3034_ _3201_/CLK _3034_/D vssd1 vssd1 vccd1 vccd1 _3034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ _2515_/Y _2534_/A _3184_/Q vssd1 vssd1 vccd1 vccd1 _2818_/X sky130_fd_sc_hd__mux2_1
X_2749_ _2341_/Y _2748_/X _3193_/Q vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__mux2_4
Xinput19 io_dat_i[9] vssd1 vssd1 vccd1 vccd1 _1511_/A sky130_fd_sc_hd__buf_1
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1982_ _3002_/X _2961_/X vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__and2_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2603_ _3211_/Q _2603_/B _2603_/C vssd1 vssd1 vccd1 vccd1 _2604_/A sky130_fd_sc_hd__nand3_1
X_2534_ _2534_/A vssd1 vssd1 vccd1 vccd1 _2534_/Y sky130_fd_sc_hd__inv_2
X_2465_ _2878_/X vssd1 vssd1 vccd1 vccd1 _2465_/Y sky130_fd_sc_hd__inv_2
X_2396_ _3017_/Q vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3017_ _3138_/CLK _3017_/D vssd1 vssd1 vccd1 vccd1 _3017_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2250_ _2249_/X _3018_/Q _2252_/S vssd1 vssd1 vccd1 vccd1 _3018_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ _3033_/Q _2990_/X _2183_/S vssd1 vssd1 vccd1 vccd1 _3033_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1965_ _2999_/X vssd1 vssd1 vccd1 vccd1 _2361_/B sky130_fd_sc_hd__buf_1
X_1896_ _1936_/B _1936_/A _1934_/A _1895_/Y vssd1 vssd1 vccd1 vccd1 _1930_/B sky130_fd_sc_hd__a31o_2
X_2517_ _3004_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _2518_/A sky130_fd_sc_hd__and2b_1
X_2448_ _2457_/A _2781_/X vssd1 vssd1 vccd1 vccd1 _2448_/Y sky130_fd_sc_hd__nand2_1
X_2379_ _2393_/A _2747_/X vssd1 vssd1 vccd1 vccd1 _2379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1750_ _2781_/X _2895_/X vssd1 vssd1 vccd1 vccd1 _1767_/A sky130_fd_sc_hd__nor2_1
X_1681_ _2789_/X _2856_/X vssd1 vssd1 vccd1 vccd1 _1681_/Y sky130_fd_sc_hd__nor2_2
X_2302_ _3075_/Q vssd1 vssd1 vccd1 vccd1 _2302_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2233_ _2233_/A _2233_/B vssd1 vssd1 vccd1 vccd1 _2233_/Y sky130_fd_sc_hd__xnor2_1
X_2164_ _2163_/Y _3041_/Q _2164_/S vssd1 vssd1 vccd1 vccd1 _3041_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2095_ _2094_/Y _2034_/Y _2035_/Y vssd1 vssd1 vccd1 vccd1 _2095_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2997_ _2368_/Y _1938_/Y _1863_/Y _1701_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _2997_/X sky130_fd_sc_hd__mux4_2
X_1948_ _3086_/Q _2765_/X _1952_/S vssd1 vssd1 vccd1 vccd1 _3086_/D sky130_fd_sc_hd__mux2_1
X_1879_ _3096_/Q _2771_/X _1880_/S vssd1 vssd1 vccd1 vccd1 _3096_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ _2920_/A0 _3125_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2920_/X sky130_fd_sc_hd__mux2_1
X_2851_ _2498_/Y _2850_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__mux2_1
X_1802_ _3114_/Q _2484_/B _1803_/S vssd1 vssd1 vccd1 vccd1 _3114_/D sky130_fd_sc_hd__mux2_1
X_2782_ _2377_/Y _2291_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__mux2_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1733_ _2769_/X _2877_/X vssd1 vssd1 vccd1 vccd1 _1791_/A sky130_fd_sc_hd__nor2_4
X_1664_ _1667_/A _1796_/S vssd1 vssd1 vccd1 vccd1 _3144_/D sky130_fd_sc_hd__nor2b_1
X_1595_ _3168_/Q vssd1 vssd1 vccd1 vccd1 _1595_/Y sky130_fd_sc_hd__inv_2
X_2216_ _2216_/A vssd1 vssd1 vccd1 vccd1 _2217_/C sky130_fd_sc_hd__inv_2
X_3196_ _3197_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2147_/A _2147_/B vssd1 vssd1 vccd1 vccd1 _2149_/C sky130_fd_sc_hd__nor2_1
XFILLER_53_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2078_ _2078_/A _2078_/B vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3074_/CLK _3050_/D vssd1 vssd1 vccd1 vccd1 _3050_/Q sky130_fd_sc_hd__dfxtp_1
X_2001_ _2017_/A _3076_/Q vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2903_ _2436_/Y _1863_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__mux2_1
X_2834_ _2516_/Y _2515_/Y _3170_/Q vssd1 vssd1 vccd1 vccd1 _2834_/X sky130_fd_sc_hd__mux2_1
X_2765_ _2408_/Y _2764_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__mux2_4
X_1716_ _3133_/Q _2500_/A _1724_/S vssd1 vssd1 vccd1 vccd1 _3133_/D sky130_fd_sc_hd__mux2_1
X_2696_ _2696_/A vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__clkbuf_1
X_1647_ _3150_/Q vssd1 vssd1 vccd1 vccd1 _2327_/A sky130_fd_sc_hd__clkbuf_2
X_1578_ _3173_/Q _1570_/X _1571_/X _1577_/Y vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3179_ _3197_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ _2550_/A _2630_/C _2626_/C vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__nand3_2
X_1501_ _1551_/A vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__buf_1
X_2481_ _2484_/A _2795_/X vssd1 vssd1 vccd1 vccd1 _2481_/Y sky130_fd_sc_hd__nand2_1
X_1432_ _1432_/A input3/X vssd1 vssd1 vccd1 vccd1 _1500_/A sky130_fd_sc_hd__nand2_4
X_3102_ _3205_/CLK _3102_/D vssd1 vssd1 vccd1 vccd1 _3102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3033_ _3201_/CLK _3033_/D vssd1 vssd1 vccd1 vccd1 _3033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2817_ _2638_/Y _2816_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2748_ _2767_/X _3145_/Q _3192_/Q vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__mux2_1
X_2679_ _2679_/A vssd1 vssd1 vccd1 vccd1 _2679_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1981_ _1995_/A _1981_/B _1995_/B vssd1 vssd1 vccd1 vccd1 _1981_/Y sky130_fd_sc_hd__nand3_4
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2602_ _2620_/C _2632_/C _3163_/Q vssd1 vssd1 vccd1 vccd1 _2602_/Y sky130_fd_sc_hd__nor3b_2
X_2533_ _2057_/Y _2532_/Y _2059_/Y _2062_/A vssd1 vssd1 vccd1 vccd1 _2534_/A sky130_fd_sc_hd__a31oi_4
X_2464_ _3096_/Q vssd1 vssd1 vccd1 vccd1 _2464_/Y sky130_fd_sc_hd__inv_2
X_2395_ _2932_/X vssd1 vssd1 vccd1 vccd1 _2395_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ _3139_/CLK _3016_/D vssd1 vssd1 vccd1 vccd1 _3016_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2180_ _3034_/Q _2313_/B _2183_/S vssd1 vssd1 vccd1 vccd1 _3034_/D sky130_fd_sc_hd__mux2_1
XFILLER_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1964_ _2998_/X _2953_/X vssd1 vssd1 vccd1 vccd1 _2010_/A sky130_fd_sc_hd__xor2_4
X_1895_ _2393_/B _2934_/X _1894_/X vssd1 vssd1 vccd1 vccd1 _1895_/Y sky130_fd_sc_hd__o21ai_1
X_2516_ _2516_/A vssd1 vssd1 vccd1 vccd1 _2516_/Y sky130_fd_sc_hd__inv_2
X_2447_ _2896_/X vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__inv_2
X_2378_ _2404_/A vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput290 _2707_/X vssd1 vssd1 vccd1 vccd1 io_wo[47] sky130_fd_sc_hd__clkbuf_2
XFILLER_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1680_ _1707_/A _1678_/Y _1679_/Y vssd1 vssd1 vccd1 vccd1 _1680_/Y sky130_fd_sc_hd__a21oi_4
X_2301_ _3036_/Q vssd1 vssd1 vccd1 vccd1 _2301_/Y sky130_fd_sc_hd__inv_2
X_2232_ _2232_/A _2232_/B vssd1 vssd1 vccd1 vccd1 _2233_/B sky130_fd_sc_hd__nand2_1
X_2163_ _2163_/A _2163_/B vssd1 vssd1 vccd1 vccd1 _2163_/Y sky130_fd_sc_hd__xnor2_1
X_2094_ _2094_/A vssd1 vssd1 vccd1 vccd1 _2094_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _2371_/Y _1942_/Y _1870_/Y _1706_/Y _3164_/Q _3165_/Q vssd1 vssd1 vccd1 vccd1
+ _2996_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1947_ _2749_/X vssd1 vssd1 vccd1 vccd1 _1952_/S sky130_fd_sc_hd__clkbuf_2
X_1878_ _3097_/Q _2773_/X _1880_/S vssd1 vssd1 vccd1 vccd1 _3097_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _2499_/Y _2377_/Y _3202_/Q vssd1 vssd1 vccd1 vccd1 _2850_/X sky130_fd_sc_hd__mux2_1
X_1801_ _3115_/Q _2795_/X _1803_/S vssd1 vssd1 vccd1 vccd1 _3115_/D sky130_fd_sc_hd__mux2_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _2447_/Y _2780_/X _3159_/Q vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__mux2_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _2831_/X vssd1 vssd1 vccd1 vccd1 _1732_/Y sky130_fd_sc_hd__inv_2
X_1663_ _2785_/X vssd1 vssd1 vccd1 vccd1 _1796_/S sky130_fd_sc_hd__buf_2
X_1594_ _1587_/X _1588_/Y _1673_/A _1593_/Y vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__a211oi_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2215_ _3006_/X _2847_/X vssd1 vssd1 vccd1 vccd1 _2216_/A sky130_fd_sc_hd__and2b_1
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3195_ _3197_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2146_ _2149_/B vssd1 vssd1 vccd1 vccd1 _2146_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2077_ _2082_/B _2082_/A _2076_/Y vssd1 vssd1 vccd1 vccd1 _2078_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2979_ _2293_/Y _2978_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__mux2_2
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2000_ _2000_/A _2000_/B vssd1 vssd1 vccd1 vccd1 _2000_/X sky130_fd_sc_hd__xor2_1
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _2902_/A0 _3119_/Q _3160_/Q vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2833_ _2495_/Y _2832_/X _3173_/Q vssd1 vssd1 vccd1 vccd1 _2833_/X sky130_fd_sc_hd__mux2_4
X_2764_ _2263_/Y _2409_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__mux2_1
X_1715_ _1728_/S vssd1 vssd1 vccd1 vccd1 _1724_/S sky130_fd_sc_hd__buf_2
X_2695_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1646_ _3151_/Q _1642_/X _1635_/X _1645_/Y vssd1 vssd1 vccd1 vccd1 _3151_/D sky130_fd_sc_hd__o211a_1
X_1577_ _1565_/X _1584_/B _1629_/B vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3178_ _3211_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
X_2129_ _2983_/X _2813_/X _2123_/A _2128_/Y vssd1 vssd1 vccd1 vccd1 _2129_/Y sky130_fd_sc_hd__a2bb2oi_1
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2480_ _2866_/X vssd1 vssd1 vccd1 vccd1 _2480_/Y sky130_fd_sc_hd__inv_2
X_1500_ _1500_/A vssd1 vssd1 vccd1 vccd1 _1551_/A sky130_fd_sc_hd__buf_2
X_1431_ input1/X input2/X vssd1 vssd1 vccd1 vccd1 _1433_/A sky130_fd_sc_hd__nand2_1
X_3101_ _3205_/CLK _3101_/D vssd1 vssd1 vccd1 vccd1 _3101_/Q sky130_fd_sc_hd__dfxtp_1
X_3032_ _3166_/CLK _3032_/D vssd1 vssd1 vccd1 vccd1 _3032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2816_ _2639_/Y _2165_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2816_/X sky130_fd_sc_hd__mux2_1
X_2747_ _2376_/Y _2746_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__mux2_2
X_2678_ _2678_/A vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__clkbuf_1
X_1629_ _1636_/A _1629_/B vssd1 vssd1 vccd1 vccd1 _1629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1980_ _1980_/A _1980_/B vssd1 vssd1 vccd1 vccd1 _1995_/B sky130_fd_sc_hd__nor2_4
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2601_ _2406_/Y _2542_/Y _2597_/Y _2599_/Y _2600_/Y vssd1 vssd1 vccd1 vccd1 _2601_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2532_ _2532_/A vssd1 vssd1 vccd1 vccd1 _2532_/Y sky130_fd_sc_hd__inv_2
X_2463_ _2466_/A _2771_/X vssd1 vssd1 vccd1 vccd1 _2463_/Y sky130_fd_sc_hd__nand2_1
X_2394_ _3066_/Q vssd1 vssd1 vccd1 vccd1 _2394_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3015_ _3139_/CLK _3015_/D vssd1 vssd1 vccd1 vccd1 _3015_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3122_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1963_ _1957_/X _1961_/Y _1962_/Y vssd1 vssd1 vccd1 vccd1 _2010_/B sky130_fd_sc_hd__o21bai_2
X_1894_ _2393_/B _2934_/X _2737_/X _2931_/X vssd1 vssd1 vccd1 vccd1 _1894_/X sky130_fd_sc_hd__a211o_1
X_2515_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__inv_2
X_2446_ _3102_/Q vssd1 vssd1 vccd1 vccd1 _2446_/Y sky130_fd_sc_hd__inv_2
X_2377_ _3022_/Q vssd1 vssd1 vccd1 vccd1 _2377_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput280 _2698_/X vssd1 vssd1 vccd1 vccd1 io_wo[38] sky130_fd_sc_hd__clkbuf_2
Xoutput291 _2708_/X vssd1 vssd1 vccd1 vccd1 io_wo[48] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2300_ _2313_/A _2993_/X vssd1 vssd1 vccd1 vccd1 _2300_/Y sky130_fd_sc_hd__nand2_1
X_2231_ _3005_/X _2849_/X vssd1 vssd1 vccd1 vccd1 _2233_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2162_ _2161_/X _3042_/Q _2164_/S vssd1 vssd1 vccd1 vccd1 _3042_/D sky130_fd_sc_hd__mux2_1
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2093_ _2177_/S _2090_/Y _2091_/X _2092_/Y vssd1 vssd1 vccd1 vccd1 _3056_/D sky130_fd_sc_hd__o22ai_4
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2995_ _2291_/Y _1956_/Y _1881_/Y _1729_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2995_/X sky130_fd_sc_hd__mux4_2
X_1946_ _2025_/S _1942_/Y _1944_/X _1945_/Y vssd1 vssd1 vccd1 vccd1 _3087_/D sky130_fd_sc_hd__o22ai_1
X_1877_ _3098_/Q _2457_/B _1880_/S vssd1 vssd1 vccd1 vccd1 _3098_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2429_ _2908_/X vssd1 vssd1 vccd1 vccd1 _2429_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1800_ _3116_/Q _2478_/B _1803_/S vssd1 vssd1 vccd1 vccd1 _3116_/D sky130_fd_sc_hd__mux2_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _2382_/Y _2295_/Y _3158_/Q vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__mux2_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ _2769_/X _2877_/X vssd1 vssd1 vccd1 vccd1 _1731_/Y sky130_fd_sc_hd__nand2_2
X_1662_ _1667_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _3145_/D sky130_fd_sc_hd__nor2b_1
X_1593_ _1593_/A _1606_/B _1603_/C vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__nor3_2
X_3194_ _3197_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_2
X_2214_ _2214_/A vssd1 vssd1 vccd1 vccd1 _2225_/C sky130_fd_sc_hd__inv_2
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2145_ _3045_/Q vssd1 vssd1 vccd1 vccd1 _2145_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _2992_/X _2973_/X vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2978_ _2294_/Y _2032_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__mux2_1
X_1929_ _1670_/X _1923_/Y _1928_/Y vssd1 vssd1 vccd1 vccd1 _3092_/D sky130_fd_sc_hd__o21ai_1
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3197_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2901_ _2439_/Y _2900_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2832_ _2496_/Y _2540_/A _3172_/Q vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2763_ _2413_/Y _2762_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__mux2_2
X_1714_ _3005_/X vssd1 vssd1 vccd1 vccd1 _2500_/A sky130_fd_sc_hd__inv_2
X_2694_ _2694_/A vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1645_ _1650_/A _1645_/B vssd1 vssd1 vccd1 vccd1 _1645_/Y sky130_fd_sc_hd__nand2_1
X_1576_ _3174_/Q _1570_/X _1571_/X _1575_/Y vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__o211a_1
X_3177_ _3193_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2128_ _2983_/X _2813_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _2128_/Y sky130_fd_sc_hd__a21oi_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2059_ _2070_/B vssd1 vssd1 vccd1 vccd1 _2059_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1430_ _3210_/Q vssd1 vssd1 vccd1 vccd1 _2404_/A sky130_fd_sc_hd__clkbuf_2
X_3100_ _3205_/CLK _3100_/D vssd1 vssd1 vccd1 vccd1 _3100_/Q sky130_fd_sc_hd__dfxtp_1
X_3031_ _3166_/CLK _3031_/D vssd1 vssd1 vccd1 vccd1 _3031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2815_ _2640_/Y _2814_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2746_ _1729_/Y _2377_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__mux2_1
X_2677_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__clkbuf_1
X_1628_ _3158_/Q _1626_/X _1623_/X _1627_/Y vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__o211a_1
X_1559_ _3180_/Q _1556_/X _1557_/X _1558_/Y vssd1 vssd1 vccd1 vccd1 _3180_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _2600_/A _2600_/B _3162_/Q vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__nand3_2
X_2531_ _1981_/Y _2530_/Y _1983_/Y _1986_/A vssd1 vssd1 vccd1 vccd1 _2535_/A sky130_fd_sc_hd__a31oi_4
X_2462_ _2881_/X vssd1 vssd1 vccd1 vccd1 _2462_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2393_ _2393_/A _2393_/B vssd1 vssd1 vccd1 vccd1 _2393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _3205_/CLK _3014_/D vssd1 vssd1 vccd1 vccd1 _3014_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2729_ _2348_/Y _2728_/X _3197_/Q vssd1 vssd1 vccd1 vccd1 _2729_/X sky130_fd_sc_hd__mux2_4
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1962_ _2997_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _1962_/Y sky130_fd_sc_hd__nor2_1
X_1893_ _1893_/A _1893_/B vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__nor2_1
X_2514_ _3170_/Q vssd1 vssd1 vccd1 vccd1 _2514_/Y sky130_fd_sc_hd__inv_2
X_2445_ _2457_/A _2783_/X vssd1 vssd1 vccd1 vccd1 _2445_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _2947_/X vssd1 vssd1 vccd1 vccd1 _2376_/Y sky130_fd_sc_hd__inv_2
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput270 _2689_/X vssd1 vssd1 vccd1 vccd1 io_wo[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput281 _2699_/X vssd1 vssd1 vccd1 vccd1 io_wo[39] sky130_fd_sc_hd__clkbuf_2
Xoutput292 _2709_/X vssd1 vssd1 vccd1 vccd1 io_wo[49] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2230_ _2230_/A _2230_/B vssd1 vssd1 vccd1 vccd1 _3022_/D sky130_fd_sc_hd__nand2_1
X_2161_ _2161_/A _2161_/B vssd1 vssd1 vccd1 vccd1 _2161_/X sky130_fd_sc_hd__xor2_1
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2092_ _2038_/Y _2033_/X _2037_/Y _2727_/X vssd1 vssd1 vccd1 vccd1 _2092_/Y sky130_fd_sc_hd__o31ai_4
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2994_ _2295_/Y _1992_/Y _1917_/Y _1766_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2994_/X sky130_fd_sc_hd__mux4_2
X_1945_ _2827_/X _1885_/Y _1943_/Y _2026_/A vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__o31ai_1
X_1876_ _3099_/Q _2777_/X _1880_/S vssd1 vssd1 vccd1 vccd1 _3099_/D sky130_fd_sc_hd__mux2_1
XFILLER_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2428_ _3082_/Q vssd1 vssd1 vccd1 vccd1 _2428_/Y sky130_fd_sc_hd__inv_2
X_2359_ _3106_/Q vssd1 vssd1 vccd1 vccd1 _2359_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1730_ _2771_/X _2880_/X vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__and2_1
X_1661_ _2767_/X vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__clkbuf_2
X_1592_ _2608_/A vssd1 vssd1 vccd1 vccd1 _1603_/C sky130_fd_sc_hd__buf_2
X_3193_ _3193_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2213_ _3005_/X _2849_/X vssd1 vssd1 vccd1 vccd1 _2214_/A sky130_fd_sc_hd__and2b_1
X_2144_ _2107_/Y _2184_/S _2143_/Y vssd1 vssd1 vccd1 vccd1 _3046_/D sky130_fd_sc_hd__o21ai_1
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2075_ _3060_/Q vssd1 vssd1 vccd1 vccd1 _2075_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2977_ _2296_/Y _2976_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__mux2_1
X_1928_ _1928_/A _2025_/S vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__nand2_1
X_1859_ _1859_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2900_ _2440_/Y _1870_/Y _3208_/Q vssd1 vssd1 vccd1 vccd1 _2900_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _2468_/Y _2830_/X _3175_/Q vssd1 vssd1 vccd1 vccd1 _2831_/X sky130_fd_sc_hd__mux2_1
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2762_ _2340_/Y _2414_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _3134_/Q _2498_/A _2244_/B vssd1 vssd1 vccd1 vccd1 _3134_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2693_ _2693_/A vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__clkbuf_1
X_1644_ _2372_/A _1642_/X _1635_/X _1643_/Y vssd1 vssd1 vccd1 vccd1 _3152_/D sky130_fd_sc_hd__o211a_1
X_1575_ _1565_/X _1584_/B _1627_/B vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3176_ _3209_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2127_ _2163_/A _2161_/A vssd1 vssd1 vccd1 vccd1 _2127_/Y sky130_fd_sc_hd__nor2_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2994_/X _2977_/X vssd1 vssd1 vccd1 vccd1 _2070_/B sky130_fd_sc_hd__and2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3030_ _3166_/CLK _3030_/D vssd1 vssd1 vccd1 vccd1 _3030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2814_ _2641_/Y _2642_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__mux2_1
X_2745_ _2381_/Y _2744_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__mux2_1
X_2676_ _2676_/A vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__clkbuf_1
X_1627_ _1627_/A _1627_/B vssd1 vssd1 vccd1 vccd1 _1627_/Y sky130_fd_sc_hd__nand2_1
X_1558_ _1551_/X _1558_/B _1643_/B vssd1 vssd1 vccd1 vccd1 _1558_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1489_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__clkbuf_2
X_3159_ _3193_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2530_/A vssd1 vssd1 vccd1 vccd1 _2530_/Y sky130_fd_sc_hd__inv_2
X_2461_ _3097_/Q vssd1 vssd1 vccd1 vccd1 _2461_/Y sky130_fd_sc_hd__inv_2
X_2392_ _3018_/Q vssd1 vssd1 vccd1 vccd1 _2392_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3013_ _3139_/CLK _3013_/D vssd1 vssd1 vccd1 vccd1 _3013_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2728_ _2731_/X _3141_/Q _3196_/Q vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__mux2_1
X_2659_ _3211_/Q _1451_/A _1459_/A _2658_/Y vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1961_ _2019_/A _1959_/Y _1960_/Y vssd1 vssd1 vccd1 vccd1 _1961_/Y sky130_fd_sc_hd__a21oi_4
X_1892_ _2739_/X _2934_/X vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__and2_1
X_2513_ _3127_/Q vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2444_ _2466_/A vssd1 vssd1 vccd1 vccd1 _2457_/A sky130_fd_sc_hd__clkbuf_2
X_2375_ _2375_/A vssd1 vssd1 vccd1 vccd1 _2375_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput260 _2661_/X vssd1 vssd1 vccd1 vccd1 io_wo[1] sky130_fd_sc_hd__clkbuf_2
Xoutput271 _2662_/X vssd1 vssd1 vccd1 vccd1 io_wo[2] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_0 _2295_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput282 _2663_/X vssd1 vssd1 vccd1 vccd1 io_wo[3] sky130_fd_sc_hd__clkbuf_2
Xoutput293 _2664_/X vssd1 vssd1 vccd1 vccd1 io_wo[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2160_ _2163_/B _2125_/B _2125_/A vssd1 vssd1 vccd1 vccd1 _2161_/B sky130_fd_sc_hd__a21boi_1
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2091_ _2038_/Y _2033_/X _2037_/Y vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2299_/Y _2298_/Y _1923_/Y _1772_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2993_/X sky130_fd_sc_hd__mux4_2
X_1944_ _1885_/Y _1943_/Y _2827_/X vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1875_ _2767_/X vssd1 vssd1 vccd1 vccd1 _1880_/S sky130_fd_sc_hd__buf_2
X_2427_ _2427_/A _2427_/B vssd1 vssd1 vccd1 vccd1 _2427_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2358_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2358_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2289_ _2289_/A _2289_/B vssd1 vssd1 vccd1 vccd1 _2289_/X sky130_fd_sc_hd__xor2_1
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _1667_/A _1659_/X vssd1 vssd1 vccd1 vccd1 _3146_/D sky130_fd_sc_hd__nor2b_1
XFILLER_50_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1591_ _2551_/A _2552_/A vssd1 vssd1 vccd1 vccd1 _2608_/A sky130_fd_sc_hd__nand2_2
X_3192_ _3193_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2212_ _2244_/C _2212_/B vssd1 vssd1 vccd1 vccd1 _2217_/A sky130_fd_sc_hd__nand2_1
X_2143_ _2140_/Y _2141_/X _2150_/A vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2074_ _1672_/X _2069_/Y _2073_/Y vssd1 vssd1 vccd1 vccd1 _3061_/D sky130_fd_sc_hd__o21ai_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2976_ _2297_/Y _2069_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__mux2_1
X_1927_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2025_/S sky130_fd_sc_hd__clkbuf_2
X_1858_ _2755_/X _2907_/X _1857_/Y vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1789_ _1735_/Y _1730_/X _1734_/Y _2767_/X vssd1 vssd1 vccd1 vccd1 _1789_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2830_ _2469_/Y _2539_/A _3174_/Q vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__mux2_1
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _2417_/Y _2760_/X _3161_/Q vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__mux2_4
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1712_ _2803_/X vssd1 vssd1 vccd1 vccd1 _2244_/B sky130_fd_sc_hd__buf_2
X_2692_ _2692_/A vssd1 vssd1 vccd1 vccd1 _2692_/X sky130_fd_sc_hd__clkbuf_1
X_1643_ _1650_/A _1643_/B vssd1 vssd1 vccd1 vccd1 _1643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1574_ _2542_/A vssd1 vssd1 vccd1 vccd1 _1584_/B sky130_fd_sc_hd__clkbuf_2
X_3175_ _3209_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
X_2126_ _2983_/X _2813_/X vssd1 vssd1 vccd1 vccd1 _2161_/A sky130_fd_sc_hd__xnor2_2
XFILLER_19_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2072_/A _2057_/B _2072_/B vssd1 vssd1 vccd1 vccd1 _2057_/Y sky130_fd_sc_hd__nand3_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _2350_/Y _2958_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__mux2_2
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2813_ _2643_/Y _2812_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2813_/X sky130_fd_sc_hd__mux2_2
X_2744_ _1766_/Y _2382_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__mux2_1
X_2675_ _2675_/A vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__clkbuf_1
X_1626_ _1626_/A vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__clkbuf_2
X_1557_ _1557_/A vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__clkbuf_2
X_1488_ _1488_/A vssd1 vssd1 vccd1 vccd1 _1635_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3158_ _3189_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_4
X_2109_ _2985_/X _2809_/X vssd1 vssd1 vccd1 vccd1 _2132_/B sky130_fd_sc_hd__and2_1
X_3089_ _3110_/CLK _3089_/D vssd1 vssd1 vccd1 vccd1 _3089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2460_ _2466_/A _2773_/X vssd1 vssd1 vccd1 vccd1 _2460_/Y sky130_fd_sc_hd__nand2_1
X_2391_ _2935_/X vssd1 vssd1 vccd1 vccd1 _2391_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3012_ _3139_/CLK _3012_/D vssd1 vssd1 vccd1 vccd1 _3012_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2727_ _2355_/Y _2726_/X _3199_/Q vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__mux2_4
X_2658_ _2658_/A _2658_/B vssd1 vssd1 vccd1 vccd1 _2658_/Y sky130_fd_sc_hd__nand2_1
X_1609_ input5/X _1609_/B _2608_/A vssd1 vssd1 vccd1 vccd1 _1609_/Y sky130_fd_sc_hd__nor3_1
X_2589_ _2600_/A _2600_/B _3160_/Q vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__nand3_2
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _2996_/X _2949_/X vssd1 vssd1 vccd1 vccd1 _1960_/Y sky130_fd_sc_hd__nor2_4
X_1891_ _2393_/B _2934_/X vssd1 vssd1 vccd1 vccd1 _1893_/A sky130_fd_sc_hd__nor2_1
X_2512_ _2512_/A _2550_/A vssd1 vssd1 vccd1 vccd1 _2512_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2443_ _2899_/X vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__inv_2
X_2374_ _3180_/Q vssd1 vssd1 vccd1 vccd1 _2374_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput250 _2670_/X vssd1 vssd1 vccd1 vccd1 io_wo[10] sky130_fd_sc_hd__clkbuf_2
Xoutput261 _2680_/X vssd1 vssd1 vccd1 vccd1 io_wo[20] sky130_fd_sc_hd__clkbuf_2
Xoutput294 _2710_/X vssd1 vssd1 vccd1 vccd1 io_wo[50] sky130_fd_sc_hd__clkbuf_2
Xoutput272 _2690_/X vssd1 vssd1 vccd1 vccd1 io_wo[30] sky130_fd_sc_hd__clkbuf_2
Xoutput283 _2700_/X vssd1 vssd1 vccd1 vccd1 io_wo[40] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_1 _2662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2090_ _3056_/Q vssd1 vssd1 vccd1 vccd1 _2090_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _3138_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2992_ _2303_/Y _2302_/Y _2304_/Y _2305_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2992_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1943_ _1943_/A vssd1 vssd1 vccd1 vccd1 _1943_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1874_ _3100_/Q _2779_/X _1874_/S vssd1 vssd1 vccd1 vccd1 _3100_/D sky130_fd_sc_hd__mux2_1
X_2426_ _2426_/A vssd1 vssd1 vccd1 vccd1 _2426_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2357_ _3051_/Q vssd1 vssd1 vccd1 vccd1 _2357_/Y sky130_fd_sc_hd__inv_2
X_2288_ _1691_/A _1691_/B _2287_/Y vssd1 vssd1 vccd1 vccd1 _2289_/B sky130_fd_sc_hd__o21bai_1
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1590_/A vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__clkbuf_2
X_3191_ _3193_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
X_2211_ _2237_/A _2211_/B vssd1 vssd1 vccd1 vccd1 _2212_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2142_ _2725_/X vssd1 vssd1 vccd1 vccd1 _2150_/A sky130_fd_sc_hd__inv_2
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2073_ _2071_/Y _2072_/X _2066_/A vssd1 vssd1 vccd1 vccd1 _2073_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2975_ _2300_/Y _2974_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2975_/X sky130_fd_sc_hd__mux2_2
X_1926_ _1926_/A _1926_/B vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__xnor2_1
X_1857_ _1861_/B _1861_/A vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1788_ _1735_/Y _1730_/X _1734_/Y vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__o21a_1
X_2409_ _2409_/A vssd1 vssd1 vccd1 vccd1 _2409_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _2347_/Y _2418_/Y _3160_/Q vssd1 vssd1 vccd1 vccd1 _2760_/X sky130_fd_sc_hd__mux2_1
X_1711_ _3004_/X vssd1 vssd1 vccd1 vccd1 _2498_/A sky130_fd_sc_hd__inv_2
X_2691_ _2691_/A vssd1 vssd1 vccd1 vccd1 _2691_/X sky130_fd_sc_hd__clkbuf_1
X_1642_ _2658_/A vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__buf_1
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1573_ _3175_/Q _1570_/X _1571_/X _1572_/Y vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__o211a_1
XFILLER_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3174_ _3205_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
X_2125_ _2125_/A _2125_/B vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2056_/A _2056_/B vssd1 vssd1 vccd1 vccd1 _2072_/B sky130_fd_sc_hd__nor2_4
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _2351_/Y _2298_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2958_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1909_ _2747_/X _2946_/X vssd1 vssd1 vccd1 vccd1 _1911_/A sky130_fd_sc_hd__nor2_4
X_2889_ _2454_/Y _2888_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__mux2_4
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput150 io_i_7_in1[2] vssd1 vssd1 vccd1 vccd1 _2430_/A sky130_fd_sc_hd__buf_1
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2812_ _2644_/Y _2645_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2812_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2743_ _2385_/Y _2742_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2743_/X sky130_fd_sc_hd__mux2_4
X_2674_ _2674_/A vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__clkbuf_1
X_1625_ _3159_/Q _1613_/X _1623_/X _1624_/Y vssd1 vssd1 vccd1 vccd1 _3159_/D sky130_fd_sc_hd__o211a_1
X_1556_ _1570_/A vssd1 vssd1 vccd1 vccd1 _1556_/X sky130_fd_sc_hd__clkbuf_2
X_1487_ _3201_/Q _1479_/X _1459_/X _1486_/Y vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ _3189_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2108_ _2725_/X vssd1 vssd1 vccd1 vccd1 _2184_/S sky130_fd_sc_hd__clkbuf_2
X_3088_ _3110_/CLK _3088_/D vssd1 vssd1 vccd1 vccd1 _3088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _2033_/X _2037_/Y _2038_/Y vssd1 vssd1 vccd1 vccd1 _2088_/B sky130_fd_sc_hd__o21bai_4
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3166_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _3067_/Q vssd1 vssd1 vccd1 vccd1 _2390_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3011_ input85/X _2438_/A _2326_/A _3011_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3011_/X sky130_fd_sc_hd__mux4_2
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2726_ _2729_/X _3147_/Q _3198_/Q vssd1 vssd1 vccd1 vccd1 _2726_/X sky130_fd_sc_hd__mux2_1
X_2657_ _2987_/X _2805_/X _2656_/Y vssd1 vssd1 vccd1 vccd1 _2657_/Y sky130_fd_sc_hd__a21oi_4
X_1608_ _3164_/Q vssd1 vssd1 vccd1 vccd1 _1608_/Y sky130_fd_sc_hd__inv_2
X_2588_ _3208_/Q _2610_/B _2626_/C vssd1 vssd1 vccd1 vccd1 _2588_/Y sky130_fd_sc_hd__nand3_2
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1539_ _2598_/A _2551_/A _1551_/A vssd1 vssd1 vccd1 vccd1 _1570_/A sky130_fd_sc_hd__nor3_4
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3209_ _3209_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1890_ _2739_/X vssd1 vssd1 vccd1 vccd1 _2393_/B sky130_fd_sc_hd__buf_1
X_2511_ _3128_/Q vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__inv_2
X_2442_ _2442_/A vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2373_ _3047_/Q vssd1 vssd1 vccd1 vccd1 _2373_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2709_/A vssd1 vssd1 vccd1 vccd1 _2709_/X sky130_fd_sc_hd__clkbuf_2
Xoutput240 _3039_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput251 _2671_/X vssd1 vssd1 vccd1 vccd1 io_wo[11] sky130_fd_sc_hd__clkbuf_2
Xoutput262 _2681_/X vssd1 vssd1 vccd1 vccd1 io_wo[21] sky130_fd_sc_hd__clkbuf_2
Xoutput295 _2711_/X vssd1 vssd1 vccd1 vccd1 io_wo[51] sky130_fd_sc_hd__clkbuf_2
XFILLER_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput273 _2691_/X vssd1 vssd1 vccd1 vccd1 io_wo[31] sky130_fd_sc_hd__clkbuf_2
Xoutput284 _2701_/X vssd1 vssd1 vccd1 vccd1 io_wo[41] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_2 _2695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ _2310_/Y _2309_/Y _2311_/Y _2312_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2991_/X sky130_fd_sc_hd__mux4_2
X_1942_ _3087_/Q vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__inv_2
X_1873_ _3101_/Q _2781_/X _1874_/S vssd1 vssd1 vccd1 vccd1 _3101_/D sky130_fd_sc_hd__mux2_1
X_2425_ _2911_/X vssd1 vssd1 vccd1 vccd1 _2425_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2356_ _2361_/A _3000_/X vssd1 vssd1 vccd1 vccd1 _2356_/Y sky130_fd_sc_hd__nand2_1
X_2287_ _2795_/X _2865_/X vssd1 vssd1 vccd1 vccd1 _2287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2210_ _2847_/X _3006_/X vssd1 vssd1 vccd1 vccd1 _2211_/B sky130_fd_sc_hd__and2b_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3190_ _3193_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2141_ _2141_/A _2141_/B _2141_/C vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__and3_1
X_2072_ _2072_/A _2072_/B _2072_/C vssd1 vssd1 vccd1 vccd1 _2072_/X sky130_fd_sc_hd__and3_1
XFILLER_34_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2974_ _2301_/Y _2075_/Y _3150_/Q vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__mux2_1
X_1925_ _1930_/B _1930_/A _1924_/Y vssd1 vssd1 vccd1 vccd1 _1926_/B sky130_fd_sc_hd__a21oi_1
X_1856_ _1855_/X _3107_/Q _1862_/S vssd1 vssd1 vccd1 vccd1 _3107_/D sky130_fd_sc_hd__mux2_1
X_1787_ _3120_/Q vssd1 vssd1 vccd1 vccd1 _1787_/Y sky130_fd_sc_hd__inv_2
X_2408_ _2923_/X vssd1 vssd1 vccd1 vccd1 _2408_/Y sky130_fd_sc_hd__inv_2
X_2339_ _2339_/A vssd1 vssd1 vccd1 vccd1 _2339_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1710_ _1796_/S _1706_/Y _1708_/X _1709_/Y vssd1 vssd1 vccd1 vccd1 _3135_/D sky130_fd_sc_hd__o22ai_1
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2690_/X sky130_fd_sc_hd__clkbuf_1
X_1641_ _3152_/Q vssd1 vssd1 vccd1 vccd1 _2372_/A sky130_fd_sc_hd__buf_2
X_1572_ _1565_/X _1572_/B _1624_/B vssd1 vssd1 vccd1 vccd1 _1572_/Y sky130_fd_sc_hd__nand3b_1
X_3173_ _3189_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
X_2124_ _2982_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _2125_/B sky130_fd_sc_hd__nand2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2993_/X _2975_/X _2992_/X _2973_/X vssd1 vssd1 vccd1 vccd1 _2056_/B sky130_fd_sc_hd__a211oi_4
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _2356_/Y _2956_/X _3153_/Q vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__mux2_4
X_2888_ _2455_/Y _2305_/Y _3206_/Q vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__mux2_1
X_1908_ _1918_/B vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__inv_2
X_1839_ _2749_/X vssd1 vssd1 vccd1 vccd1 _1848_/A sky130_fd_sc_hd__inv_2
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput140 io_i_6_in1[1] vssd1 vssd1 vccd1 vccd1 _2323_/A sky130_fd_sc_hd__buf_1
Xinput151 io_i_7_in1[3] vssd1 vssd1 vccd1 vccd1 _2426_/A sky130_fd_sc_hd__buf_1
XFILLER_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2811_ _2646_/Y _2810_/X _3149_/Q vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__mux2_2
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ _1772_/Y _2236_/Y _3162_/Q vssd1 vssd1 vccd1 vccd1 _2742_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _2673_/A vssd1 vssd1 vccd1 vccd1 _2673_/X sky130_fd_sc_hd__clkbuf_1
X_1624_ _1627_/A _1624_/B vssd1 vssd1 vccd1 vccd1 _1624_/Y sky130_fd_sc_hd__nand2_1
X_1555_ _3181_/Q _1540_/X _1541_/X _1554_/Y vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1486_ _1609_/B _1498_/B _1650_/B vssd1 vssd1 vccd1 vccd1 _1486_/Y sky130_fd_sc_hd__nand3b_1
X_3156_ _3189_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_4
X_3087_ _3092_/CLK _3087_/D vssd1 vssd1 vccd1 vccd1 _3087_/Q sky130_fd_sc_hd__dfxtp_1
X_2107_ _3046_/Q vssd1 vssd1 vccd1 vccd1 _2107_/Y sky130_fd_sc_hd__inv_2
X_2038_ _2989_/X _2967_/X vssd1 vssd1 vccd1 vccd1 _2038_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ input86/X _2434_/A _2323_/A _3010_/A3 _3154_/Q _3155_/Q vssd1 vssd1 vccd1
+ vccd1 _3010_/X sky130_fd_sc_hd__mux4_2
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2725_ _2541_/Y _2724_/X _3201_/Q vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__mux2_8
X_2656_ _2987_/X _2805_/X _2141_/C _2141_/A vssd1 vssd1 vccd1 vccd1 _2656_/Y sky130_fd_sc_hd__a2bb2oi_2
X_1607_ _1587_/X _1605_/Y _1655_/A _1606_/Y vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__a211oi_2
X_2587_ _2593_/B _3192_/Q _2618_/C vssd1 vssd1 vccd1 vccd1 _2587_/Y sky130_fd_sc_hd__nand3b_4
X_1538_ input1/X vssd1 vssd1 vccd1 vccd1 _2551_/A sky130_fd_sc_hd__inv_2
X_1469_ _3203_/Q _1458_/X _1459_/X _1468_/Y vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3208_ _3209_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_4
X_3139_ _3139_/CLK _3139_/D vssd1 vssd1 vccd1 vccd1 _3139_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2510_ _2510_/A _2550_/A vssd1 vssd1 vccd1 vccd1 _2510_/Y sky130_fd_sc_hd__nand2_1
X_2441_ _3176_/Q vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2372_ _2372_/A _2996_/X vssd1 vssd1 vccd1 vccd1 _2372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2708_ _2708_/A vssd1 vssd1 vccd1 vccd1 _2708_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput241 _3040_/Q vssd1 vssd1 vccd1 vccd1 io_o_7_out[1] sky130_fd_sc_hd__clkbuf_2
Xoutput230 _2534_/Y vssd1 vssd1 vccd1 vccd1 io_o_6_co sky130_fd_sc_hd__clkbuf_2
Xoutput252 _2672_/X vssd1 vssd1 vccd1 vccd1 io_wo[12] sky130_fd_sc_hd__clkbuf_2
X_2639_ _3024_/Q vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput263 _2682_/X vssd1 vssd1 vccd1 vccd1 io_wo[22] sky130_fd_sc_hd__clkbuf_2
Xoutput274 _2692_/X vssd1 vssd1 vccd1 vccd1 io_wo[32] sky130_fd_sc_hd__clkbuf_2
Xoutput285 _2702_/X vssd1 vssd1 vccd1 vccd1 io_wo[42] sky130_fd_sc_hd__clkbuf_2
Xoutput296 _2712_/X vssd1 vssd1 vccd1 vccd1 io_wo[52] sky130_fd_sc_hd__clkbuf_2
XINSDIODE2_3 _2664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2990_ _2317_/Y _2316_/Y _2318_/Y _2319_/Y _3166_/Q _3167_/Q vssd1 vssd1 vccd1 vccd1
+ _2990_/X sky130_fd_sc_hd__mux4_2
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1670_/X _1938_/Y _1939_/X _1940_/Y vssd1 vssd1 vccd1 vccd1 _3088_/D sky130_fd_sc_hd__o22ai_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1872_ _3102_/Q _2783_/X _1874_/S vssd1 vssd1 vccd1 vccd1 _3102_/D sky130_fd_sc_hd__mux2_1
X_2424_ _3083_/Q vssd1 vssd1 vccd1 vccd1 _2424_/Y sky130_fd_sc_hd__inv_2
X_2355_ _2541_/A _3198_/Q vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__nand2_1
X_2286_ _2285_/X _3013_/Q _2290_/S vssd1 vssd1 vccd1 vccd1 _3013_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2140_ _2141_/A _2141_/C _2141_/B vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _2072_/A _2072_/B _2072_/C vssd1 vssd1 vccd1 vccd1 _2071_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2973_ _2306_/Y _2972_/X _3151_/Q vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__mux2_4
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _2741_/X _2937_/X vssd1 vssd1 vccd1 vccd1 _1924_/Y sky130_fd_sc_hd__nor2_1
X_1855_ _1855_/A _1855_/B vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__xor2_1
X_1786_ _1785_/X _3121_/Q _1786_/S vssd1 vssd1 vccd1 vccd1 _3121_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2407_ _2407_/A vssd1 vssd1 vccd1 vccd1 _2407_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2338_ _3054_/Q vssd1 vssd1 vccd1 vccd1 _2338_/Y sky130_fd_sc_hd__inv_2
X_2269_ _2478_/B _2868_/X _2795_/X _2865_/X vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__a211o_1
XFILLER_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1640_ _3153_/Q _1458_/X _1635_/X _1639_/Y vssd1 vssd1 vccd1 vccd1 _3153_/D sky130_fd_sc_hd__o211a_1
X_1571_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _3205_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
X_2123_ _2123_/A _2123_/B vssd1 vssd1 vccd1 vccd1 _2125_/A sky130_fd_sc_hd__nand2_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _2070_/A vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__inv_2
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2956_ _2357_/Y _2302_/Y _3152_/Q vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__mux2_1
X_2887_ _2887_/A0 _3138_/Q _3158_/Q vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__mux2_1
X_1907_ _2745_/X _2943_/X vssd1 vssd1 vccd1 vccd1 _1918_/B sky130_fd_sc_hd__and2_1
X_1838_ _2526_/A _1836_/A _1833_/Y _1831_/Y vssd1 vssd1 vccd1 vccd1 _1838_/X sky130_fd_sc_hd__o211a_1
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1769_ _1769_/A _1769_/B _1769_/C vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__and3_1
XFILLER_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput141 io_i_6_in1[2] vssd1 vssd1 vccd1 vccd1 _2317_/A sky130_fd_sc_hd__buf_1
Xinput130 io_i_5_in1[0] vssd1 vssd1 vccd1 vccd1 _2371_/A sky130_fd_sc_hd__clkbuf_1
Xinput152 io_i_7_in1[4] vssd1 vssd1 vccd1 vccd1 _2422_/A sky130_fd_sc_hd__buf_1
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _2647_/Y _2648_/Y _3148_/Q vssd1 vssd1 vccd1 vccd1 _2810_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2741_ _2388_/Y _2740_/X _3163_/Q vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__mux2_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2672_ _2672_/A vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__clkbuf_1
X_1623_ _1635_/A vssd1 vssd1 vccd1 vccd1 _1623_/X sky130_fd_sc_hd__clkbuf_2
X_1554_ _1551_/X _1558_/B _1639_/B vssd1 vssd1 vccd1 vccd1 _1554_/Y sky130_fd_sc_hd__nand3b_1
X_1485_ _1593_/A vssd1 vssd1 vccd1 vccd1 _1650_/B sky130_fd_sc_hd__inv_2
.ends

