magic
tech sky130A
magscale 1 2
timestamp 1624054006
<< locali >>
rect 38945 92531 38979 93245
rect 26801 86683 26835 86921
rect 30849 80155 30883 80393
rect 30941 80087 30975 80325
rect 38945 67643 38979 68221
rect 33425 62135 33459 62305
rect 38945 57307 38979 58361
rect 26249 56695 26283 56865
rect 29285 43707 29319 43945
rect 36185 41055 36219 41225
rect 36185 39967 36219 40069
rect 36185 38879 36219 39049
rect 35725 36703 35759 36873
rect 26157 33847 26191 34153
rect 24777 31671 24811 31909
rect 35909 30107 35943 30345
rect 16037 19159 16071 19261
rect 22017 3383 22051 3689
rect 27169 3451 27203 3689
<< viali >>
rect 2697 117385 2731 117419
rect 23857 117385 23891 117419
rect 27261 117385 27295 117419
rect 29929 117385 29963 117419
rect 31125 117385 31159 117419
rect 34345 117385 34379 117419
rect 28549 117317 28583 117351
rect 2053 117249 2087 117283
rect 4537 117249 4571 117283
rect 6009 117249 6043 117283
rect 8585 117249 8619 117283
rect 9873 117249 9907 117283
rect 11345 117249 11379 117283
rect 13277 117249 13311 117283
rect 15209 117249 15243 117283
rect 16681 117249 16715 117283
rect 18613 117249 18647 117283
rect 20545 117249 20579 117283
rect 26617 117249 26651 117283
rect 31953 117249 31987 117283
rect 35357 117249 35391 117283
rect 36553 117249 36587 117283
rect 5273 117181 5307 117215
rect 7849 117181 7883 117215
rect 10609 117181 10643 117215
rect 12541 117181 12575 117215
rect 14013 117181 14047 117215
rect 15761 117181 15795 117215
rect 17693 117181 17727 117215
rect 19165 117181 19199 117215
rect 23029 117181 23063 117215
rect 26433 117181 26467 117215
rect 29837 117181 29871 117215
rect 32689 117181 32723 117215
rect 36369 117181 36403 117215
rect 37381 117181 37415 117215
rect 1869 117113 1903 117147
rect 2605 117113 2639 117147
rect 4353 117113 4387 117147
rect 5089 117113 5123 117147
rect 5825 117113 5859 117147
rect 7021 117113 7055 117147
rect 8401 117113 8435 117147
rect 9689 117113 9723 117147
rect 10425 117113 10459 117147
rect 11161 117113 11195 117147
rect 12357 117113 12391 117147
rect 13093 117113 13127 117147
rect 13829 117113 13863 117147
rect 15025 117113 15059 117147
rect 16497 117113 16531 117147
rect 18429 117113 18463 117147
rect 20361 117113 20395 117147
rect 21097 117113 21131 117147
rect 21833 117113 21867 117147
rect 23213 117113 23247 117147
rect 23765 117113 23799 117147
rect 24501 117113 24535 117147
rect 25697 117113 25731 117147
rect 27169 117113 27203 117147
rect 28365 117113 28399 117147
rect 29101 117113 29135 117147
rect 31033 117113 31067 117147
rect 31769 117113 31803 117147
rect 32505 117113 32539 117147
rect 34253 117113 34287 117147
rect 35173 117113 35207 117147
rect 37933 117113 37967 117147
rect 7113 117045 7147 117079
rect 15853 117045 15887 117079
rect 17785 117045 17819 117079
rect 19257 117045 19291 117079
rect 21189 117045 21223 117079
rect 21925 117045 21959 117079
rect 24593 117045 24627 117079
rect 25789 117045 25823 117079
rect 29193 117045 29227 117079
rect 1961 116841 1995 116875
rect 4169 116841 4203 116875
rect 7021 116841 7055 116875
rect 7757 116841 7791 116875
rect 9229 116841 9263 116875
rect 9965 116841 9999 116875
rect 12265 116841 12299 116875
rect 13001 116841 13035 116875
rect 14473 116841 14507 116875
rect 15945 116841 15979 116875
rect 17509 116841 17543 116875
rect 18245 116841 18279 116875
rect 19717 116841 19751 116875
rect 20453 116841 20487 116875
rect 21189 116841 21223 116875
rect 22753 116841 22787 116875
rect 24409 116841 24443 116875
rect 25145 116841 25179 116875
rect 26617 116841 26651 116875
rect 28733 116841 28767 116875
rect 31585 116841 31619 116875
rect 34805 116841 34839 116875
rect 35541 116841 35575 116875
rect 2789 116773 2823 116807
rect 4997 116773 5031 116807
rect 8401 116773 8435 116807
rect 10793 116773 10827 116807
rect 13829 116773 13863 116807
rect 15301 116773 15335 116807
rect 19073 116773 19107 116807
rect 22644 116773 22678 116807
rect 28089 116773 28123 116807
rect 33425 116773 33459 116807
rect 36369 116773 36403 116807
rect 1869 116705 1903 116739
rect 2605 116705 2639 116739
rect 3341 116705 3375 116739
rect 4077 116705 4111 116739
rect 4813 116705 4847 116739
rect 5549 116705 5583 116739
rect 6929 116705 6963 116739
rect 7665 116705 7699 116739
rect 9137 116705 9171 116739
rect 9873 116705 9907 116739
rect 10609 116705 10643 116739
rect 12173 116705 12207 116739
rect 12909 116705 12943 116739
rect 13645 116705 13679 116739
rect 14381 116705 14415 116739
rect 15117 116705 15151 116739
rect 15853 116705 15887 116739
rect 17417 116705 17451 116739
rect 18153 116705 18187 116739
rect 18889 116705 18923 116739
rect 19625 116705 19659 116739
rect 20361 116705 20395 116739
rect 21097 116705 21131 116739
rect 23397 116705 23431 116739
rect 24317 116705 24351 116739
rect 25053 116705 25087 116739
rect 25789 116705 25823 116739
rect 26525 116705 26559 116739
rect 27905 116705 27939 116739
rect 28641 116705 28675 116739
rect 29285 116705 29319 116739
rect 30941 116705 30975 116739
rect 33241 116705 33275 116739
rect 33977 116705 34011 116739
rect 34713 116705 34747 116739
rect 35449 116705 35483 116739
rect 36185 116705 36219 116739
rect 36921 116705 36955 116739
rect 5733 116637 5767 116671
rect 29653 116637 29687 116671
rect 31309 116637 31343 116671
rect 29745 116569 29779 116603
rect 34161 116569 34195 116603
rect 3433 116501 3467 116535
rect 8493 116501 8527 116535
rect 23489 116501 23523 116535
rect 25881 116501 25915 116535
rect 29423 116501 29457 116535
rect 29561 116501 29595 116535
rect 31079 116501 31113 116535
rect 31217 116501 31251 116535
rect 37013 116501 37047 116535
rect 2421 116297 2455 116331
rect 3157 116297 3191 116331
rect 5641 116297 5675 116331
rect 6377 116297 6411 116331
rect 7849 116297 7883 116331
rect 10609 116297 10643 116331
rect 11345 116297 11379 116331
rect 15761 116297 15795 116331
rect 20177 116297 20211 116331
rect 21465 116297 21499 116331
rect 22201 116297 22235 116331
rect 23305 116297 23339 116331
rect 24041 116297 24075 116331
rect 26065 116297 26099 116331
rect 27629 116297 27663 116331
rect 33333 116297 33367 116331
rect 35909 116297 35943 116331
rect 4997 116229 5031 116263
rect 7205 116229 7239 116263
rect 16589 116229 16623 116263
rect 25421 116229 25455 116263
rect 28457 116229 28491 116263
rect 30757 116229 30791 116263
rect 31953 116229 31987 116263
rect 33149 116229 33183 116263
rect 36737 116229 36771 116263
rect 9505 116161 9539 116195
rect 11897 116161 11931 116195
rect 13185 116161 13219 116195
rect 17049 116161 17083 116195
rect 30628 116161 30662 116195
rect 30849 116161 30883 116195
rect 30941 116161 30975 116195
rect 32045 116161 32079 116195
rect 33241 116161 33275 116195
rect 34805 116161 34839 116195
rect 37841 116161 37875 116195
rect 12541 116093 12575 116127
rect 14749 116093 14783 116127
rect 18337 116093 18371 116127
rect 20085 116093 20119 116127
rect 22109 116093 22143 116127
rect 23213 116093 23247 116127
rect 26617 116093 26651 116127
rect 26801 116093 26835 116127
rect 31824 116093 31858 116127
rect 33020 116093 33054 116127
rect 36553 116093 36587 116127
rect 37657 116093 37691 116127
rect 2329 116025 2363 116059
rect 3065 116025 3099 116059
rect 4813 116025 4847 116059
rect 5549 116025 5583 116059
rect 6285 116025 6319 116059
rect 7021 116025 7055 116059
rect 7757 116025 7791 116059
rect 10517 116025 10551 116059
rect 11253 116025 11287 116059
rect 15669 116025 15703 116059
rect 16405 116025 16439 116059
rect 17693 116025 17727 116059
rect 21373 116025 21407 116059
rect 23949 116025 23983 116059
rect 25973 116025 26007 116059
rect 26985 116025 27019 116059
rect 27537 116025 27571 116059
rect 28273 116025 28307 116059
rect 29009 116025 29043 116059
rect 30481 116025 30515 116059
rect 31677 116025 31711 116059
rect 32873 116025 32907 116059
rect 34621 116025 34655 116059
rect 35817 116025 35851 116059
rect 29101 115957 29135 115991
rect 32321 115957 32355 115991
rect 4445 115753 4479 115787
rect 5181 115753 5215 115787
rect 8309 115753 8343 115787
rect 8861 115753 8895 115787
rect 9505 115753 9539 115787
rect 10149 115753 10183 115787
rect 13369 115753 13403 115787
rect 14565 115753 14599 115787
rect 18429 115753 18463 115787
rect 26525 115753 26559 115787
rect 27997 115753 28031 115787
rect 29653 115753 29687 115787
rect 30389 115753 30423 115787
rect 30941 115753 30975 115787
rect 31585 115753 31619 115787
rect 36001 115753 36035 115787
rect 36737 115753 36771 115787
rect 2789 115685 2823 115719
rect 3801 115685 3835 115719
rect 10793 115685 10827 115719
rect 15209 115685 15243 115719
rect 19073 115685 19107 115719
rect 30297 115685 30331 115719
rect 33885 115685 33919 115719
rect 35357 115685 35391 115719
rect 1869 115617 1903 115651
rect 2605 115617 2639 115651
rect 3617 115617 3651 115651
rect 4353 115617 4387 115651
rect 5089 115617 5123 115651
rect 7021 115617 7055 115651
rect 8217 115617 8251 115651
rect 12265 115617 12299 115651
rect 12909 115617 12943 115651
rect 17509 115617 17543 115651
rect 20545 115617 20579 115651
rect 21189 115617 21223 115651
rect 22753 115617 22787 115651
rect 24041 115617 24075 115651
rect 24685 115617 24719 115651
rect 25513 115617 25547 115651
rect 26433 115617 26467 115651
rect 27905 115617 27939 115651
rect 28733 115617 28767 115651
rect 29561 115617 29595 115651
rect 31125 115617 31159 115651
rect 31769 115617 31803 115651
rect 33701 115617 33735 115651
rect 34437 115617 34471 115651
rect 35173 115617 35207 115651
rect 35909 115617 35943 115651
rect 36645 115617 36679 115651
rect 15853 115549 15887 115583
rect 19901 115481 19935 115515
rect 28549 115481 28583 115515
rect 34621 115481 34655 115515
rect 1961 115413 1995 115447
rect 23397 115413 23431 115447
rect 1961 115209 1995 115243
rect 4445 115209 4479 115243
rect 5089 115209 5123 115243
rect 7113 115209 7147 115243
rect 8125 115209 8159 115243
rect 9689 115209 9723 115243
rect 10333 115209 10367 115243
rect 10977 115209 11011 115243
rect 11621 115209 11655 115243
rect 13001 115209 13035 115243
rect 13645 115209 13679 115243
rect 14933 115209 14967 115243
rect 15577 115209 15611 115243
rect 16221 115209 16255 115243
rect 16865 115209 16899 115243
rect 17509 115209 17543 115243
rect 18797 115209 18831 115243
rect 20177 115209 20211 115243
rect 20637 115209 20671 115243
rect 21649 115209 21683 115243
rect 22109 115209 22143 115243
rect 25421 115209 25455 115243
rect 26065 115209 26099 115243
rect 27813 115209 27847 115243
rect 31125 115209 31159 115243
rect 31769 115209 31803 115243
rect 32413 115209 32447 115243
rect 34713 115209 34747 115243
rect 37105 115209 37139 115243
rect 2789 115141 2823 115175
rect 5825 115141 5859 115175
rect 22753 115141 22787 115175
rect 29009 115141 29043 115175
rect 34069 115141 34103 115175
rect 36461 115141 36495 115175
rect 6469 115073 6503 115107
rect 18153 115073 18187 115107
rect 33333 115073 33367 115107
rect 2605 115005 2639 115039
rect 12265 115005 12299 115039
rect 20821 115005 20855 115039
rect 22293 115005 22327 115039
rect 22937 115005 22971 115039
rect 23581 115005 23615 115039
rect 24317 115005 24351 115039
rect 26709 115005 26743 115039
rect 28549 115005 28583 115039
rect 29193 115005 29227 115039
rect 30665 115005 30699 115039
rect 31309 115005 31343 115039
rect 31953 115005 31987 115039
rect 32597 115005 32631 115039
rect 37657 115005 37691 115039
rect 1869 114937 1903 114971
rect 5641 114937 5675 114971
rect 8033 114937 8067 114971
rect 27721 114937 27755 114971
rect 33149 114937 33183 114971
rect 33885 114937 33919 114971
rect 34621 114937 34655 114971
rect 36277 114937 36311 114971
rect 37013 114937 37047 114971
rect 37933 114937 37967 114971
rect 12081 114869 12115 114903
rect 23397 114869 23431 114903
rect 24133 114869 24167 114903
rect 26525 114869 26559 114903
rect 28365 114869 28399 114903
rect 30481 114869 30515 114903
rect 10333 114665 10367 114699
rect 12725 114665 12759 114699
rect 14013 114665 14047 114699
rect 15945 114665 15979 114699
rect 17325 114665 17359 114699
rect 18245 114665 18279 114699
rect 20821 114665 20855 114699
rect 21465 114665 21499 114699
rect 22569 114665 22603 114699
rect 24041 114665 24075 114699
rect 27997 114665 28031 114699
rect 29285 114665 29319 114699
rect 30573 114665 30607 114699
rect 31953 114665 31987 114699
rect 1869 114597 1903 114631
rect 35725 114597 35759 114631
rect 35909 114597 35943 114631
rect 2605 114529 2639 114563
rect 3341 114529 3375 114563
rect 9229 114529 9263 114563
rect 9689 114529 9723 114563
rect 10517 114529 10551 114563
rect 11161 114529 11195 114563
rect 12265 114529 12299 114563
rect 12909 114529 12943 114563
rect 13553 114529 13587 114563
rect 14197 114529 14231 114563
rect 14841 114529 14875 114563
rect 15485 114529 15519 114563
rect 16129 114529 16163 114563
rect 17509 114529 17543 114563
rect 18061 114529 18095 114563
rect 18705 114529 18739 114563
rect 19533 114529 19567 114563
rect 19993 114529 20027 114563
rect 21005 114529 21039 114563
rect 21649 114529 21683 114563
rect 22753 114529 22787 114563
rect 23213 114529 23247 114563
rect 24225 114529 24259 114563
rect 25145 114529 25179 114563
rect 25789 114529 25823 114563
rect 26433 114529 26467 114563
rect 28181 114529 28215 114563
rect 28825 114529 28859 114563
rect 29469 114529 29503 114563
rect 30113 114529 30147 114563
rect 30757 114529 30791 114563
rect 31401 114529 31435 114563
rect 32137 114529 32171 114563
rect 33517 114529 33551 114563
rect 34253 114529 34287 114563
rect 34989 114529 35023 114563
rect 36461 114529 36495 114563
rect 37105 114529 37139 114563
rect 2053 114461 2087 114495
rect 2789 114461 2823 114495
rect 4169 114461 4203 114495
rect 5089 114461 5123 114495
rect 7021 114461 7055 114495
rect 7665 114461 7699 114495
rect 8585 114461 8619 114495
rect 33701 114461 33735 114495
rect 35173 114461 35207 114495
rect 36645 114461 36679 114495
rect 12081 114393 12115 114427
rect 15301 114393 15335 114427
rect 18889 114393 18923 114427
rect 19349 114393 19383 114427
rect 24961 114393 24995 114427
rect 25605 114393 25639 114427
rect 26249 114393 26283 114427
rect 29929 114393 29963 114427
rect 31217 114393 31251 114427
rect 34437 114393 34471 114427
rect 3433 114325 3467 114359
rect 5733 114325 5767 114359
rect 9045 114325 9079 114359
rect 9873 114325 9907 114359
rect 10977 114325 11011 114359
rect 13369 114325 13403 114359
rect 14657 114325 14691 114359
rect 28641 114325 28675 114359
rect 37289 114325 37323 114359
rect 3065 114121 3099 114155
rect 4445 114121 4479 114155
rect 5825 114121 5859 114155
rect 7021 114121 7055 114155
rect 9505 114121 9539 114155
rect 18337 114121 18371 114155
rect 21557 114121 21591 114155
rect 25237 114121 25271 114155
rect 26249 114121 26283 114155
rect 29285 114121 29319 114155
rect 30481 114121 30515 114155
rect 31769 114121 31803 114155
rect 32505 114121 32539 114155
rect 33701 114121 33735 114155
rect 34713 114121 34747 114155
rect 38025 114121 38059 114155
rect 5089 114053 5123 114087
rect 8125 114053 8159 114087
rect 15761 114053 15795 114087
rect 17693 114053 17727 114087
rect 31125 114053 31159 114087
rect 36645 114053 36679 114087
rect 37381 113985 37415 114019
rect 7665 113917 7699 113951
rect 8309 113917 8343 113951
rect 9689 113917 9723 113951
rect 15945 113917 15979 113951
rect 16589 113917 16623 113951
rect 17877 113917 17911 113951
rect 18521 113917 18555 113951
rect 20177 113917 20211 113951
rect 20821 113917 20855 113951
rect 21741 113917 21775 113951
rect 22201 113917 22235 113951
rect 22845 113917 22879 113951
rect 23489 113917 23523 113951
rect 24133 113917 24167 113951
rect 25421 113917 25455 113951
rect 26433 113917 26467 113951
rect 29469 113917 29503 113951
rect 30665 113917 30699 113951
rect 31309 113917 31343 113951
rect 31953 113917 31987 113951
rect 32689 113917 32723 113951
rect 33885 113917 33919 113951
rect 37197 113917 37231 113951
rect 1869 113849 1903 113883
rect 34621 113849 34655 113883
rect 36461 113849 36495 113883
rect 37933 113849 37967 113883
rect 1961 113781 1995 113815
rect 7481 113781 7515 113815
rect 16405 113781 16439 113815
rect 4629 113577 4663 113611
rect 6837 113577 6871 113611
rect 30757 113577 30791 113611
rect 33057 113577 33091 113611
rect 35081 113577 35115 113611
rect 35909 113509 35943 113543
rect 36645 113509 36679 113543
rect 1501 113441 1535 113475
rect 2329 113441 2363 113475
rect 2973 113441 3007 113475
rect 3433 113441 3467 113475
rect 4813 113441 4847 113475
rect 5457 113441 5491 113475
rect 7021 113441 7055 113475
rect 7665 113441 7699 113475
rect 8301 113441 8335 113475
rect 8769 113441 8803 113475
rect 24593 113441 24627 113475
rect 25237 113441 25271 113475
rect 30941 113441 30975 113475
rect 31585 113441 31619 113475
rect 33241 113441 33275 113475
rect 33885 113441 33919 113475
rect 34989 113441 35023 113475
rect 35725 113441 35759 113475
rect 36461 113441 36495 113475
rect 37197 113441 37231 113475
rect 5273 113305 5307 113339
rect 7481 113305 7515 113339
rect 8125 113305 8159 113339
rect 31401 113305 31435 113339
rect 33701 113305 33735 113339
rect 37381 113305 37415 113339
rect 31401 113033 31435 113067
rect 33333 113033 33367 113067
rect 33977 113033 34011 113067
rect 36553 113033 36587 113067
rect 28273 112965 28307 112999
rect 1869 112829 1903 112863
rect 2697 112829 2731 112863
rect 4261 112829 4295 112863
rect 4905 112829 4939 112863
rect 5549 112829 5583 112863
rect 6193 112829 6227 112863
rect 6837 112829 6871 112863
rect 7481 112829 7515 112863
rect 28181 112829 28215 112863
rect 28457 112829 28491 112863
rect 31585 112829 31619 112863
rect 33517 112829 33551 112863
rect 34161 112829 34195 112863
rect 37197 112829 37231 112863
rect 37933 112829 37967 112863
rect 36461 112761 36495 112795
rect 37381 112761 37415 112795
rect 38117 112761 38151 112795
rect 2145 112693 2179 112727
rect 28641 112693 28675 112727
rect 36553 112489 36587 112523
rect 37381 112421 37415 112455
rect 1869 112353 1903 112387
rect 36461 112353 36495 112387
rect 37197 112353 37231 112387
rect 1961 112149 1995 112183
rect 37657 111741 37691 111775
rect 37933 111673 37967 111707
rect 31769 111401 31803 111435
rect 36553 111401 36587 111435
rect 1409 111265 1443 111299
rect 31585 111265 31619 111299
rect 36461 111265 36495 111299
rect 37197 111265 37231 111299
rect 1685 111197 1719 111231
rect 37381 111129 37415 111163
rect 37473 110653 37507 110687
rect 1869 110585 1903 110619
rect 37841 110585 37875 110619
rect 1961 110517 1995 110551
rect 37197 110177 37231 110211
rect 37381 110041 37415 110075
rect 2053 109565 2087 109599
rect 37197 109565 37231 109599
rect 1869 109497 1903 109531
rect 37933 109497 37967 109531
rect 38117 109497 38151 109531
rect 37289 109429 37323 109463
rect 8677 109225 8711 109259
rect 8493 109089 8527 109123
rect 37197 109089 37231 109123
rect 37381 109021 37415 109055
rect 1961 108681 1995 108715
rect 38117 108477 38151 108511
rect 1869 108409 1903 108443
rect 37933 108409 37967 108443
rect 1869 108001 1903 108035
rect 37197 108001 37231 108035
rect 2053 107865 2087 107899
rect 37289 107797 37323 107831
rect 37197 107389 37231 107423
rect 37381 107321 37415 107355
rect 37933 107321 37967 107355
rect 38025 107253 38059 107287
rect 1961 107049 1995 107083
rect 1869 106913 1903 106947
rect 37197 106913 37231 106947
rect 37381 106777 37415 106811
rect 1685 106369 1719 106403
rect 37565 106369 37599 106403
rect 1777 106301 1811 106335
rect 1961 106301 1995 106335
rect 37289 106301 37323 106335
rect 37197 105825 37231 105859
rect 37289 105621 37323 105655
rect 26341 105417 26375 105451
rect 32229 105417 32263 105451
rect 1409 105213 1443 105247
rect 25237 105213 25271 105247
rect 25697 105213 25731 105247
rect 26065 105213 26099 105247
rect 32045 105213 32079 105247
rect 37197 105213 37231 105247
rect 37933 105145 37967 105179
rect 1593 105077 1627 105111
rect 37289 105077 37323 105111
rect 38025 105077 38059 105111
rect 25973 104873 26007 104907
rect 1869 104737 1903 104771
rect 24869 104737 24903 104771
rect 25329 104737 25363 104771
rect 25697 104737 25731 104771
rect 37197 104737 37231 104771
rect 1961 104533 1995 104567
rect 37289 104533 37323 104567
rect 29561 104329 29595 104363
rect 29377 104125 29411 104159
rect 37197 104057 37231 104091
rect 37381 104057 37415 104091
rect 37933 104057 37967 104091
rect 38025 103989 38059 104023
rect 12541 103785 12575 103819
rect 21281 103785 21315 103819
rect 21649 103785 21683 103819
rect 1869 103717 1903 103751
rect 21490 103717 21524 103751
rect 25145 103717 25179 103751
rect 12541 103649 12575 103683
rect 13093 103649 13127 103683
rect 13277 103649 13311 103683
rect 24961 103649 24995 103683
rect 37197 103649 37231 103683
rect 21005 103581 21039 103615
rect 21373 103581 21407 103615
rect 37381 103581 37415 103615
rect 2053 103513 2087 103547
rect 6377 103241 6411 103275
rect 7021 103173 7055 103207
rect 26617 103173 26651 103207
rect 37565 103105 37599 103139
rect 6193 103037 6227 103071
rect 6837 103037 6871 103071
rect 37289 103037 37323 103071
rect 1869 102969 1903 103003
rect 2053 102969 2087 103003
rect 26433 102969 26467 103003
rect 7849 102697 7883 102731
rect 12449 102697 12483 102731
rect 26801 102697 26835 102731
rect 7665 102561 7699 102595
rect 12357 102561 12391 102595
rect 26709 102561 26743 102595
rect 37197 102561 37231 102595
rect 12081 102493 12115 102527
rect 12566 102493 12600 102527
rect 12725 102425 12759 102459
rect 37289 102357 37323 102391
rect 11897 102085 11931 102119
rect 13461 102085 13495 102119
rect 11529 102017 11563 102051
rect 13185 102017 13219 102051
rect 1869 101949 1903 101983
rect 11253 101949 11287 101983
rect 12817 101949 12851 101983
rect 2053 101881 2087 101915
rect 11738 101881 11772 101915
rect 13302 101881 13336 101915
rect 37933 101881 37967 101915
rect 11621 101813 11655 101847
rect 13093 101813 13127 101847
rect 38025 101813 38059 101847
rect 5917 101609 5951 101643
rect 12449 101609 12483 101643
rect 12725 101609 12759 101643
rect 23305 101609 23339 101643
rect 12357 101541 12391 101575
rect 1869 101473 1903 101507
rect 5733 101473 5767 101507
rect 12081 101473 12115 101507
rect 23213 101473 23247 101507
rect 37197 101473 37231 101507
rect 12566 101405 12600 101439
rect 2053 101337 2087 101371
rect 37289 101269 37323 101303
rect 37933 100861 37967 100895
rect 37197 100793 37231 100827
rect 37381 100793 37415 100827
rect 38025 100725 38059 100759
rect 23121 100521 23155 100555
rect 1869 100453 1903 100487
rect 23029 100385 23063 100419
rect 37197 100385 37231 100419
rect 1961 100181 1995 100215
rect 37289 100181 37323 100215
rect 34713 99977 34747 100011
rect 33977 99909 34011 99943
rect 33793 99773 33827 99807
rect 34621 99773 34655 99807
rect 1869 99705 1903 99739
rect 2053 99705 2087 99739
rect 21925 99705 21959 99739
rect 22109 99705 22143 99739
rect 33609 99705 33643 99739
rect 34437 99705 34471 99739
rect 37933 99705 37967 99739
rect 38025 99637 38059 99671
rect 13277 99297 13311 99331
rect 37197 99297 37231 99331
rect 12909 99229 12943 99263
rect 13185 99229 13219 99263
rect 13369 99229 13403 99263
rect 13553 99093 13587 99127
rect 37289 99093 37323 99127
rect 21465 98821 21499 98855
rect 22201 98821 22235 98855
rect 1869 98685 1903 98719
rect 37197 98685 37231 98719
rect 2053 98617 2087 98651
rect 21281 98617 21315 98651
rect 22017 98617 22051 98651
rect 37381 98617 37415 98651
rect 37933 98617 37967 98651
rect 38025 98549 38059 98583
rect 5181 98345 5215 98379
rect 1869 98209 1903 98243
rect 4997 98209 5031 98243
rect 37197 98209 37231 98243
rect 2053 98073 2087 98107
rect 37289 98005 37323 98039
rect 16589 97733 16623 97767
rect 16405 97597 16439 97631
rect 37933 97597 37967 97631
rect 14841 97529 14875 97563
rect 15117 97461 15151 97495
rect 38025 97461 38059 97495
rect 1869 97121 1903 97155
rect 37197 97121 37231 97155
rect 1961 96917 1995 96951
rect 37289 96917 37323 96951
rect 18337 96713 18371 96747
rect 18245 96509 18279 96543
rect 37197 96509 37231 96543
rect 37933 96509 37967 96543
rect 1869 96441 1903 96475
rect 18061 96441 18095 96475
rect 38117 96441 38151 96475
rect 1961 96373 1995 96407
rect 37381 96373 37415 96407
rect 37197 96033 37231 96067
rect 37381 95829 37415 95863
rect 1961 95625 1995 95659
rect 38117 95557 38151 95591
rect 1869 95421 1903 95455
rect 22845 95421 22879 95455
rect 23305 95421 23339 95455
rect 23673 95421 23707 95455
rect 37289 95421 37323 95455
rect 37933 95421 37967 95455
rect 23949 95285 23983 95319
rect 37473 95285 37507 95319
rect 1869 94945 1903 94979
rect 37197 94945 37231 94979
rect 1961 94741 1995 94775
rect 37381 94741 37415 94775
rect 38117 94469 38151 94503
rect 37289 94333 37323 94367
rect 37933 94333 37967 94367
rect 37473 94197 37507 94231
rect 1869 93857 1903 93891
rect 2053 93857 2087 93891
rect 37289 93245 37323 93279
rect 37933 93245 37967 93279
rect 38945 93245 38979 93279
rect 1869 93177 1903 93211
rect 1961 93109 1995 93143
rect 37473 93109 37507 93143
rect 38117 93109 38151 93143
rect 37197 92769 37231 92803
rect 37381 92565 37415 92599
rect 38945 92497 38979 92531
rect 20177 92361 20211 92395
rect 38117 92293 38151 92327
rect 1869 92157 1903 92191
rect 37289 92157 37323 92191
rect 37933 92157 37967 92191
rect 20085 92089 20119 92123
rect 1961 92021 1995 92055
rect 37473 92021 37507 92055
rect 10885 91817 10919 91851
rect 15853 91817 15887 91851
rect 1869 91681 1903 91715
rect 10793 91681 10827 91715
rect 15761 91681 15795 91715
rect 1961 91477 1995 91511
rect 38117 91273 38151 91307
rect 37473 91205 37507 91239
rect 33057 91137 33091 91171
rect 28365 91069 28399 91103
rect 28458 91069 28492 91103
rect 28641 91069 28675 91103
rect 28871 91069 28905 91103
rect 32597 91069 32631 91103
rect 32689 91069 32723 91103
rect 32965 91069 32999 91103
rect 37289 91069 37323 91103
rect 37933 91069 37967 91103
rect 28733 91001 28767 91035
rect 31953 91001 31987 91035
rect 29009 90933 29043 90967
rect 18245 90729 18279 90763
rect 28641 90661 28675 90695
rect 1869 90593 1903 90627
rect 18153 90593 18187 90627
rect 28365 90593 28399 90627
rect 28458 90593 28492 90627
rect 28733 90593 28767 90627
rect 28871 90593 28905 90627
rect 31585 90593 31619 90627
rect 31953 90593 31987 90627
rect 32137 90593 32171 90627
rect 33057 90593 33091 90627
rect 37197 90593 37231 90627
rect 31677 90525 31711 90559
rect 1961 90389 1995 90423
rect 29009 90389 29043 90423
rect 31033 90389 31067 90423
rect 33241 90389 33275 90423
rect 37381 90389 37415 90423
rect 38117 90117 38151 90151
rect 32781 90049 32815 90083
rect 33149 90049 33183 90083
rect 18705 89981 18739 90015
rect 28365 89981 28399 90015
rect 28458 89981 28492 90015
rect 28641 89981 28675 90015
rect 28830 89981 28864 90015
rect 32689 89981 32723 90015
rect 33057 89981 33091 90015
rect 37289 89981 37323 90015
rect 37933 89981 37967 90015
rect 19073 89913 19107 89947
rect 28733 89913 28767 89947
rect 32045 89913 32079 89947
rect 29009 89845 29043 89879
rect 37473 89845 37507 89879
rect 28917 89641 28951 89675
rect 1869 89573 1903 89607
rect 28273 89505 28307 89539
rect 28366 89505 28400 89539
rect 28549 89505 28583 89539
rect 28641 89505 28675 89539
rect 28779 89505 28813 89539
rect 31585 89505 31619 89539
rect 31953 89505 31987 89539
rect 32137 89505 32171 89539
rect 33701 89505 33735 89539
rect 34069 89505 34103 89539
rect 34161 89505 34195 89539
rect 31493 89437 31527 89471
rect 33609 89437 33643 89471
rect 2053 89369 2087 89403
rect 31033 89301 31067 89335
rect 33149 89301 33183 89335
rect 28917 89097 28951 89131
rect 33057 88961 33091 88995
rect 23581 88893 23615 88927
rect 28273 88893 28307 88927
rect 28366 88893 28400 88927
rect 28779 88893 28813 88927
rect 32597 88893 32631 88927
rect 32689 88893 32723 88927
rect 32965 88893 32999 88927
rect 37289 88893 37323 88927
rect 37933 88893 37967 88927
rect 1869 88825 1903 88859
rect 2053 88825 2087 88859
rect 23765 88825 23799 88859
rect 28549 88825 28583 88859
rect 28641 88825 28675 88859
rect 31953 88825 31987 88859
rect 37473 88757 37507 88791
rect 38117 88757 38151 88791
rect 28733 88553 28767 88587
rect 37381 88553 37415 88587
rect 28089 88417 28123 88451
rect 28182 88417 28216 88451
rect 28365 88417 28399 88451
rect 28457 88417 28491 88451
rect 28595 88417 28629 88451
rect 29193 88417 29227 88451
rect 29286 88417 29320 88451
rect 29469 88417 29503 88451
rect 29561 88417 29595 88451
rect 29699 88417 29733 88451
rect 30941 88417 30975 88451
rect 31585 88417 31619 88451
rect 31953 88417 31987 88451
rect 32137 88417 32171 88451
rect 33701 88417 33735 88451
rect 33793 88417 33827 88451
rect 34069 88417 34103 88451
rect 34253 88417 34287 88451
rect 37197 88417 37231 88451
rect 31493 88349 31527 88383
rect 29837 88213 29871 88247
rect 33149 88213 33183 88247
rect 28733 88009 28767 88043
rect 27629 87941 27663 87975
rect 30941 87941 30975 87975
rect 38117 87941 38151 87975
rect 32045 87873 32079 87907
rect 32597 87873 32631 87907
rect 1869 87805 1903 87839
rect 26985 87805 27019 87839
rect 27078 87805 27112 87839
rect 27491 87805 27525 87839
rect 28089 87805 28123 87839
rect 28182 87805 28216 87839
rect 28595 87805 28629 87839
rect 30757 87805 30791 87839
rect 32137 87805 32171 87839
rect 32505 87805 32539 87839
rect 37289 87805 37323 87839
rect 37933 87805 37967 87839
rect 2053 87737 2087 87771
rect 27261 87737 27295 87771
rect 27353 87737 27387 87771
rect 28365 87737 28399 87771
rect 28457 87737 28491 87771
rect 31493 87737 31527 87771
rect 33241 87737 33275 87771
rect 33333 87669 33367 87703
rect 37473 87669 37507 87703
rect 28641 87465 28675 87499
rect 33241 87465 33275 87499
rect 28365 87397 28399 87431
rect 29285 87397 29319 87431
rect 1869 87329 1903 87363
rect 23397 87329 23431 87363
rect 27997 87329 28031 87363
rect 28090 87329 28124 87363
rect 28273 87329 28307 87363
rect 28503 87329 28537 87363
rect 29929 87329 29963 87363
rect 30297 87329 30331 87363
rect 30481 87329 30515 87363
rect 31585 87329 31619 87363
rect 31953 87329 31987 87363
rect 33057 87329 33091 87363
rect 30021 87261 30055 87295
rect 31493 87261 31527 87295
rect 32045 87261 32079 87295
rect 23581 87193 23615 87227
rect 1961 87125 1995 87159
rect 31033 87125 31067 87159
rect 26801 86921 26835 86955
rect 27537 86921 27571 86955
rect 23029 86717 23063 86751
rect 23213 86717 23247 86751
rect 23949 86717 23983 86751
rect 31585 86785 31619 86819
rect 32137 86785 32171 86819
rect 26893 86717 26927 86751
rect 26986 86717 27020 86751
rect 27169 86717 27203 86751
rect 27261 86717 27295 86751
rect 27399 86717 27433 86751
rect 27997 86717 28031 86751
rect 28090 86717 28124 86751
rect 28365 86717 28399 86751
rect 28503 86717 28537 86751
rect 31677 86717 31711 86751
rect 32045 86717 32079 86751
rect 32965 86717 32999 86751
rect 33057 86717 33091 86751
rect 33241 86717 33275 86751
rect 33333 86717 33367 86751
rect 33793 86717 33827 86751
rect 37289 86717 37323 86751
rect 37933 86717 37967 86751
rect 22569 86649 22603 86683
rect 22661 86649 22695 86683
rect 23121 86649 23155 86683
rect 24133 86649 24167 86683
rect 26801 86649 26835 86683
rect 28273 86649 28307 86683
rect 31033 86649 31067 86683
rect 28641 86581 28675 86615
rect 32781 86581 32815 86615
rect 33977 86581 34011 86615
rect 37473 86581 37507 86615
rect 38117 86581 38151 86615
rect 19993 86377 20027 86411
rect 26801 86377 26835 86411
rect 28641 86377 28675 86411
rect 29745 86377 29779 86411
rect 33241 86377 33275 86411
rect 1869 86309 1903 86343
rect 29469 86309 29503 86343
rect 19901 86241 19935 86275
rect 23397 86241 23431 86275
rect 26709 86241 26743 86275
rect 27997 86241 28031 86275
rect 28090 86241 28124 86275
rect 28273 86241 28307 86275
rect 28365 86241 28399 86275
rect 28503 86241 28537 86275
rect 29101 86241 29135 86275
rect 29194 86241 29228 86275
rect 29377 86241 29411 86275
rect 29605 86241 29639 86275
rect 30205 86241 30239 86275
rect 31507 86241 31541 86275
rect 31953 86241 31987 86275
rect 33057 86241 33091 86275
rect 37197 86241 37231 86275
rect 31585 86173 31619 86207
rect 32045 86173 32079 86207
rect 2053 86105 2087 86139
rect 30389 86105 30423 86139
rect 23581 86037 23615 86071
rect 31033 86037 31067 86071
rect 37381 86037 37415 86071
rect 37473 85765 37507 85799
rect 1869 85629 1903 85663
rect 27813 85629 27847 85663
rect 27906 85629 27940 85663
rect 28089 85629 28123 85663
rect 28319 85629 28353 85663
rect 28917 85629 28951 85663
rect 29065 85629 29099 85663
rect 29285 85629 29319 85663
rect 29423 85629 29457 85663
rect 31401 85629 31435 85663
rect 31493 85629 31527 85663
rect 31769 85629 31803 85663
rect 31953 85629 31987 85663
rect 32689 85629 32723 85663
rect 32781 85629 32815 85663
rect 32965 85629 32999 85663
rect 33057 85629 33091 85663
rect 33517 85629 33551 85663
rect 37289 85629 37323 85663
rect 37933 85629 37967 85663
rect 2053 85561 2087 85595
rect 28181 85561 28215 85595
rect 29193 85561 29227 85595
rect 30757 85561 30791 85595
rect 28457 85493 28491 85527
rect 29561 85493 29595 85527
rect 32505 85493 32539 85527
rect 33701 85493 33735 85527
rect 38117 85493 38151 85527
rect 26801 85289 26835 85323
rect 30205 85289 30239 85323
rect 33517 85289 33551 85323
rect 28089 85221 28123 85255
rect 29193 85221 29227 85255
rect 23213 85153 23247 85187
rect 26709 85153 26743 85187
rect 27813 85153 27847 85187
rect 27906 85153 27940 85187
rect 28181 85153 28215 85187
rect 28319 85153 28353 85187
rect 28917 85153 28951 85187
rect 29010 85153 29044 85187
rect 29285 85153 29319 85187
rect 29423 85153 29457 85187
rect 30021 85153 30055 85187
rect 31401 85153 31435 85187
rect 31769 85153 31803 85187
rect 33425 85153 33459 85187
rect 31493 85085 31527 85119
rect 31861 85085 31895 85119
rect 23397 85017 23431 85051
rect 29561 85017 29595 85051
rect 30849 85017 30883 85051
rect 28457 84949 28491 84983
rect 29193 84677 29227 84711
rect 38117 84677 38151 84711
rect 31585 84609 31619 84643
rect 32689 84609 32723 84643
rect 1869 84541 1903 84575
rect 27813 84541 27847 84575
rect 27906 84541 27940 84575
rect 28181 84541 28215 84575
rect 28319 84541 28353 84575
rect 29009 84541 29043 84575
rect 31125 84541 31159 84575
rect 31217 84541 31251 84575
rect 31493 84541 31527 84575
rect 32781 84541 32815 84575
rect 33149 84541 33183 84575
rect 33333 84541 33367 84575
rect 37289 84541 37323 84575
rect 37933 84541 37967 84575
rect 2053 84473 2087 84507
rect 28089 84473 28123 84507
rect 30481 84473 30515 84507
rect 32137 84473 32171 84507
rect 28457 84405 28491 84439
rect 37473 84405 37507 84439
rect 28457 84201 28491 84235
rect 28089 84133 28123 84167
rect 1869 84065 1903 84099
rect 27813 84065 27847 84099
rect 27906 84065 27940 84099
rect 28181 84065 28215 84099
rect 28278 84065 28312 84099
rect 28917 84065 28951 84099
rect 29653 84065 29687 84099
rect 31033 84065 31067 84099
rect 31401 84065 31435 84099
rect 31585 84065 31619 84099
rect 37197 84065 37231 84099
rect 30941 83997 30975 84031
rect 2053 83929 2087 83963
rect 29101 83861 29135 83895
rect 29837 83861 29871 83895
rect 30481 83861 30515 83895
rect 37381 83861 37415 83895
rect 30573 83657 30607 83691
rect 29469 83589 29503 83623
rect 27537 83453 27571 83487
rect 27630 83453 27664 83487
rect 27813 83453 27847 83487
rect 28043 83453 28077 83487
rect 29285 83453 29319 83487
rect 31125 83453 31159 83487
rect 31217 83453 31251 83487
rect 31493 83453 31527 83487
rect 31677 83453 31711 83487
rect 37289 83453 37323 83487
rect 37933 83453 37967 83487
rect 27905 83385 27939 83419
rect 28181 83317 28215 83351
rect 37473 83317 37507 83351
rect 38117 83317 38151 83351
rect 28089 83045 28123 83079
rect 1409 82977 1443 83011
rect 27813 82977 27847 83011
rect 27906 82977 27940 83011
rect 28181 82977 28215 83011
rect 28278 82977 28312 83011
rect 30665 82977 30699 83011
rect 31033 82977 31067 83011
rect 31125 82977 31159 83011
rect 1685 82909 1719 82943
rect 30021 82909 30055 82943
rect 30757 82909 30791 82943
rect 28457 82841 28491 82875
rect 27997 82569 28031 82603
rect 29101 82569 29135 82603
rect 37473 82501 37507 82535
rect 31585 82433 31619 82467
rect 27353 82365 27387 82399
rect 27446 82365 27480 82399
rect 27859 82365 27893 82399
rect 28457 82365 28491 82399
rect 28550 82365 28584 82399
rect 28733 82365 28767 82399
rect 28963 82365 28997 82399
rect 31125 82365 31159 82399
rect 31217 82365 31251 82399
rect 31493 82365 31527 82399
rect 37289 82365 37323 82399
rect 37933 82365 37967 82399
rect 1869 82297 1903 82331
rect 27629 82297 27663 82331
rect 27721 82297 27755 82331
rect 28825 82297 28859 82331
rect 30481 82297 30515 82331
rect 1961 82229 1995 82263
rect 38117 82229 38151 82263
rect 28733 81889 28767 81923
rect 29101 81889 29135 81923
rect 29193 81889 29227 81923
rect 30389 81889 30423 81923
rect 30757 81889 30791 81923
rect 37197 81889 37231 81923
rect 28641 81821 28675 81855
rect 30481 81821 30515 81855
rect 30849 81821 30883 81855
rect 29837 81753 29871 81787
rect 28181 81685 28215 81719
rect 37381 81685 37415 81719
rect 29469 81345 29503 81379
rect 31585 81345 31619 81379
rect 1869 81277 1903 81311
rect 29009 81277 29043 81311
rect 29101 81277 29135 81311
rect 29377 81277 29411 81311
rect 31125 81277 31159 81311
rect 31217 81277 31251 81311
rect 31493 81277 31527 81311
rect 32781 81277 32815 81311
rect 32873 81277 32907 81311
rect 33149 81277 33183 81311
rect 33333 81277 33367 81311
rect 37289 81277 37323 81311
rect 37933 81277 37967 81311
rect 2053 81209 2087 81243
rect 28365 81209 28399 81243
rect 30481 81209 30515 81243
rect 32137 81209 32171 81243
rect 37473 81141 37507 81175
rect 38117 81141 38151 81175
rect 1409 80801 1443 80835
rect 27813 80801 27847 80835
rect 27906 80801 27940 80835
rect 28089 80801 28123 80835
rect 28181 80801 28215 80835
rect 28319 80801 28353 80835
rect 30205 80801 30239 80835
rect 30573 80801 30607 80835
rect 30757 80801 30791 80835
rect 31309 80801 31343 80835
rect 31493 80801 31527 80835
rect 31585 80801 31619 80835
rect 31769 80801 31803 80835
rect 31856 80801 31890 80835
rect 30113 80733 30147 80767
rect 28457 80665 28491 80699
rect 1593 80597 1627 80631
rect 29653 80597 29687 80631
rect 27813 80393 27847 80427
rect 30849 80393 30883 80427
rect 28917 80325 28951 80359
rect 27169 80189 27203 80223
rect 27262 80189 27296 80223
rect 27675 80189 27709 80223
rect 28273 80189 28307 80223
rect 28366 80189 28400 80223
rect 28549 80189 28583 80223
rect 28779 80189 28813 80223
rect 27445 80121 27479 80155
rect 27537 80121 27571 80155
rect 28641 80121 28675 80155
rect 30849 80121 30883 80155
rect 30941 80325 30975 80359
rect 37473 80325 37507 80359
rect 31309 80189 31343 80223
rect 31401 80189 31435 80223
rect 31585 80189 31619 80223
rect 31677 80189 31711 80223
rect 37289 80189 37323 80223
rect 37933 80189 37967 80223
rect 30941 80053 30975 80087
rect 31125 80053 31159 80087
rect 38117 80053 38151 80087
rect 26525 79781 26559 79815
rect 28089 79781 28123 79815
rect 28181 79781 28215 79815
rect 1409 79713 1443 79747
rect 26249 79713 26283 79747
rect 26342 79713 26376 79747
rect 26617 79713 26651 79747
rect 26714 79713 26748 79747
rect 27813 79713 27847 79747
rect 27933 79713 27967 79747
rect 28319 79713 28353 79747
rect 30205 79713 30239 79747
rect 30573 79713 30607 79747
rect 37197 79713 37231 79747
rect 30297 79645 30331 79679
rect 30665 79645 30699 79679
rect 28457 79577 28491 79611
rect 37381 79577 37415 79611
rect 1593 79509 1627 79543
rect 26893 79509 26927 79543
rect 29653 79509 29687 79543
rect 38117 79305 38151 79339
rect 28825 79237 28859 79271
rect 29561 79237 29595 79271
rect 27077 79101 27111 79135
rect 27170 79101 27204 79135
rect 27445 79101 27479 79135
rect 27583 79101 27617 79135
rect 28181 79101 28215 79135
rect 28274 79101 28308 79135
rect 28549 79101 28583 79135
rect 28687 79101 28721 79135
rect 37933 79101 37967 79135
rect 1869 79033 1903 79067
rect 2053 79033 2087 79067
rect 27353 79033 27387 79067
rect 28457 79033 28491 79067
rect 29377 79033 29411 79067
rect 27721 78965 27755 78999
rect 28089 78693 28123 78727
rect 37197 78693 37231 78727
rect 27813 78625 27847 78659
rect 27906 78625 27940 78659
rect 28181 78625 28215 78659
rect 28319 78625 28353 78659
rect 29469 78625 29503 78659
rect 29193 78557 29227 78591
rect 28457 78489 28491 78523
rect 37289 78421 37323 78455
rect 29377 78217 29411 78251
rect 1869 78013 1903 78047
rect 28089 78013 28123 78047
rect 37197 78013 37231 78047
rect 29285 77945 29319 77979
rect 37933 77945 37967 77979
rect 1961 77877 1995 77911
rect 28181 77877 28215 77911
rect 37289 77877 37323 77911
rect 38025 77877 38059 77911
rect 1409 77537 1443 77571
rect 37197 77537 37231 77571
rect 1593 77333 1627 77367
rect 37289 77333 37323 77367
rect 25513 77061 25547 77095
rect 29285 77061 29319 77095
rect 25329 76857 25363 76891
rect 29101 76857 29135 76891
rect 37933 76857 37967 76891
rect 38025 76789 38059 76823
rect 1409 76449 1443 76483
rect 24777 76449 24811 76483
rect 37197 76449 37231 76483
rect 1593 76245 1627 76279
rect 24961 76245 24995 76279
rect 37289 76245 37323 76279
rect 25237 75837 25271 75871
rect 37197 75837 37231 75871
rect 1869 75769 1903 75803
rect 37933 75769 37967 75803
rect 1961 75701 1995 75735
rect 25421 75701 25455 75735
rect 37289 75701 37323 75735
rect 38025 75701 38059 75735
rect 37197 75361 37231 75395
rect 37289 75157 37323 75191
rect 1869 74749 1903 74783
rect 2053 74681 2087 74715
rect 37933 74681 37967 74715
rect 38025 74613 38059 74647
rect 1869 74273 1903 74307
rect 37197 74273 37231 74307
rect 2053 74137 2087 74171
rect 37289 74069 37323 74103
rect 29377 73865 29411 73899
rect 29193 73661 29227 73695
rect 37197 73661 37231 73695
rect 37933 73593 37967 73627
rect 37289 73525 37323 73559
rect 38025 73525 38059 73559
rect 1869 73185 1903 73219
rect 2053 73185 2087 73219
rect 37197 73185 37231 73219
rect 37289 72981 37323 73015
rect 37933 72573 37967 72607
rect 1869 72505 1903 72539
rect 2053 72505 2087 72539
rect 38025 72437 38059 72471
rect 37197 72097 37231 72131
rect 37381 71961 37415 71995
rect 33977 71689 34011 71723
rect 1869 71485 1903 71519
rect 33793 71485 33827 71519
rect 37197 71485 37231 71519
rect 37381 71485 37415 71519
rect 2053 71417 2087 71451
rect 37933 71417 37967 71451
rect 38117 71417 38151 71451
rect 1869 71009 1903 71043
rect 37197 71009 37231 71043
rect 2053 70873 2087 70907
rect 37381 70873 37415 70907
rect 38117 70465 38151 70499
rect 37933 70397 37967 70431
rect 1869 69921 1903 69955
rect 37197 69921 37231 69955
rect 2053 69785 2087 69819
rect 37289 69717 37323 69751
rect 37381 69377 37415 69411
rect 38117 69309 38151 69343
rect 37197 69241 37231 69275
rect 37933 69241 37967 69275
rect 1869 68901 1903 68935
rect 37197 68833 37231 68867
rect 2053 68697 2087 68731
rect 37381 68629 37415 68663
rect 1869 68221 1903 68255
rect 37289 68221 37323 68255
rect 37933 68221 37967 68255
rect 38945 68221 38979 68255
rect 2053 68153 2087 68187
rect 37473 68085 37507 68119
rect 38117 68085 38151 68119
rect 37197 67745 37231 67779
rect 37381 67609 37415 67643
rect 38945 67609 38979 67643
rect 37473 67269 37507 67303
rect 1409 67133 1443 67167
rect 37289 67133 37323 67167
rect 37933 67133 37967 67167
rect 1593 66997 1627 67031
rect 38117 66997 38151 67031
rect 1409 66657 1443 66691
rect 1593 66453 1627 66487
rect 37473 66181 37507 66215
rect 37289 66045 37323 66079
rect 37933 66045 37967 66079
rect 38117 65909 38151 65943
rect 1409 65569 1443 65603
rect 37197 65569 37231 65603
rect 1593 65365 1627 65399
rect 37381 65365 37415 65399
rect 1593 65093 1627 65127
rect 37473 65093 37507 65127
rect 1409 64957 1443 64991
rect 37289 64957 37323 64991
rect 37933 64957 37967 64991
rect 38117 64821 38151 64855
rect 34621 64617 34655 64651
rect 34345 64481 34379 64515
rect 34529 64481 34563 64515
rect 15301 64073 15335 64107
rect 34253 64073 34287 64107
rect 1409 63869 1443 63903
rect 34161 63869 34195 63903
rect 37289 63869 37323 63903
rect 37933 63869 37967 63903
rect 15209 63801 15243 63835
rect 33977 63801 34011 63835
rect 1593 63733 1627 63767
rect 37473 63733 37507 63767
rect 38117 63733 38151 63767
rect 35449 63529 35483 63563
rect 36461 63529 36495 63563
rect 34713 63461 34747 63495
rect 36185 63461 36219 63495
rect 1409 63393 1443 63427
rect 33149 63393 33183 63427
rect 33333 63393 33367 63427
rect 33701 63393 33735 63427
rect 34161 63393 34195 63427
rect 34345 63393 34379 63427
rect 35173 63393 35207 63427
rect 35357 63393 35391 63427
rect 36369 63393 36403 63427
rect 37197 63393 37231 63427
rect 1593 63189 1627 63223
rect 37381 63189 37415 63223
rect 33057 62985 33091 63019
rect 34069 62985 34103 63019
rect 32965 62781 32999 62815
rect 33977 62781 34011 62815
rect 37289 62781 37323 62815
rect 37933 62781 37967 62815
rect 32781 62713 32815 62747
rect 33793 62713 33827 62747
rect 37473 62645 37507 62679
rect 38117 62645 38151 62679
rect 30021 62441 30055 62475
rect 34069 62373 34103 62407
rect 1409 62305 1443 62339
rect 29929 62305 29963 62339
rect 30757 62305 30791 62339
rect 30941 62305 30975 62339
rect 33425 62305 33459 62339
rect 33517 62305 33551 62339
rect 33701 62305 33735 62339
rect 34805 62305 34839 62339
rect 34989 62305 35023 62339
rect 35357 62305 35391 62339
rect 1593 62101 1627 62135
rect 33425 62101 33459 62135
rect 1409 61693 1443 61727
rect 37289 61693 37323 61727
rect 37933 61693 37967 61727
rect 1593 61557 1627 61591
rect 37473 61557 37507 61591
rect 38117 61557 38151 61591
rect 37197 61217 37231 61251
rect 37381 61013 37415 61047
rect 34437 60809 34471 60843
rect 1409 60605 1443 60639
rect 25973 60605 26007 60639
rect 26157 60605 26191 60639
rect 26341 60605 26375 60639
rect 26525 60605 26559 60639
rect 34253 60605 34287 60639
rect 37289 60605 37323 60639
rect 37933 60605 37967 60639
rect 1593 60469 1627 60503
rect 25973 60469 26007 60503
rect 37473 60469 37507 60503
rect 38117 60469 38151 60503
rect 1409 60129 1443 60163
rect 37197 60129 37231 60163
rect 1593 59925 1627 59959
rect 37381 59925 37415 59959
rect 37105 59653 37139 59687
rect 26249 59517 26283 59551
rect 26525 59517 26559 59551
rect 26801 59517 26835 59551
rect 26985 59517 27019 59551
rect 36921 59517 36955 59551
rect 37565 59517 37599 59551
rect 37749 59517 37783 59551
rect 37979 59517 38013 59551
rect 37837 59449 37871 59483
rect 26341 59381 26375 59415
rect 38117 59381 38151 59415
rect 10241 59109 10275 59143
rect 1409 59041 1443 59075
rect 12265 59041 12299 59075
rect 36461 59041 36495 59075
rect 37197 59041 37231 59075
rect 10425 58973 10459 59007
rect 12081 58973 12115 59007
rect 37381 58905 37415 58939
rect 1593 58837 1627 58871
rect 12449 58837 12483 58871
rect 36645 58837 36679 58871
rect 27169 58633 27203 58667
rect 12817 58497 12851 58531
rect 1409 58429 1443 58463
rect 12081 58429 12115 58463
rect 12173 58429 12207 58463
rect 13001 58429 13035 58463
rect 26617 58429 26651 58463
rect 26893 58429 26927 58463
rect 26985 58429 27019 58463
rect 36553 58429 36587 58463
rect 36829 58429 36863 58463
rect 36921 58429 36955 58463
rect 37565 58429 37599 58463
rect 37841 58429 37875 58463
rect 37933 58429 37967 58463
rect 26801 58361 26835 58395
rect 36737 58361 36771 58395
rect 37749 58361 37783 58395
rect 38945 58361 38979 58395
rect 1593 58293 1627 58327
rect 12357 58293 12391 58327
rect 13185 58293 13219 58327
rect 37105 58293 37139 58327
rect 38117 58293 38151 58327
rect 12081 57953 12115 57987
rect 12265 57953 12299 57987
rect 12449 57953 12483 57987
rect 36461 57953 36495 57987
rect 37197 57953 37231 57987
rect 37381 57817 37415 57851
rect 36553 57749 36587 57783
rect 27169 57545 27203 57579
rect 37105 57477 37139 57511
rect 1409 57341 1443 57375
rect 26617 57341 26651 57375
rect 26801 57341 26835 57375
rect 26893 57341 26927 57375
rect 27031 57341 27065 57375
rect 29193 57341 29227 57375
rect 36921 57341 36955 57375
rect 37565 57341 37599 57375
rect 37933 57341 37967 57375
rect 29009 57273 29043 57307
rect 37749 57273 37783 57307
rect 37841 57273 37875 57307
rect 38945 57273 38979 57307
rect 1593 57205 1627 57239
rect 38117 57205 38151 57239
rect 26617 56933 26651 56967
rect 36461 56933 36495 56967
rect 1409 56865 1443 56899
rect 26249 56865 26283 56899
rect 26341 56865 26375 56899
rect 26479 56865 26513 56899
rect 26733 56865 26767 56899
rect 37197 56865 37231 56899
rect 36645 56797 36679 56831
rect 26893 56729 26927 56763
rect 37381 56729 37415 56763
rect 1593 56661 1627 56695
rect 26249 56661 26283 56695
rect 27261 56457 27295 56491
rect 36829 56457 36863 56491
rect 37473 56457 37507 56491
rect 26709 56253 26743 56287
rect 26985 56253 27019 56287
rect 27077 56253 27111 56287
rect 36185 56253 36219 56287
rect 36278 56253 36312 56287
rect 36461 56253 36495 56287
rect 36691 56253 36725 56287
rect 26893 56185 26927 56219
rect 36553 56185 36587 56219
rect 37381 56185 37415 56219
rect 35633 55913 35667 55947
rect 36461 55845 36495 55879
rect 1409 55777 1443 55811
rect 34805 55777 34839 55811
rect 35541 55777 35575 55811
rect 36185 55777 36219 55811
rect 36278 55777 36312 55811
rect 36553 55777 36587 55811
rect 36691 55777 36725 55811
rect 36829 55641 36863 55675
rect 1593 55573 1627 55607
rect 34989 55573 35023 55607
rect 29193 55369 29227 55403
rect 1409 55165 1443 55199
rect 29101 55165 29135 55199
rect 34621 55165 34655 55199
rect 36185 55165 36219 55199
rect 36333 55165 36367 55199
rect 36691 55165 36725 55199
rect 37565 55165 37599 55199
rect 37933 55165 37967 55199
rect 36461 55097 36495 55131
rect 36553 55097 36587 55131
rect 37749 55097 37783 55131
rect 37841 55097 37875 55131
rect 1593 55029 1627 55063
rect 34805 55029 34839 55063
rect 36829 55029 36863 55063
rect 38117 55029 38151 55063
rect 35725 54825 35759 54859
rect 36461 54757 36495 54791
rect 35541 54689 35575 54723
rect 36185 54689 36219 54723
rect 36278 54689 36312 54723
rect 36553 54689 36587 54723
rect 36691 54689 36725 54723
rect 36829 54485 36863 54519
rect 36277 54281 36311 54315
rect 36921 54213 36955 54247
rect 1409 54077 1443 54111
rect 36461 54077 36495 54111
rect 37105 54077 37139 54111
rect 37565 54077 37599 54111
rect 37933 54077 37967 54111
rect 37749 54009 37783 54043
rect 37841 54009 37875 54043
rect 1593 53941 1627 53975
rect 38117 53941 38151 53975
rect 36553 53737 36587 53771
rect 37197 53737 37231 53771
rect 1409 53601 1443 53635
rect 36737 53601 36771 53635
rect 37381 53601 37415 53635
rect 1593 53397 1627 53431
rect 27077 53193 27111 53227
rect 36093 53125 36127 53159
rect 26525 52989 26559 53023
rect 26898 52989 26932 53023
rect 35909 52989 35943 53023
rect 36553 52989 36587 53023
rect 36921 52989 36955 53023
rect 37565 52989 37599 53023
rect 37749 52989 37783 53023
rect 37933 52989 37967 53023
rect 26709 52921 26743 52955
rect 26801 52921 26835 52955
rect 36737 52921 36771 52955
rect 36829 52921 36863 52955
rect 37841 52921 37875 52955
rect 37105 52853 37139 52887
rect 38117 52853 38151 52887
rect 36553 52649 36587 52683
rect 37197 52649 37231 52683
rect 1869 52513 1903 52547
rect 36737 52513 36771 52547
rect 37381 52513 37415 52547
rect 2053 52445 2087 52479
rect 2053 52037 2087 52071
rect 27077 52037 27111 52071
rect 26525 51901 26559 51935
rect 26801 51901 26835 51935
rect 26898 51901 26932 51935
rect 37565 51901 37599 51935
rect 37933 51901 37967 51935
rect 1869 51833 1903 51867
rect 26709 51833 26743 51867
rect 37749 51833 37783 51867
rect 37841 51833 37875 51867
rect 38117 51765 38151 51799
rect 19809 51561 19843 51595
rect 23121 51561 23155 51595
rect 24961 51561 24995 51595
rect 29837 51561 29871 51595
rect 37197 51561 37231 51595
rect 26525 51493 26559 51527
rect 28825 51493 28859 51527
rect 34989 51493 35023 51527
rect 19533 51425 19567 51459
rect 23029 51425 23063 51459
rect 24685 51425 24719 51459
rect 26249 51425 26283 51459
rect 26433 51425 26467 51459
rect 26622 51425 26656 51459
rect 27905 51425 27939 51459
rect 29193 51425 29227 51459
rect 29745 51425 29779 51459
rect 34621 51425 34655 51459
rect 36553 51425 36587 51459
rect 37381 51425 37415 51459
rect 36737 51289 36771 51323
rect 26801 51221 26835 51255
rect 28181 51221 28215 51255
rect 20729 51017 20763 51051
rect 22569 51017 22603 51051
rect 23581 51017 23615 51051
rect 25421 51017 25455 51051
rect 27077 51017 27111 51051
rect 30849 51017 30883 51051
rect 32873 51017 32907 51051
rect 37933 51017 37967 51051
rect 2053 50949 2087 50983
rect 1869 50813 1903 50847
rect 23489 50813 23523 50847
rect 26525 50813 26559 50847
rect 26898 50813 26932 50847
rect 28273 50813 28307 50847
rect 28549 50813 28583 50847
rect 28825 50813 28859 50847
rect 28917 50813 28951 50847
rect 36737 50813 36771 50847
rect 36830 50813 36864 50847
rect 37013 50813 37047 50847
rect 37241 50813 37275 50847
rect 38117 50813 38151 50847
rect 20453 50745 20487 50779
rect 22477 50745 22511 50779
rect 25329 50745 25363 50779
rect 26709 50745 26743 50779
rect 26801 50745 26835 50779
rect 30573 50745 30607 50779
rect 32781 50745 32815 50779
rect 37105 50745 37139 50779
rect 28365 50677 28399 50711
rect 37381 50677 37415 50711
rect 25329 50473 25363 50507
rect 7297 50337 7331 50371
rect 25237 50337 25271 50371
rect 36093 50337 36127 50371
rect 36737 50337 36771 50371
rect 36885 50337 36919 50371
rect 37013 50337 37047 50371
rect 37105 50337 37139 50371
rect 37243 50337 37277 50371
rect 36277 50201 36311 50235
rect 7481 50133 7515 50167
rect 37381 50133 37415 50167
rect 27077 49929 27111 49963
rect 36093 49929 36127 49963
rect 37933 49929 37967 49963
rect 2053 49861 2087 49895
rect 1869 49725 1903 49759
rect 26525 49725 26559 49759
rect 26898 49725 26932 49759
rect 36277 49725 36311 49759
rect 36737 49725 36771 49759
rect 36830 49725 36864 49759
rect 37013 49725 37047 49759
rect 37243 49725 37277 49759
rect 38117 49725 38151 49759
rect 26709 49657 26743 49691
rect 26801 49657 26835 49691
rect 37105 49657 37139 49691
rect 37381 49589 37415 49623
rect 2053 49317 2087 49351
rect 36921 49317 36955 49351
rect 1869 49249 1903 49283
rect 23121 49249 23155 49283
rect 23397 49249 23431 49283
rect 23857 49249 23891 49283
rect 35633 49249 35667 49283
rect 35817 49249 35851 49283
rect 35909 49249 35943 49283
rect 36001 49249 36035 49283
rect 36645 49249 36679 49283
rect 36738 49249 36772 49283
rect 37013 49249 37047 49283
rect 37151 49249 37185 49283
rect 23949 49181 23983 49215
rect 24225 49113 24259 49147
rect 36185 49045 36219 49079
rect 37289 49045 37323 49079
rect 36001 48841 36035 48875
rect 38025 48841 38059 48875
rect 7205 48637 7239 48671
rect 36185 48637 36219 48671
rect 36645 48637 36679 48671
rect 36738 48637 36772 48671
rect 37151 48637 37185 48671
rect 36921 48569 36955 48603
rect 37013 48569 37047 48603
rect 37933 48569 37967 48603
rect 7389 48501 7423 48535
rect 37289 48501 37323 48535
rect 1869 48229 1903 48263
rect 2053 48229 2087 48263
rect 37013 48229 37047 48263
rect 37105 48229 37139 48263
rect 8769 48161 8803 48195
rect 35541 48161 35575 48195
rect 36369 48161 36403 48195
rect 36829 48161 36863 48195
rect 37197 48161 37231 48195
rect 8585 48093 8619 48127
rect 35725 48025 35759 48059
rect 36185 48025 36219 48059
rect 8953 47957 8987 47991
rect 37381 47957 37415 47991
rect 26893 47753 26927 47787
rect 36093 47753 36127 47787
rect 1685 47617 1719 47651
rect 8217 47617 8251 47651
rect 9505 47617 9539 47651
rect 1409 47549 1443 47583
rect 7113 47549 7147 47583
rect 8401 47549 8435 47583
rect 9689 47549 9723 47583
rect 26341 47549 26375 47583
rect 26714 47549 26748 47583
rect 35909 47549 35943 47583
rect 36553 47549 36587 47583
rect 36829 47549 36863 47583
rect 36921 47549 36955 47583
rect 37565 47549 37599 47583
rect 37841 47549 37875 47583
rect 37933 47549 37967 47583
rect 8585 47481 8619 47515
rect 26525 47481 26559 47515
rect 26617 47481 26651 47515
rect 36737 47481 36771 47515
rect 37749 47481 37783 47515
rect 7297 47413 7331 47447
rect 9873 47413 9907 47447
rect 37105 47413 37139 47447
rect 38117 47413 38151 47447
rect 35449 47209 35483 47243
rect 35909 47209 35943 47243
rect 26525 47141 26559 47175
rect 7573 47073 7607 47107
rect 8401 47073 8435 47107
rect 9229 47073 9263 47107
rect 10057 47073 10091 47107
rect 26249 47073 26283 47107
rect 26433 47073 26467 47107
rect 26622 47073 26656 47107
rect 35265 47073 35299 47107
rect 36093 47073 36127 47107
rect 36553 47073 36587 47107
rect 7389 47005 7423 47039
rect 8217 47005 8251 47039
rect 9045 47005 9079 47039
rect 9873 47005 9907 47039
rect 7757 46937 7791 46971
rect 8585 46937 8619 46971
rect 10241 46937 10275 46971
rect 26801 46937 26835 46971
rect 36737 46937 36771 46971
rect 9413 46869 9447 46903
rect 26893 46665 26927 46699
rect 36185 46597 36219 46631
rect 37105 46597 37139 46631
rect 1409 46529 1443 46563
rect 1685 46529 1719 46563
rect 7021 46461 7055 46495
rect 8217 46461 8251 46495
rect 8401 46461 8435 46495
rect 9505 46461 9539 46495
rect 9689 46461 9723 46495
rect 26341 46461 26375 46495
rect 26714 46461 26748 46495
rect 36369 46461 36403 46495
rect 37565 46461 37599 46495
rect 37933 46461 37967 46495
rect 26525 46393 26559 46427
rect 26617 46393 26651 46427
rect 36921 46393 36955 46427
rect 37749 46393 37783 46427
rect 37841 46393 37875 46427
rect 7205 46325 7239 46359
rect 8585 46325 8619 46359
rect 9873 46325 9907 46359
rect 38117 46325 38151 46359
rect 35265 46121 35299 46155
rect 35909 46121 35943 46155
rect 37197 46121 37231 46155
rect 2053 46053 2087 46087
rect 1869 45985 1903 46019
rect 9137 45985 9171 46019
rect 26249 45985 26283 46019
rect 26433 45985 26467 46019
rect 26525 45985 26559 46019
rect 26622 45985 26656 46019
rect 35449 45985 35483 46019
rect 36093 45985 36127 46019
rect 36553 45985 36587 46019
rect 36701 45985 36735 46019
rect 36829 45985 36863 46019
rect 36921 45985 36955 46019
rect 37057 45985 37091 46019
rect 8953 45917 8987 45951
rect 26801 45849 26835 45883
rect 9321 45781 9355 45815
rect 7757 45577 7791 45611
rect 37841 45577 37875 45611
rect 36001 45509 36035 45543
rect 8217 45441 8251 45475
rect 7573 45373 7607 45407
rect 8401 45373 8435 45407
rect 9505 45373 9539 45407
rect 9689 45373 9723 45407
rect 26341 45373 26375 45407
rect 26714 45373 26748 45407
rect 35817 45373 35851 45407
rect 36461 45373 36495 45407
rect 36554 45373 36588 45407
rect 36737 45373 36771 45407
rect 36967 45373 37001 45407
rect 37749 45373 37783 45407
rect 26525 45305 26559 45339
rect 26617 45305 26651 45339
rect 26910 45305 26944 45339
rect 36829 45305 36863 45339
rect 8585 45237 8619 45271
rect 9873 45237 9907 45271
rect 37105 45237 37139 45271
rect 24225 45033 24259 45067
rect 34713 45033 34747 45067
rect 35357 45033 35391 45067
rect 1869 44965 1903 44999
rect 2053 44965 2087 44999
rect 26893 44965 26927 44999
rect 28917 44965 28951 44999
rect 8033 44897 8067 44931
rect 8861 44897 8895 44931
rect 9689 44897 9723 44931
rect 10517 44897 10551 44931
rect 24041 44897 24075 44931
rect 26709 44897 26743 44931
rect 29745 44897 29779 44931
rect 29929 44897 29963 44931
rect 30205 44897 30239 44931
rect 34529 44897 34563 44931
rect 35173 44897 35207 44931
rect 35817 44897 35851 44931
rect 36461 44897 36495 44931
rect 36554 44897 36588 44931
rect 36737 44897 36771 44931
rect 36829 44897 36863 44931
rect 36967 44897 37001 44931
rect 7849 44829 7883 44863
rect 8677 44829 8711 44863
rect 9505 44829 9539 44863
rect 10333 44829 10367 44863
rect 29837 44829 29871 44863
rect 30021 44829 30055 44863
rect 9873 44761 9907 44795
rect 8217 44693 8251 44727
rect 9045 44693 9079 44727
rect 10701 44693 10735 44727
rect 29009 44693 29043 44727
rect 29561 44693 29595 44727
rect 36001 44693 36035 44727
rect 37105 44693 37139 44727
rect 26985 44489 27019 44523
rect 34621 44489 34655 44523
rect 35909 44489 35943 44523
rect 2053 44421 2087 44455
rect 29193 44421 29227 44455
rect 38117 44421 38151 44455
rect 9505 44353 9539 44387
rect 1869 44285 1903 44319
rect 7389 44285 7423 44319
rect 7573 44285 7607 44319
rect 8217 44285 8251 44319
rect 8401 44285 8435 44319
rect 9689 44285 9723 44319
rect 29101 44285 29135 44319
rect 29285 44285 29319 44319
rect 29377 44285 29411 44319
rect 29561 44285 29595 44319
rect 34805 44285 34839 44319
rect 36461 44285 36495 44319
rect 36554 44285 36588 44319
rect 36737 44285 36771 44319
rect 36967 44285 37001 44319
rect 37565 44285 37599 44319
rect 37749 44285 37783 44319
rect 37933 44285 37967 44319
rect 8585 44217 8619 44251
rect 26893 44217 26927 44251
rect 28273 44217 28307 44251
rect 35817 44217 35851 44251
rect 36829 44217 36863 44251
rect 37841 44217 37875 44251
rect 7757 44149 7791 44183
rect 9873 44149 9907 44183
rect 28365 44149 28399 44183
rect 28917 44149 28951 44183
rect 37105 44149 37139 44183
rect 9229 43945 9263 43979
rect 29285 43945 29319 43979
rect 35265 43945 35299 43979
rect 37013 43945 37047 43979
rect 8217 43809 8251 43843
rect 8401 43809 8435 43843
rect 9045 43809 9079 43843
rect 36645 43877 36679 43911
rect 29561 43809 29595 43843
rect 29837 43809 29871 43843
rect 30033 43809 30067 43843
rect 35081 43809 35115 43843
rect 35909 43809 35943 43843
rect 36369 43809 36403 43843
rect 36517 43809 36551 43843
rect 36737 43809 36771 43843
rect 36834 43809 36868 43843
rect 29754 43741 29788 43775
rect 29285 43673 29319 43707
rect 29653 43673 29687 43707
rect 8585 43605 8619 43639
rect 29377 43605 29411 43639
rect 35725 43605 35759 43639
rect 27077 43401 27111 43435
rect 34621 43401 34655 43435
rect 36829 43401 36863 43435
rect 2053 43265 2087 43299
rect 1869 43197 1903 43231
rect 26525 43197 26559 43231
rect 26898 43197 26932 43231
rect 29101 43197 29135 43231
rect 29193 43197 29227 43231
rect 29285 43197 29319 43231
rect 29377 43197 29411 43231
rect 29561 43197 29595 43231
rect 34805 43197 34839 43231
rect 35725 43197 35759 43231
rect 37565 43197 37599 43231
rect 37749 43197 37783 43231
rect 37979 43197 38013 43231
rect 26709 43129 26743 43163
rect 26801 43129 26835 43163
rect 36737 43129 36771 43163
rect 37841 43129 37875 43163
rect 28917 43061 28951 43095
rect 35909 43061 35943 43095
rect 38117 43061 38151 43095
rect 26433 42789 26467 42823
rect 26525 42789 26559 42823
rect 37105 42789 37139 42823
rect 1869 42721 1903 42755
rect 2053 42721 2087 42755
rect 26249 42721 26283 42755
rect 26645 42721 26679 42755
rect 26818 42721 26852 42755
rect 34897 42721 34931 42755
rect 35725 42721 35759 42755
rect 36185 42721 36219 42755
rect 36829 42721 36863 42755
rect 37013 42721 37047 42755
rect 37243 42721 37277 42755
rect 35081 42585 35115 42619
rect 35541 42585 35575 42619
rect 36369 42517 36403 42551
rect 37381 42517 37415 42551
rect 25973 42313 26007 42347
rect 28365 42313 28399 42347
rect 34621 42313 34655 42347
rect 26525 42177 26559 42211
rect 37289 42177 37323 42211
rect 7941 42109 7975 42143
rect 8125 42109 8159 42143
rect 26801 42109 26835 42143
rect 27813 42109 27847 42143
rect 27997 42109 28031 42143
rect 28089 42109 28123 42143
rect 28186 42109 28220 42143
rect 29009 42109 29043 42143
rect 34805 42109 34839 42143
rect 36277 42109 36311 42143
rect 36461 42109 36495 42143
rect 36553 42109 36587 42143
rect 36645 42109 36679 42143
rect 37565 42109 37599 42143
rect 25881 42041 25915 42075
rect 8309 41973 8343 42007
rect 29101 41973 29135 42007
rect 36829 41973 36863 42007
rect 34621 41769 34655 41803
rect 35449 41769 35483 41803
rect 36093 41769 36127 41803
rect 1869 41701 1903 41735
rect 26433 41701 26467 41735
rect 28825 41701 28859 41735
rect 36001 41701 36035 41735
rect 8125 41633 8159 41667
rect 8953 41633 8987 41667
rect 26249 41633 26283 41667
rect 26525 41633 26559 41667
rect 26622 41633 26656 41667
rect 29561 41633 29595 41667
rect 34805 41633 34839 41667
rect 35265 41633 35299 41667
rect 36737 41633 36771 41667
rect 7941 41565 7975 41599
rect 8769 41565 8803 41599
rect 36921 41565 36955 41599
rect 2053 41497 2087 41531
rect 26801 41497 26835 41531
rect 29745 41497 29779 41531
rect 8309 41429 8343 41463
rect 9137 41429 9171 41463
rect 28917 41429 28951 41463
rect 27077 41225 27111 41259
rect 34805 41225 34839 41259
rect 36185 41225 36219 41259
rect 2053 41157 2087 41191
rect 9505 41089 9539 41123
rect 1869 41021 1903 41055
rect 7941 41021 7975 41055
rect 8033 41021 8067 41055
rect 9689 41021 9723 41055
rect 26525 41021 26559 41055
rect 26898 41021 26932 41055
rect 34621 41021 34655 41055
rect 36185 41021 36219 41055
rect 36277 41021 36311 41055
rect 36370 41021 36404 41055
rect 36742 41021 36776 41055
rect 37565 41021 37599 41055
rect 37841 41021 37875 41055
rect 37933 41021 37967 41055
rect 26709 40953 26743 40987
rect 26801 40953 26835 40987
rect 28733 40953 28767 40987
rect 36553 40953 36587 40987
rect 36645 40953 36679 40987
rect 37749 40953 37783 40987
rect 8217 40885 8251 40919
rect 9873 40885 9907 40919
rect 28825 40885 28859 40919
rect 36921 40885 36955 40919
rect 38117 40885 38151 40919
rect 24869 40681 24903 40715
rect 35633 40681 35667 40715
rect 24225 40613 24259 40647
rect 29000 40613 29034 40647
rect 36553 40613 36587 40647
rect 8033 40545 8067 40579
rect 8677 40545 8711 40579
rect 8861 40545 8895 40579
rect 22569 40545 22603 40579
rect 24685 40545 24719 40579
rect 35173 40545 35207 40579
rect 35817 40545 35851 40579
rect 36277 40545 36311 40579
rect 36370 40545 36404 40579
rect 36645 40545 36679 40579
rect 36742 40545 36776 40579
rect 7849 40477 7883 40511
rect 22845 40477 22879 40511
rect 28733 40477 28767 40511
rect 34989 40409 35023 40443
rect 8217 40341 8251 40375
rect 9045 40341 9079 40375
rect 30113 40341 30147 40375
rect 36921 40341 36955 40375
rect 36185 40069 36219 40103
rect 2053 40001 2087 40035
rect 8033 40001 8067 40035
rect 1869 39933 1903 39967
rect 8217 39933 8251 39967
rect 28089 39933 28123 39967
rect 28356 39933 28390 39967
rect 34621 39933 34655 39967
rect 36185 39933 36219 39967
rect 36277 39933 36311 39967
rect 36370 39933 36404 39967
rect 36553 39933 36587 39967
rect 36742 39933 36776 39967
rect 37565 39933 37599 39967
rect 37749 39933 37783 39967
rect 37933 39933 37967 39967
rect 36645 39865 36679 39899
rect 37841 39865 37875 39899
rect 8401 39797 8435 39831
rect 29469 39797 29503 39831
rect 34805 39797 34839 39831
rect 36921 39797 36955 39831
rect 38117 39797 38151 39831
rect 1961 39593 1995 39627
rect 35081 39593 35115 39627
rect 28448 39525 28482 39559
rect 30380 39525 30414 39559
rect 36553 39525 36587 39559
rect 1869 39457 1903 39491
rect 30113 39457 30147 39491
rect 34437 39457 34471 39491
rect 34897 39457 34931 39491
rect 35633 39457 35667 39491
rect 36277 39457 36311 39491
rect 36425 39457 36459 39491
rect 36645 39457 36679 39491
rect 36742 39457 36776 39491
rect 28181 39389 28215 39423
rect 31493 39321 31527 39355
rect 34253 39321 34287 39355
rect 36921 39321 36955 39355
rect 29561 39253 29595 39287
rect 35725 39253 35759 39287
rect 23581 39049 23615 39083
rect 29469 39049 29503 39083
rect 34805 39049 34839 39083
rect 36185 39049 36219 39083
rect 22293 38981 22327 39015
rect 21649 38845 21683 38879
rect 21797 38845 21831 38879
rect 22114 38845 22148 38879
rect 23029 38845 23063 38879
rect 23397 38845 23431 38879
rect 25237 38845 25271 38879
rect 25421 38845 25455 38879
rect 28641 38845 28675 38879
rect 29377 38845 29411 38879
rect 34621 38845 34655 38879
rect 36185 38845 36219 38879
rect 36277 38845 36311 38879
rect 36425 38845 36459 38879
rect 36742 38845 36776 38879
rect 37565 38845 37599 38879
rect 37933 38845 37967 38879
rect 21925 38777 21959 38811
rect 22017 38777 22051 38811
rect 23213 38777 23247 38811
rect 23305 38777 23339 38811
rect 36553 38777 36587 38811
rect 36645 38777 36679 38811
rect 37749 38777 37783 38811
rect 37841 38777 37875 38811
rect 25329 38709 25363 38743
rect 28733 38709 28767 38743
rect 36921 38709 36955 38743
rect 38117 38709 38151 38743
rect 34805 38505 34839 38539
rect 35449 38505 35483 38539
rect 36277 38505 36311 38539
rect 1869 38437 1903 38471
rect 2053 38437 2087 38471
rect 22845 38437 22879 38471
rect 22937 38437 22971 38471
rect 24124 38437 24158 38471
rect 26433 38437 26467 38471
rect 37013 38437 37047 38471
rect 22569 38369 22603 38403
rect 22707 38369 22741 38403
rect 23075 38369 23109 38403
rect 26249 38369 26283 38403
rect 26525 38369 26559 38403
rect 26622 38369 26656 38403
rect 28917 38369 28951 38403
rect 29101 38369 29135 38403
rect 29377 38369 29411 38403
rect 34989 38369 35023 38403
rect 35633 38369 35667 38403
rect 36185 38369 36219 38403
rect 36829 38369 36863 38403
rect 37105 38369 37139 38403
rect 37197 38369 37231 38403
rect 23857 38301 23891 38335
rect 29193 38301 29227 38335
rect 23213 38233 23247 38267
rect 26801 38233 26835 38267
rect 29009 38233 29043 38267
rect 25237 38165 25271 38199
rect 28733 38165 28767 38199
rect 37381 38165 37415 38199
rect 26801 37961 26835 37995
rect 36369 37961 36403 37995
rect 2053 37893 2087 37927
rect 22385 37893 22419 37927
rect 23489 37893 23523 37927
rect 28825 37893 28859 37927
rect 38117 37893 38151 37927
rect 28917 37825 28951 37859
rect 29009 37825 29043 37859
rect 21741 37757 21775 37791
rect 21889 37757 21923 37791
rect 22206 37757 22240 37791
rect 22845 37757 22879 37791
rect 22938 37757 22972 37791
rect 23310 37757 23344 37791
rect 24133 37757 24167 37791
rect 24317 37757 24351 37791
rect 26249 37757 26283 37791
rect 26525 37757 26559 37791
rect 26622 37757 26656 37791
rect 28733 37757 28767 37791
rect 29193 37757 29227 37791
rect 36185 37757 36219 37791
rect 36921 37757 36955 37791
rect 37565 37757 37599 37791
rect 37749 37757 37783 37791
rect 37933 37757 37967 37791
rect 1869 37689 1903 37723
rect 22017 37689 22051 37723
rect 22109 37689 22143 37723
rect 23121 37689 23155 37723
rect 23213 37689 23247 37723
rect 26433 37689 26467 37723
rect 37105 37689 37139 37723
rect 37841 37689 37875 37723
rect 24225 37621 24259 37655
rect 28549 37621 28583 37655
rect 28365 37417 28399 37451
rect 35725 37417 35759 37451
rect 36185 37417 36219 37451
rect 24133 37349 24167 37383
rect 24338 37349 24372 37383
rect 26433 37349 26467 37383
rect 26525 37349 26559 37383
rect 37105 37349 37139 37383
rect 22937 37281 22971 37315
rect 23213 37281 23247 37315
rect 26249 37281 26283 37315
rect 26622 37281 26656 37315
rect 28549 37281 28583 37315
rect 28733 37281 28767 37315
rect 28825 37281 28859 37315
rect 29009 37281 29043 37315
rect 29653 37281 29687 37315
rect 29837 37281 29871 37315
rect 30113 37281 30147 37315
rect 35541 37281 35575 37315
rect 36369 37281 36403 37315
rect 36829 37281 36863 37315
rect 37013 37281 37047 37315
rect 37197 37281 37231 37315
rect 23581 37213 23615 37247
rect 29745 37213 29779 37247
rect 29929 37213 29963 37247
rect 23029 37145 23063 37179
rect 24501 37145 24535 37179
rect 26801 37145 26835 37179
rect 28641 37145 28675 37179
rect 24317 37077 24351 37111
rect 29469 37077 29503 37111
rect 37381 37077 37415 37111
rect 1593 36873 1627 36907
rect 23489 36873 23523 36907
rect 26801 36873 26835 36907
rect 35725 36873 35759 36907
rect 38117 36873 38151 36907
rect 21557 36737 21591 36771
rect 23949 36737 23983 36771
rect 28457 36737 28491 36771
rect 28549 36737 28583 36771
rect 1409 36669 1443 36703
rect 21281 36669 21315 36703
rect 23673 36669 23707 36703
rect 23765 36669 23799 36703
rect 24041 36669 24075 36703
rect 26249 36669 26283 36703
rect 26525 36669 26559 36703
rect 26622 36669 26656 36703
rect 28365 36669 28399 36703
rect 28641 36669 28675 36703
rect 28825 36669 28859 36703
rect 35725 36669 35759 36703
rect 35909 36669 35943 36703
rect 36553 36669 36587 36703
rect 36967 36669 37001 36703
rect 37565 36669 37599 36703
rect 37933 36669 37967 36703
rect 26433 36601 26467 36635
rect 36737 36601 36771 36635
rect 36829 36601 36863 36635
rect 37749 36601 37783 36635
rect 37841 36601 37875 36635
rect 22661 36533 22695 36567
rect 28181 36533 28215 36567
rect 36001 36533 36035 36567
rect 37105 36533 37139 36567
rect 1593 36329 1627 36363
rect 34805 36329 34839 36363
rect 35265 36329 35299 36363
rect 36277 36261 36311 36295
rect 37381 36261 37415 36295
rect 1409 36193 1443 36227
rect 21465 36193 21499 36227
rect 21557 36193 21591 36227
rect 23388 36193 23422 36227
rect 26249 36193 26283 36227
rect 26387 36193 26421 36227
rect 26525 36193 26559 36227
rect 26622 36193 26656 36227
rect 26818 36193 26852 36227
rect 34621 36193 34655 36227
rect 35449 36193 35483 36227
rect 35909 36193 35943 36227
rect 36057 36193 36091 36227
rect 36185 36193 36219 36227
rect 36374 36193 36408 36227
rect 37197 36193 37231 36227
rect 23121 36125 23155 36159
rect 36553 36057 36587 36091
rect 24501 35989 24535 36023
rect 22753 35785 22787 35819
rect 34621 35785 34655 35819
rect 22937 35649 22971 35683
rect 22661 35581 22695 35615
rect 23949 35581 23983 35615
rect 34805 35581 34839 35615
rect 35909 35581 35943 35615
rect 36002 35581 36036 35615
rect 36277 35581 36311 35615
rect 36374 35581 36408 35615
rect 37105 35581 37139 35615
rect 37198 35581 37232 35615
rect 37570 35581 37604 35615
rect 22937 35513 22971 35547
rect 36185 35513 36219 35547
rect 37381 35513 37415 35547
rect 37473 35513 37507 35547
rect 24041 35445 24075 35479
rect 36553 35445 36587 35479
rect 37749 35445 37783 35479
rect 1593 35241 1627 35275
rect 23489 35241 23523 35275
rect 36737 35241 36771 35275
rect 35449 35173 35483 35207
rect 36369 35173 36403 35207
rect 1409 35105 1443 35139
rect 23397 35105 23431 35139
rect 27813 35105 27847 35139
rect 28080 35105 28114 35139
rect 36093 35105 36127 35139
rect 36241 35105 36275 35139
rect 36461 35105 36495 35139
rect 36558 35105 36592 35139
rect 37197 35105 37231 35139
rect 29193 34901 29227 34935
rect 35541 34901 35575 34935
rect 37381 34901 37415 34935
rect 1593 34697 1627 34731
rect 25237 34629 25271 34663
rect 28089 34629 28123 34663
rect 28917 34629 28951 34663
rect 34805 34629 34839 34663
rect 26709 34561 26743 34595
rect 29101 34561 29135 34595
rect 1409 34493 1443 34527
rect 25421 34493 25455 34527
rect 26249 34493 26283 34527
rect 26976 34493 27010 34527
rect 28825 34493 28859 34527
rect 29009 34493 29043 34527
rect 29285 34493 29319 34527
rect 34621 34493 34655 34527
rect 36093 34493 36127 34527
rect 36186 34493 36220 34527
rect 36369 34493 36403 34527
rect 36558 34493 36592 34527
rect 37565 34493 37599 34527
rect 37841 34493 37875 34527
rect 37933 34493 37967 34527
rect 36461 34425 36495 34459
rect 37749 34425 37783 34459
rect 26065 34357 26099 34391
rect 28641 34357 28675 34391
rect 36737 34357 36771 34391
rect 38117 34357 38151 34391
rect 26157 34153 26191 34187
rect 29193 34153 29227 34187
rect 29929 34153 29963 34187
rect 37197 34153 37231 34187
rect 25421 34017 25455 34051
rect 36369 34085 36403 34119
rect 26433 34017 26467 34051
rect 26893 34017 26927 34051
rect 27813 34017 27847 34051
rect 28080 34017 28114 34051
rect 29837 34017 29871 34051
rect 35633 34017 35667 34051
rect 36093 34017 36127 34051
rect 36186 34017 36220 34051
rect 36461 34017 36495 34051
rect 36599 34017 36633 34051
rect 37381 34017 37415 34051
rect 26617 33949 26651 33983
rect 26709 33949 26743 33983
rect 26525 33881 26559 33915
rect 25605 33813 25639 33847
rect 26157 33813 26191 33847
rect 26249 33813 26283 33847
rect 35449 33813 35483 33847
rect 36737 33813 36771 33847
rect 25789 33609 25823 33643
rect 38117 33609 38151 33643
rect 2053 33541 2087 33575
rect 28273 33541 28307 33575
rect 37289 33541 37323 33575
rect 28549 33473 28583 33507
rect 28733 33473 28767 33507
rect 1869 33405 1903 33439
rect 25237 33405 25271 33439
rect 25610 33405 25644 33439
rect 26341 33405 26375 33439
rect 26608 33405 26642 33439
rect 28457 33405 28491 33439
rect 28641 33405 28675 33439
rect 28908 33405 28942 33439
rect 36093 33405 36127 33439
rect 36186 33405 36220 33439
rect 36558 33405 36592 33439
rect 37473 33405 37507 33439
rect 37933 33405 37967 33439
rect 25421 33337 25455 33371
rect 25513 33337 25547 33371
rect 36369 33337 36403 33371
rect 36461 33337 36495 33371
rect 27721 33269 27755 33303
rect 36737 33269 36771 33303
rect 1593 33065 1627 33099
rect 29193 33065 29227 33099
rect 35633 33065 35667 33099
rect 37197 33065 37231 33099
rect 28058 32997 28092 33031
rect 36369 32997 36403 33031
rect 1409 32929 1443 32963
rect 25145 32929 25179 32963
rect 25329 32929 25363 32963
rect 25421 32929 25455 32963
rect 25518 32929 25552 32963
rect 26433 32929 26467 32963
rect 26709 32929 26743 32963
rect 26893 32929 26927 32963
rect 27813 32929 27847 32963
rect 35449 32929 35483 32963
rect 36093 32929 36127 32963
rect 36241 32929 36275 32963
rect 36461 32929 36495 32963
rect 36558 32929 36592 32963
rect 37381 32929 37415 32963
rect 26617 32861 26651 32895
rect 25697 32793 25731 32827
rect 26525 32793 26559 32827
rect 36737 32793 36771 32827
rect 26249 32725 26283 32759
rect 25973 32521 26007 32555
rect 28181 32521 28215 32555
rect 36277 32521 36311 32555
rect 37105 32521 37139 32555
rect 23857 32453 23891 32487
rect 26893 32385 26927 32419
rect 26985 32385 27019 32419
rect 25421 32317 25455 32351
rect 25794 32317 25828 32351
rect 26709 32317 26743 32351
rect 26801 32317 26835 32351
rect 27169 32317 27203 32351
rect 27629 32317 27663 32351
rect 27813 32317 27847 32351
rect 28002 32317 28036 32351
rect 36093 32317 36127 32351
rect 36921 32317 36955 32351
rect 37565 32317 37599 32351
rect 37933 32317 37967 32351
rect 23673 32249 23707 32283
rect 25605 32249 25639 32283
rect 25697 32249 25731 32283
rect 27905 32249 27939 32283
rect 37749 32249 37783 32283
rect 37841 32249 37875 32283
rect 26525 32181 26559 32215
rect 38117 32181 38151 32215
rect 1593 31977 1627 32011
rect 28373 31977 28407 32011
rect 35725 31977 35759 32011
rect 36369 31977 36403 32011
rect 24777 31909 24811 31943
rect 26249 31909 26283 31943
rect 27997 31909 28031 31943
rect 28089 31909 28123 31943
rect 37013 31909 37047 31943
rect 37105 31909 37139 31943
rect 1409 31841 1443 31875
rect 22569 31841 22603 31875
rect 22661 31841 22695 31875
rect 24869 31841 24903 31875
rect 25053 31841 25087 31875
rect 25145 31841 25179 31875
rect 25242 31841 25276 31875
rect 25973 31841 26007 31875
rect 26157 31841 26191 31875
rect 26393 31841 26427 31875
rect 27813 31841 27847 31875
rect 28186 31841 28220 31875
rect 35541 31841 35575 31875
rect 36185 31841 36219 31875
rect 36829 31841 36863 31875
rect 37197 31841 37231 31875
rect 25421 31705 25455 31739
rect 26525 31705 26559 31739
rect 24777 31637 24811 31671
rect 37381 31637 37415 31671
rect 1593 31433 1627 31467
rect 27629 31433 27663 31467
rect 28365 31433 28399 31467
rect 26249 31365 26283 31399
rect 26341 31297 26375 31331
rect 26433 31297 26467 31331
rect 1409 31229 1443 31263
rect 26157 31229 26191 31263
rect 26617 31229 26651 31263
rect 27077 31229 27111 31263
rect 27497 31229 27531 31263
rect 28181 31229 28215 31263
rect 36553 31229 36587 31263
rect 36921 31229 36955 31263
rect 37565 31229 37599 31263
rect 37841 31229 37875 31263
rect 37933 31229 37967 31263
rect 25329 31161 25363 31195
rect 27261 31161 27295 31195
rect 27353 31161 27387 31195
rect 36737 31161 36771 31195
rect 36829 31161 36863 31195
rect 37749 31161 37783 31195
rect 25421 31093 25455 31127
rect 25973 31093 26007 31127
rect 37105 31093 37139 31127
rect 38117 31093 38151 31127
rect 36093 30889 36127 30923
rect 36553 30889 36587 30923
rect 37381 30889 37415 30923
rect 25596 30821 25630 30855
rect 27813 30753 27847 30787
rect 35909 30753 35943 30787
rect 36737 30753 36771 30787
rect 37197 30753 37231 30787
rect 25329 30685 25363 30719
rect 26709 30549 26743 30583
rect 27997 30549 28031 30583
rect 35909 30345 35943 30379
rect 36645 30345 36679 30379
rect 1593 30277 1627 30311
rect 26617 30277 26651 30311
rect 27169 30209 27203 30243
rect 1409 30141 1443 30175
rect 25237 30141 25271 30175
rect 27436 30141 27470 30175
rect 36001 30141 36035 30175
rect 36094 30141 36128 30175
rect 36231 30141 36265 30175
rect 36369 30141 36403 30175
rect 36466 30141 36500 30175
rect 37565 30141 37599 30175
rect 37841 30141 37875 30175
rect 37933 30141 37967 30175
rect 25504 30073 25538 30107
rect 35909 30073 35943 30107
rect 37749 30073 37783 30107
rect 28549 30005 28583 30039
rect 38117 30005 38151 30039
rect 19441 29801 19475 29835
rect 37197 29801 37231 29835
rect 19165 29733 19199 29767
rect 24584 29733 24618 29767
rect 36369 29733 36403 29767
rect 18797 29665 18831 29699
rect 18945 29665 18979 29699
rect 19073 29665 19107 29699
rect 19262 29665 19296 29699
rect 22753 29665 22787 29699
rect 22937 29665 22971 29699
rect 23213 29665 23247 29699
rect 24317 29665 24351 29699
rect 26433 29665 26467 29699
rect 26709 29665 26743 29699
rect 26893 29665 26927 29699
rect 35357 29665 35391 29699
rect 36001 29665 36035 29699
rect 36149 29665 36183 29699
rect 36277 29665 36311 29699
rect 36466 29665 36500 29699
rect 37381 29665 37415 29699
rect 23029 29597 23063 29631
rect 26525 29597 26559 29631
rect 26617 29597 26651 29631
rect 22845 29529 22879 29563
rect 25697 29529 25731 29563
rect 36645 29529 36679 29563
rect 22569 29461 22603 29495
rect 26249 29461 26283 29495
rect 35541 29461 35575 29495
rect 1593 29257 1627 29291
rect 37289 29257 37323 29291
rect 37933 29257 37967 29291
rect 27721 29189 27755 29223
rect 23581 29121 23615 29155
rect 24041 29121 24075 29155
rect 27445 29121 27479 29155
rect 27922 29121 27956 29155
rect 1409 29053 1443 29087
rect 18436 29053 18470 29087
rect 18522 29053 18556 29087
rect 18894 29053 18928 29087
rect 22385 29053 22419 29087
rect 22477 29053 22511 29087
rect 22661 29053 22695 29087
rect 23765 29053 23799 29087
rect 23857 29053 23891 29087
rect 23949 29053 23983 29087
rect 24225 29053 24259 29087
rect 27629 29053 27663 29087
rect 27813 29053 27847 29087
rect 28101 29053 28135 29087
rect 35909 29053 35943 29087
rect 36002 29053 36036 29087
rect 36374 29053 36408 29087
rect 37473 29053 37507 29087
rect 38117 29053 38151 29087
rect 18705 28985 18739 29019
rect 18797 28985 18831 29019
rect 25237 28985 25271 29019
rect 26985 28985 27019 29019
rect 36185 28985 36219 29019
rect 36277 28985 36311 29019
rect 19073 28917 19107 28951
rect 22845 28917 22879 28951
rect 36553 28917 36587 28951
rect 19349 28713 19383 28747
rect 20453 28713 20487 28747
rect 37381 28713 37415 28747
rect 18981 28645 19015 28679
rect 20085 28645 20119 28679
rect 36277 28645 36311 28679
rect 1685 28577 1719 28611
rect 18694 28577 18728 28611
rect 18798 28577 18832 28611
rect 19073 28577 19107 28611
rect 19170 28577 19204 28611
rect 19809 28577 19843 28611
rect 19957 28577 19991 28611
rect 20177 28577 20211 28611
rect 20274 28577 20308 28611
rect 22569 28577 22603 28611
rect 22825 28577 22859 28611
rect 25237 28577 25271 28611
rect 25504 28577 25538 28611
rect 35909 28577 35943 28611
rect 36002 28577 36036 28611
rect 36185 28577 36219 28611
rect 36415 28577 36449 28611
rect 37197 28577 37231 28611
rect 1409 28509 1443 28543
rect 23949 28373 23983 28407
rect 26617 28373 26651 28407
rect 36553 28373 36587 28407
rect 19073 28169 19107 28203
rect 37289 28169 37323 28203
rect 38117 28169 38151 28203
rect 27169 28101 27203 28135
rect 36553 28101 36587 28135
rect 26157 28033 26191 28067
rect 26249 28033 26283 28067
rect 18429 27965 18463 27999
rect 18577 27965 18611 27999
rect 18935 27965 18969 27999
rect 21005 27965 21039 27999
rect 22845 27965 22879 27999
rect 25973 27965 26007 27999
rect 26065 27965 26099 27999
rect 26433 27965 26467 27999
rect 27077 27965 27111 27999
rect 27261 27965 27295 27999
rect 27370 27965 27404 27999
rect 27537 27965 27571 27999
rect 35909 27965 35943 27999
rect 36002 27965 36036 27999
rect 36277 27965 36311 27999
rect 36374 27965 36408 27999
rect 37473 27965 37507 27999
rect 37933 27965 37967 27999
rect 18705 27897 18739 27931
rect 18797 27897 18831 27931
rect 21272 27897 21306 27931
rect 23112 27897 23146 27931
rect 36185 27897 36219 27931
rect 22385 27829 22419 27863
rect 24225 27829 24259 27863
rect 25789 27829 25823 27863
rect 26893 27829 26927 27863
rect 19809 27625 19843 27659
rect 36185 27625 36219 27659
rect 1869 27557 1903 27591
rect 2053 27557 2087 27591
rect 20536 27557 20570 27591
rect 22814 27557 22848 27591
rect 24409 27557 24443 27591
rect 19441 27489 19475 27523
rect 24748 27489 24782 27523
rect 25789 27489 25823 27523
rect 25973 27489 26007 27523
rect 26065 27489 26099 27523
rect 26249 27489 26283 27523
rect 26709 27489 26743 27523
rect 36001 27489 36035 27523
rect 19533 27421 19567 27455
rect 20269 27421 20303 27455
rect 22569 27421 22603 27455
rect 25605 27353 25639 27387
rect 25881 27353 25915 27387
rect 19625 27285 19659 27319
rect 21649 27285 21683 27319
rect 23949 27285 23983 27319
rect 24547 27285 24581 27319
rect 24685 27285 24719 27319
rect 25053 27285 25087 27319
rect 26893 27285 26927 27319
rect 37473 27081 37507 27115
rect 38117 27081 38151 27115
rect 2053 27013 2087 27047
rect 21373 27013 21407 27047
rect 19993 26945 20027 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 21833 26877 21867 26911
rect 22100 26877 22134 26911
rect 25421 26877 25455 26911
rect 25513 26877 25547 26911
rect 25881 26877 25915 26911
rect 37289 26877 37323 26911
rect 37933 26877 37967 26911
rect 1869 26809 1903 26843
rect 20260 26809 20294 26843
rect 24133 26809 24167 26843
rect 23213 26741 23247 26775
rect 24225 26741 24259 26775
rect 25237 26741 25271 26775
rect 20085 26537 20119 26571
rect 21281 26537 21315 26571
rect 20637 26469 20671 26503
rect 23480 26469 23514 26503
rect 18521 26401 18555 26435
rect 18961 26401 18995 26435
rect 25412 26401 25446 26435
rect 18705 26333 18739 26367
rect 21005 26333 21039 26367
rect 23213 26333 23247 26367
rect 25145 26333 25179 26367
rect 20802 26265 20836 26299
rect 24593 26265 24627 26299
rect 26525 26265 26559 26299
rect 20913 26197 20947 26231
rect 18705 25993 18739 26027
rect 22293 25993 22327 26027
rect 24225 25993 24259 26027
rect 26617 25993 26651 26027
rect 38117 25993 38151 26027
rect 2053 25925 2087 25959
rect 37473 25925 37507 25959
rect 20913 25857 20947 25891
rect 25237 25857 25271 25891
rect 1869 25789 1903 25823
rect 18061 25789 18095 25823
rect 18154 25789 18188 25823
rect 18526 25789 18560 25823
rect 21180 25789 21214 25823
rect 22845 25789 22879 25823
rect 25504 25789 25538 25823
rect 37289 25789 37323 25823
rect 37933 25789 37967 25823
rect 18337 25721 18371 25755
rect 18429 25721 18463 25755
rect 23112 25721 23146 25755
rect 18521 25449 18555 25483
rect 23949 25449 23983 25483
rect 37381 25449 37415 25483
rect 2053 25381 2087 25415
rect 18245 25381 18279 25415
rect 19248 25381 19282 25415
rect 22836 25381 22870 25415
rect 1869 25313 1903 25347
rect 17877 25313 17911 25347
rect 18025 25313 18059 25347
rect 18153 25313 18187 25347
rect 18342 25313 18376 25347
rect 18981 25313 19015 25347
rect 21373 25313 21407 25347
rect 24961 25313 24995 25347
rect 25145 25313 25179 25347
rect 25237 25313 25271 25347
rect 25421 25313 25455 25347
rect 26065 25313 26099 25347
rect 26341 25313 26375 25347
rect 26525 25313 26559 25347
rect 37197 25313 37231 25347
rect 22569 25245 22603 25279
rect 26249 25245 26283 25279
rect 21557 25177 21591 25211
rect 25053 25177 25087 25211
rect 26157 25177 26191 25211
rect 20361 25109 20395 25143
rect 24777 25109 24811 25143
rect 25881 25109 25915 25143
rect 23949 24837 23983 24871
rect 25513 24837 25547 24871
rect 23673 24769 23707 24803
rect 24050 24769 24084 24803
rect 16865 24701 16899 24735
rect 17013 24701 17047 24735
rect 17330 24701 17364 24735
rect 17969 24701 18003 24735
rect 18062 24701 18096 24735
rect 18434 24701 18468 24735
rect 20269 24701 20303 24735
rect 21097 24701 21131 24735
rect 21189 24701 21223 24735
rect 21373 24701 21407 24735
rect 23857 24701 23891 24735
rect 24133 24701 24167 24735
rect 24317 24701 24351 24735
rect 25421 24701 25455 24735
rect 25605 24701 25639 24735
rect 25697 24701 25731 24735
rect 25881 24701 25915 24735
rect 37933 24701 37967 24735
rect 17141 24633 17175 24667
rect 17233 24633 17267 24667
rect 18245 24633 18279 24667
rect 18337 24633 18371 24667
rect 20085 24633 20119 24667
rect 21925 24633 21959 24667
rect 22661 24633 22695 24667
rect 17509 24565 17543 24599
rect 18613 24565 18647 24599
rect 22017 24565 22051 24599
rect 22753 24565 22787 24599
rect 25237 24565 25271 24599
rect 38117 24565 38151 24599
rect 21557 24361 21591 24395
rect 37381 24361 37415 24395
rect 1869 24293 1903 24327
rect 2053 24293 2087 24327
rect 17877 24293 17911 24327
rect 18880 24293 18914 24327
rect 17509 24225 17543 24259
rect 17602 24225 17636 24259
rect 17785 24225 17819 24259
rect 17974 24225 18008 24259
rect 18613 24225 18647 24259
rect 21465 24225 21499 24259
rect 24685 24225 24719 24259
rect 37197 24225 37231 24259
rect 24501 24089 24535 24123
rect 18153 24021 18187 24055
rect 19993 24021 20027 24055
rect 37289 23817 37323 23851
rect 37933 23817 37967 23851
rect 2053 23749 2087 23783
rect 18705 23749 18739 23783
rect 1869 23613 1903 23647
rect 18521 23613 18555 23647
rect 19993 23613 20027 23647
rect 21373 23613 21407 23647
rect 21557 23613 21591 23647
rect 22201 23613 22235 23647
rect 37473 23613 37507 23647
rect 38117 23613 38151 23647
rect 20085 23477 20119 23511
rect 22017 23477 22051 23511
rect 17693 23273 17727 23307
rect 18337 23273 18371 23307
rect 20177 23273 20211 23307
rect 23949 23273 23983 23307
rect 37381 23273 37415 23307
rect 19064 23205 19098 23239
rect 22836 23205 22870 23239
rect 17509 23137 17543 23171
rect 18153 23137 18187 23171
rect 21189 23137 21223 23171
rect 37197 23137 37231 23171
rect 18797 23069 18831 23103
rect 22569 23069 22603 23103
rect 21281 22933 21315 22967
rect 1593 22729 1627 22763
rect 22753 22729 22787 22763
rect 37473 22729 37507 22763
rect 38117 22729 38151 22763
rect 18613 22661 18647 22695
rect 23857 22661 23891 22695
rect 23958 22593 23992 22627
rect 1409 22525 1443 22559
rect 17969 22525 18003 22559
rect 18117 22525 18151 22559
rect 18245 22525 18279 22559
rect 18337 22525 18371 22559
rect 18434 22525 18468 22559
rect 21373 22525 21407 22559
rect 21640 22525 21674 22559
rect 23765 22525 23799 22559
rect 24058 22525 24092 22559
rect 24225 22525 24259 22559
rect 37289 22525 37323 22559
rect 37933 22525 37967 22559
rect 23581 22389 23615 22423
rect 18889 22117 18923 22151
rect 18981 22117 19015 22151
rect 1409 22049 1443 22083
rect 17785 22049 17819 22083
rect 18602 22049 18636 22083
rect 18733 22049 18767 22083
rect 19078 22049 19112 22083
rect 20177 22049 20211 22083
rect 20444 22049 20478 22083
rect 22569 22049 22603 22083
rect 22836 22049 22870 22083
rect 24685 22049 24719 22083
rect 24869 22049 24903 22083
rect 25145 22049 25179 22083
rect 37197 22049 37231 22083
rect 17417 21981 17451 22015
rect 17969 21981 18003 22015
rect 24961 21981 24995 22015
rect 1593 21913 1627 21947
rect 19257 21913 19291 21947
rect 24777 21913 24811 21947
rect 21557 21845 21591 21879
rect 23949 21845 23983 21879
rect 24501 21845 24535 21879
rect 37381 21845 37415 21879
rect 18521 21641 18555 21675
rect 20269 21641 20303 21675
rect 22201 21641 22235 21675
rect 37473 21641 37507 21675
rect 38117 21573 38151 21607
rect 20821 21505 20855 21539
rect 22753 21505 22787 21539
rect 16773 21437 16807 21471
rect 16921 21437 16955 21471
rect 17141 21437 17175 21471
rect 17238 21437 17272 21471
rect 17866 21437 17900 21471
rect 18025 21437 18059 21471
rect 18153 21437 18187 21471
rect 18342 21437 18376 21471
rect 21088 21437 21122 21471
rect 23020 21437 23054 21471
rect 37289 21437 37323 21471
rect 37933 21437 37967 21471
rect 17049 21369 17083 21403
rect 18245 21369 18279 21403
rect 20177 21369 20211 21403
rect 17417 21301 17451 21335
rect 24133 21301 24167 21335
rect 1593 21097 1627 21131
rect 18061 21029 18095 21063
rect 18153 21029 18187 21063
rect 20821 21029 20855 21063
rect 1409 20961 1443 20995
rect 17785 20961 17819 20995
rect 17878 20961 17912 20995
rect 18250 20961 18284 20995
rect 23489 20961 23523 20995
rect 23673 20961 23707 20995
rect 23949 20961 23983 20995
rect 24593 20961 24627 20995
rect 24777 20961 24811 20995
rect 25053 20961 25087 20995
rect 23765 20893 23799 20927
rect 24869 20893 24903 20927
rect 18429 20825 18463 20859
rect 23581 20825 23615 20859
rect 24685 20825 24719 20859
rect 20913 20757 20947 20791
rect 23305 20757 23339 20791
rect 24409 20757 24443 20791
rect 1593 20553 1627 20587
rect 38117 20553 38151 20587
rect 23397 20485 23431 20519
rect 23489 20417 23523 20451
rect 1409 20349 1443 20383
rect 23305 20349 23339 20383
rect 23581 20349 23615 20383
rect 23765 20349 23799 20383
rect 37289 20349 37323 20383
rect 37933 20349 37967 20383
rect 23121 20213 23155 20247
rect 37473 20213 37507 20247
rect 17601 19941 17635 19975
rect 17693 19941 17727 19975
rect 17325 19873 17359 19907
rect 17418 19873 17452 19907
rect 17790 19873 17824 19907
rect 17969 19669 18003 19703
rect 1409 19261 1443 19295
rect 16037 19261 16071 19295
rect 16129 19261 16163 19295
rect 16249 19261 16283 19295
rect 16405 19261 16439 19295
rect 16497 19261 16531 19295
rect 16594 19261 16628 19295
rect 17233 19261 17267 19295
rect 17326 19261 17360 19295
rect 17509 19261 17543 19295
rect 17698 19261 17732 19295
rect 19993 19261 20027 19295
rect 21925 19261 21959 19295
rect 22192 19261 22226 19295
rect 37289 19261 37323 19295
rect 37933 19261 37967 19295
rect 17601 19193 17635 19227
rect 20260 19193 20294 19227
rect 1593 19125 1627 19159
rect 16037 19125 16071 19159
rect 16773 19125 16807 19159
rect 17877 19125 17911 19159
rect 21373 19125 21407 19159
rect 23305 19125 23339 19159
rect 37473 19125 37507 19159
rect 38117 19125 38151 19159
rect 1593 18921 1627 18955
rect 19073 18921 19107 18955
rect 37381 18921 37415 18955
rect 16129 18853 16163 18887
rect 18705 18853 18739 18887
rect 18797 18853 18831 18887
rect 1409 18785 1443 18819
rect 15761 18785 15795 18819
rect 15909 18785 15943 18819
rect 16037 18785 16071 18819
rect 16267 18785 16301 18819
rect 17325 18785 17359 18819
rect 17418 18785 17452 18819
rect 17601 18785 17635 18819
rect 17701 18785 17735 18819
rect 17831 18785 17865 18819
rect 18429 18785 18463 18819
rect 18522 18785 18556 18819
rect 18894 18785 18928 18819
rect 19533 18785 19567 18819
rect 19800 18785 19834 18819
rect 37197 18785 37231 18819
rect 16405 18581 16439 18615
rect 17969 18581 18003 18615
rect 20913 18581 20947 18615
rect 18797 18377 18831 18411
rect 38117 18377 38151 18411
rect 19993 18241 20027 18275
rect 16589 18173 16623 18207
rect 16737 18173 16771 18207
rect 16865 18173 16899 18207
rect 16957 18173 16991 18207
rect 17054 18173 17088 18207
rect 17969 18173 18003 18207
rect 18889 18173 18923 18207
rect 20260 18173 20294 18207
rect 37933 18173 37967 18207
rect 17233 18037 17267 18071
rect 21373 18037 21407 18071
rect 1593 17833 1627 17867
rect 17969 17833 18003 17867
rect 37381 17833 37415 17867
rect 17601 17765 17635 17799
rect 17693 17765 17727 17799
rect 1409 17697 1443 17731
rect 17325 17697 17359 17731
rect 17473 17697 17507 17731
rect 17790 17697 17824 17731
rect 19809 17697 19843 17731
rect 20076 17697 20110 17731
rect 37197 17697 37231 17731
rect 21189 17493 21223 17527
rect 1593 17289 1627 17323
rect 21281 17289 21315 17323
rect 37473 17289 37507 17323
rect 38117 17221 38151 17255
rect 1409 17085 1443 17119
rect 21465 17085 21499 17119
rect 21557 17085 21591 17119
rect 21767 17085 21801 17119
rect 21925 17085 21959 17119
rect 37289 17085 37323 17119
rect 37933 17085 37967 17119
rect 21649 17017 21683 17051
rect 37289 16745 37323 16779
rect 37197 16609 37231 16643
rect 1593 16201 1627 16235
rect 37473 16201 37507 16235
rect 17233 16133 17267 16167
rect 38117 16133 38151 16167
rect 1409 15997 1443 16031
rect 16589 15997 16623 16031
rect 16737 15997 16771 16031
rect 17054 15997 17088 16031
rect 37289 15997 37323 16031
rect 37933 15997 37967 16031
rect 16865 15929 16899 15963
rect 16957 15929 16991 15963
rect 1593 15657 1627 15691
rect 17969 15657 18003 15691
rect 37289 15657 37323 15691
rect 17693 15589 17727 15623
rect 1409 15521 1443 15555
rect 15761 15521 15795 15555
rect 15854 15521 15888 15555
rect 16037 15521 16071 15555
rect 16129 15521 16163 15555
rect 16226 15521 16260 15555
rect 17325 15521 17359 15555
rect 17473 15521 17507 15555
rect 17601 15521 17635 15555
rect 17790 15521 17824 15555
rect 37197 15521 37231 15555
rect 16405 15385 16439 15419
rect 17141 15113 17175 15147
rect 18245 15113 18279 15147
rect 37473 15113 37507 15147
rect 38117 15045 38151 15079
rect 16497 14909 16531 14943
rect 16590 14909 16624 14943
rect 16773 14909 16807 14943
rect 17003 14909 17037 14943
rect 17601 14909 17635 14943
rect 17694 14909 17728 14943
rect 17877 14909 17911 14943
rect 18066 14909 18100 14943
rect 37289 14909 37323 14943
rect 37933 14909 37967 14943
rect 16865 14841 16899 14875
rect 17969 14841 18003 14875
rect 1593 14569 1627 14603
rect 1409 14433 1443 14467
rect 29009 14433 29043 14467
rect 29193 14229 29227 14263
rect 1593 14025 1627 14059
rect 37289 14025 37323 14059
rect 38117 13957 38151 13991
rect 1409 13821 1443 13855
rect 37197 13821 37231 13855
rect 37933 13821 37967 13855
rect 37197 13345 37231 13379
rect 37289 13141 37323 13175
rect 1593 12937 1627 12971
rect 38025 12937 38059 12971
rect 21005 12801 21039 12835
rect 1409 12733 1443 12767
rect 21373 12733 21407 12767
rect 21465 12665 21499 12699
rect 21741 12665 21775 12699
rect 37933 12665 37967 12699
rect 21281 12597 21315 12631
rect 1593 12393 1627 12427
rect 37289 12393 37323 12427
rect 1409 12257 1443 12291
rect 37197 12257 37231 12291
rect 38025 11849 38059 11883
rect 37197 11645 37231 11679
rect 37933 11577 37967 11611
rect 37289 11509 37323 11543
rect 1409 11169 1443 11203
rect 37197 11169 37231 11203
rect 1593 11033 1627 11067
rect 37381 11033 37415 11067
rect 37933 10489 37967 10523
rect 38025 10421 38059 10455
rect 1409 10081 1443 10115
rect 37197 10081 37231 10115
rect 1593 9877 1627 9911
rect 37289 9877 37323 9911
rect 37381 9605 37415 9639
rect 38117 9605 38151 9639
rect 1409 9469 1443 9503
rect 37197 9469 37231 9503
rect 37933 9401 37967 9435
rect 1593 9333 1627 9367
rect 37289 9129 37323 9163
rect 23397 9061 23431 9095
rect 22661 8993 22695 9027
rect 22845 8993 22879 9027
rect 23029 8993 23063 9027
rect 23305 8993 23339 9027
rect 37197 8993 37231 9027
rect 1409 8381 1443 8415
rect 38117 8381 38151 8415
rect 37933 8313 37967 8347
rect 1593 8245 1627 8279
rect 1593 8041 1627 8075
rect 1409 7905 1443 7939
rect 37197 7905 37231 7939
rect 37289 7701 37323 7735
rect 17141 7497 17175 7531
rect 38025 7497 38059 7531
rect 16865 7293 16899 7327
rect 37197 7293 37231 7327
rect 37933 7225 37967 7259
rect 37289 7157 37323 7191
rect 1409 6817 1443 6851
rect 37197 6817 37231 6851
rect 37381 6817 37415 6851
rect 1593 6681 1627 6715
rect 1593 6409 1627 6443
rect 37289 6409 37323 6443
rect 38117 6341 38151 6375
rect 1409 6205 1443 6239
rect 36461 6137 36495 6171
rect 36645 6137 36679 6171
rect 37197 6137 37231 6171
rect 37933 6137 37967 6171
rect 1593 5865 1627 5899
rect 35357 5797 35391 5831
rect 1409 5729 1443 5763
rect 2881 5729 2915 5763
rect 36093 5729 36127 5763
rect 37197 5729 37231 5763
rect 37381 5593 37415 5627
rect 2697 5525 2731 5559
rect 35449 5525 35483 5559
rect 36185 5525 36219 5559
rect 1593 5321 1627 5355
rect 2237 5321 2271 5355
rect 2973 5321 3007 5355
rect 36553 5321 36587 5355
rect 38025 5321 38059 5355
rect 37381 5253 37415 5287
rect 1409 5117 1443 5151
rect 2053 5117 2087 5151
rect 2789 5117 2823 5151
rect 31493 5117 31527 5151
rect 34069 5117 34103 5151
rect 37197 5117 37231 5151
rect 33885 5049 33919 5083
rect 34621 5049 34655 5083
rect 36461 5049 36495 5083
rect 37933 5049 37967 5083
rect 31309 4981 31343 5015
rect 34713 4981 34747 5015
rect 36553 4777 36587 4811
rect 34253 4709 34287 4743
rect 34989 4709 35023 4743
rect 35909 4709 35943 4743
rect 37381 4709 37415 4743
rect 1869 4641 1903 4675
rect 3341 4641 3375 4675
rect 14657 4641 14691 4675
rect 22753 4641 22787 4675
rect 23397 4641 23431 4675
rect 25421 4641 25455 4675
rect 26801 4641 26835 4675
rect 30297 4641 30331 4675
rect 30757 4641 30791 4675
rect 31585 4641 31619 4675
rect 33517 4641 33551 4675
rect 35725 4641 35759 4675
rect 36461 4641 36495 4675
rect 37197 4641 37231 4675
rect 33701 4573 33735 4607
rect 23213 4505 23247 4539
rect 30941 4505 30975 4539
rect 34437 4505 34471 4539
rect 1961 4437 1995 4471
rect 2697 4437 2731 4471
rect 14841 4437 14875 4471
rect 22569 4437 22603 4471
rect 25237 4437 25271 4471
rect 26617 4437 26651 4471
rect 30113 4437 30147 4471
rect 31401 4437 31435 4471
rect 35081 4437 35115 4471
rect 10241 4233 10275 4267
rect 4261 4165 4295 4199
rect 23949 4165 23983 4199
rect 26801 4165 26835 4199
rect 28549 4165 28583 4199
rect 34713 4165 34747 4199
rect 9873 4097 9907 4131
rect 36645 4097 36679 4131
rect 37381 4097 37415 4131
rect 38117 4097 38151 4131
rect 1869 4029 1903 4063
rect 2605 4029 2639 4063
rect 4445 4029 4479 4063
rect 4905 4029 4939 4063
rect 5549 4029 5583 4063
rect 6193 4029 6227 4063
rect 7113 4029 7147 4063
rect 10977 4029 11011 4063
rect 11713 4029 11747 4063
rect 15025 4029 15059 4063
rect 15945 4029 15979 4063
rect 18061 4029 18095 4063
rect 20177 4029 20211 4063
rect 20821 4029 20855 4063
rect 21557 4029 21591 4063
rect 22017 4029 22051 4063
rect 22661 4029 22695 4063
rect 23305 4029 23339 4063
rect 24133 4029 24167 4063
rect 25421 4029 25455 4063
rect 26065 4029 26099 4063
rect 26617 4029 26651 4063
rect 27261 4029 27295 4063
rect 28089 4029 28123 4063
rect 28733 4029 28767 4063
rect 29469 4029 29503 4063
rect 30849 4029 30883 4063
rect 32505 4029 32539 4063
rect 33885 4029 33919 4063
rect 34529 4029 34563 4063
rect 35909 4029 35943 4063
rect 2789 3961 2823 3995
rect 31677 3961 31711 3995
rect 33149 3961 33183 3995
rect 36461 3961 36495 3995
rect 37197 3961 37231 3995
rect 37933 3961 37967 3995
rect 1961 3893 1995 3927
rect 10241 3893 10275 3927
rect 10425 3893 10459 3927
rect 11069 3893 11103 3927
rect 11805 3893 11839 3927
rect 15117 3893 15151 3927
rect 16037 3893 16071 3927
rect 17877 3893 17911 3927
rect 19993 3893 20027 3927
rect 20637 3893 20671 3927
rect 21373 3893 21407 3927
rect 22201 3893 22235 3927
rect 22845 3893 22879 3927
rect 23489 3893 23523 3927
rect 25237 3893 25271 3927
rect 25881 3893 25915 3927
rect 27353 3893 27387 3927
rect 27905 3893 27939 3927
rect 29285 3893 29319 3927
rect 30941 3893 30975 3927
rect 31769 3893 31803 3927
rect 32321 3893 32355 3927
rect 33241 3893 33275 3927
rect 33977 3893 34011 3927
rect 35725 3893 35759 3927
rect 1961 3689 1995 3723
rect 3433 3689 3467 3723
rect 7757 3689 7791 3723
rect 8769 3689 8803 3723
rect 11069 3689 11103 3723
rect 12265 3689 12299 3723
rect 16313 3689 16347 3723
rect 22017 3689 22051 3723
rect 26249 3689 26283 3723
rect 27169 3689 27203 3723
rect 33517 3689 33551 3723
rect 34253 3689 34287 3723
rect 34989 3689 35023 3723
rect 35909 3689 35943 3723
rect 37289 3689 37323 3723
rect 1869 3621 1903 3655
rect 4077 3621 4111 3655
rect 6929 3621 6963 3655
rect 9413 3621 9447 3655
rect 10149 3621 10183 3655
rect 12909 3621 12943 3655
rect 14105 3621 14139 3655
rect 17417 3621 17451 3655
rect 18153 3621 18187 3655
rect 2605 3553 2639 3587
rect 3249 3553 3283 3587
rect 4997 3553 5031 3587
rect 5641 3553 5675 3587
rect 7573 3553 7607 3587
rect 8585 3553 8619 3587
rect 10885 3553 10919 3587
rect 12081 3553 12115 3587
rect 13829 3553 13863 3587
rect 14841 3553 14875 3587
rect 15485 3553 15519 3587
rect 16129 3553 16163 3587
rect 18889 3553 18923 3587
rect 19717 3553 19751 3587
rect 20361 3553 20395 3587
rect 21005 3553 21039 3587
rect 2789 3485 2823 3519
rect 5825 3417 5859 3451
rect 15669 3417 15703 3451
rect 20545 3417 20579 3451
rect 21189 3417 21223 3451
rect 23857 3621 23891 3655
rect 25421 3621 25455 3655
rect 22937 3553 22971 3587
rect 24685 3553 24719 3587
rect 26065 3553 26099 3587
rect 28181 3621 28215 3655
rect 28917 3621 28951 3655
rect 30481 3621 30515 3655
rect 31033 3621 31067 3655
rect 29561 3553 29595 3587
rect 30083 3553 30117 3587
rect 31217 3553 31251 3587
rect 31953 3553 31987 3587
rect 33333 3553 33367 3587
rect 34069 3553 34103 3587
rect 34805 3553 34839 3587
rect 35725 3553 35759 3587
rect 37197 3553 37231 3587
rect 27169 3417 27203 3451
rect 30021 3417 30055 3451
rect 32137 3417 32171 3451
rect 4169 3349 4203 3383
rect 5181 3349 5215 3383
rect 7021 3349 7055 3383
rect 9505 3349 9539 3383
rect 10241 3349 10275 3383
rect 13001 3349 13035 3383
rect 14933 3349 14967 3383
rect 17509 3349 17543 3383
rect 18245 3349 18279 3383
rect 18981 3349 19015 3383
rect 19533 3349 19567 3383
rect 22017 3349 22051 3383
rect 23029 3349 23063 3383
rect 23949 3349 23983 3383
rect 24501 3349 24535 3383
rect 25513 3349 25547 3383
rect 28273 3349 28307 3383
rect 29009 3349 29043 3383
rect 29929 3349 29963 3383
rect 1961 3145 1995 3179
rect 4445 3145 4479 3179
rect 7849 3145 7883 3179
rect 8585 3145 8619 3179
rect 11069 3145 11103 3179
rect 17601 3145 17635 3179
rect 18705 3145 18739 3179
rect 21005 3145 21039 3179
rect 23562 3145 23596 3179
rect 26322 3145 26356 3179
rect 29469 3145 29503 3179
rect 32413 3145 32447 3179
rect 33149 3145 33183 3179
rect 33885 3145 33919 3179
rect 38025 3145 38059 3179
rect 17490 3077 17524 3111
rect 23673 3077 23707 3111
rect 26433 3077 26467 3111
rect 26801 3077 26835 3111
rect 31033 3077 31067 3111
rect 3157 3009 3191 3043
rect 6745 3009 6779 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 15761 3009 15795 3043
rect 17693 3009 17727 3043
rect 23765 3009 23799 3043
rect 26525 3009 26559 3043
rect 31769 3009 31803 3043
rect 36001 3009 36035 3043
rect 37381 3009 37415 3043
rect 2881 2941 2915 2975
rect 4261 2941 4295 2975
rect 5089 2941 5123 2975
rect 5825 2941 5859 2975
rect 6469 2941 6503 2975
rect 7665 2941 7699 2975
rect 8401 2941 8435 2975
rect 10241 2941 10275 2975
rect 10885 2941 10919 2975
rect 11805 2941 11839 2975
rect 12909 2941 12943 2975
rect 15577 2941 15611 2975
rect 16589 2941 16623 2975
rect 17325 2941 17359 2975
rect 18521 2941 18555 2975
rect 20085 2941 20119 2975
rect 20821 2941 20855 2975
rect 21649 2941 21683 2975
rect 23397 2941 23431 2975
rect 25329 2941 25363 2975
rect 26157 2941 26191 2975
rect 27445 2941 27479 2975
rect 28181 2941 28215 2975
rect 29285 2941 29319 2975
rect 30849 2941 30883 2975
rect 32229 2941 32263 2975
rect 32965 2941 32999 2975
rect 33701 2941 33735 2975
rect 34437 2941 34471 2975
rect 35725 2941 35759 2975
rect 1869 2873 1903 2907
rect 9597 2873 9631 2907
rect 14841 2873 14875 2907
rect 18061 2873 18095 2907
rect 22385 2873 22419 2907
rect 27629 2873 27663 2907
rect 31585 2873 31619 2907
rect 37197 2873 37231 2907
rect 37933 2873 37967 2907
rect 5181 2805 5215 2839
rect 5917 2805 5951 2839
rect 9689 2805 9723 2839
rect 10425 2805 10459 2839
rect 14933 2805 14967 2839
rect 16773 2805 16807 2839
rect 20177 2805 20211 2839
rect 21741 2805 21775 2839
rect 22477 2805 22511 2839
rect 24041 2805 24075 2839
rect 25421 2805 25455 2839
rect 28273 2805 28307 2839
rect 34621 2805 34655 2839
rect 5365 2601 5399 2635
rect 8585 2601 8619 2635
rect 20453 2601 20487 2635
rect 24593 2601 24627 2635
rect 29377 2601 29411 2635
rect 32137 2601 32171 2635
rect 33793 2601 33827 2635
rect 37933 2601 37967 2635
rect 2973 2533 3007 2567
rect 4537 2533 4571 2567
rect 5273 2533 5307 2567
rect 7205 2533 7239 2567
rect 10241 2533 10275 2567
rect 12909 2533 12943 2567
rect 13829 2533 13863 2567
rect 15209 2533 15243 2567
rect 16129 2533 16163 2567
rect 17877 2533 17911 2567
rect 19165 2533 19199 2567
rect 23765 2533 23799 2567
rect 24501 2533 24535 2567
rect 27353 2533 27387 2567
rect 35081 2533 35115 2567
rect 1501 2465 1535 2499
rect 2697 2465 2731 2499
rect 4261 2465 4295 2499
rect 6929 2465 6963 2499
rect 8401 2465 8435 2499
rect 9965 2465 9999 2499
rect 10885 2465 10919 2499
rect 12633 2465 12667 2499
rect 13553 2465 13587 2499
rect 14933 2465 14967 2499
rect 15853 2465 15887 2499
rect 17601 2465 17635 2499
rect 18889 2465 18923 2499
rect 20269 2465 20303 2499
rect 21557 2465 21591 2499
rect 23489 2465 23523 2499
rect 25605 2465 25639 2499
rect 26985 2465 27019 2499
rect 28365 2465 28399 2499
rect 29193 2465 29227 2499
rect 31033 2465 31067 2499
rect 31953 2465 31987 2499
rect 33609 2465 33643 2499
rect 34805 2465 34839 2499
rect 36553 2465 36587 2499
rect 37749 2465 37783 2499
rect 2053 2397 2087 2431
rect 11069 2397 11103 2431
rect 21741 2397 21775 2431
rect 25881 2397 25915 2431
rect 28641 2397 28675 2431
rect 36737 2397 36771 2431
rect 31217 2329 31251 2363
<< metal1 >>
rect 25498 117920 25504 117972
rect 25556 117960 25562 117972
rect 31110 117960 31116 117972
rect 25556 117932 31116 117960
rect 25556 117920 25562 117932
rect 31110 117920 31116 117932
rect 31168 117920 31174 117972
rect 35250 117920 35256 117972
rect 35308 117920 35314 117972
rect 24854 117716 24860 117768
rect 24912 117756 24918 117768
rect 29822 117756 29828 117768
rect 24912 117728 29828 117756
rect 24912 117716 24918 117728
rect 29822 117716 29828 117728
rect 29880 117716 29886 117768
rect 35268 117700 35296 117920
rect 4338 117648 4344 117700
rect 4396 117688 4402 117700
rect 4890 117688 4896 117700
rect 4396 117660 4896 117688
rect 4396 117648 4402 117660
rect 4890 117648 4896 117660
rect 4948 117648 4954 117700
rect 20346 117648 20352 117700
rect 20404 117688 20410 117700
rect 24670 117688 24676 117700
rect 20404 117660 24676 117688
rect 20404 117648 20410 117660
rect 24670 117648 24676 117660
rect 24728 117648 24734 117700
rect 35250 117648 35256 117700
rect 35308 117648 35314 117700
rect 18506 117580 18512 117632
rect 18564 117620 18570 117632
rect 19058 117620 19064 117632
rect 18564 117592 19064 117620
rect 18564 117580 18570 117592
rect 19058 117580 19064 117592
rect 19116 117580 19122 117632
rect 21634 117580 21640 117632
rect 21692 117620 21698 117632
rect 27246 117620 27252 117632
rect 21692 117592 27252 117620
rect 21692 117580 21698 117592
rect 27246 117580 27252 117592
rect 27304 117580 27310 117632
rect 1104 117530 38824 117552
rect 1104 117478 4246 117530
rect 4298 117478 4310 117530
rect 4362 117478 4374 117530
rect 4426 117478 4438 117530
rect 4490 117478 34966 117530
rect 35018 117478 35030 117530
rect 35082 117478 35094 117530
rect 35146 117478 35158 117530
rect 35210 117478 38824 117530
rect 1104 117456 38824 117478
rect 290 117376 296 117428
rect 348 117416 354 117428
rect 2685 117419 2743 117425
rect 2685 117416 2697 117419
rect 348 117388 2697 117416
rect 348 117376 354 117388
rect 2685 117385 2697 117388
rect 2731 117385 2743 117419
rect 2685 117379 2743 117385
rect 16574 117376 16580 117428
rect 16632 117416 16638 117428
rect 16632 117388 18644 117416
rect 16632 117376 16638 117388
rect 1118 117308 1124 117360
rect 1176 117348 1182 117360
rect 1176 117320 4660 117348
rect 1176 117308 1182 117320
rect 106 117240 112 117292
rect 164 117280 170 117292
rect 2041 117283 2099 117289
rect 2041 117280 2053 117283
rect 164 117252 2053 117280
rect 164 117240 170 117252
rect 2041 117249 2053 117252
rect 2087 117249 2099 117283
rect 4525 117283 4583 117289
rect 4525 117280 4537 117283
rect 2041 117243 2099 117249
rect 2746 117252 4537 117280
rect 658 117172 664 117224
rect 716 117212 722 117224
rect 2746 117212 2774 117252
rect 4525 117249 4537 117252
rect 4571 117249 4583 117283
rect 4632 117280 4660 117320
rect 12802 117308 12808 117360
rect 12860 117348 12866 117360
rect 12860 117320 13676 117348
rect 12860 117308 12866 117320
rect 5997 117283 6055 117289
rect 5997 117280 6009 117283
rect 4632 117252 6009 117280
rect 4525 117243 4583 117249
rect 5997 117249 6009 117252
rect 6043 117249 6055 117283
rect 5997 117243 6055 117249
rect 8294 117240 8300 117292
rect 8352 117280 8358 117292
rect 8573 117283 8631 117289
rect 8573 117280 8585 117283
rect 8352 117252 8585 117280
rect 8352 117240 8358 117252
rect 8573 117249 8585 117252
rect 8619 117249 8631 117283
rect 8573 117243 8631 117249
rect 8938 117240 8944 117292
rect 8996 117280 9002 117292
rect 9861 117283 9919 117289
rect 9861 117280 9873 117283
rect 8996 117252 9873 117280
rect 8996 117240 9002 117252
rect 9861 117249 9873 117252
rect 9907 117249 9919 117283
rect 9861 117243 9919 117249
rect 10226 117240 10232 117292
rect 10284 117280 10290 117292
rect 11333 117283 11391 117289
rect 11333 117280 11345 117283
rect 10284 117252 11345 117280
rect 10284 117240 10290 117252
rect 11333 117249 11345 117252
rect 11379 117249 11391 117283
rect 11333 117243 11391 117249
rect 11514 117240 11520 117292
rect 11572 117280 11578 117292
rect 13265 117283 13323 117289
rect 13265 117280 13277 117283
rect 11572 117252 13277 117280
rect 11572 117240 11578 117252
rect 13265 117249 13277 117252
rect 13311 117249 13323 117283
rect 13648 117280 13676 117320
rect 13998 117308 14004 117360
rect 14056 117348 14062 117360
rect 14056 117320 15332 117348
rect 14056 117308 14062 117320
rect 15197 117283 15255 117289
rect 15197 117280 15209 117283
rect 13648 117252 15209 117280
rect 13265 117243 13323 117249
rect 15197 117249 15209 117252
rect 15243 117249 15255 117283
rect 15304 117280 15332 117320
rect 15378 117308 15384 117360
rect 15436 117348 15442 117360
rect 18616 117348 18644 117388
rect 19794 117376 19800 117428
rect 19852 117416 19858 117428
rect 20254 117416 20260 117428
rect 19852 117388 20260 117416
rect 19852 117376 19858 117388
rect 20254 117376 20260 117388
rect 20312 117376 20318 117428
rect 20990 117376 20996 117428
rect 21048 117416 21054 117428
rect 21048 117388 22094 117416
rect 21048 117376 21054 117388
rect 15436 117320 16804 117348
rect 18616 117320 18736 117348
rect 15436 117308 15442 117320
rect 16669 117283 16727 117289
rect 16669 117280 16681 117283
rect 15304 117252 16681 117280
rect 15197 117243 15255 117249
rect 16669 117249 16681 117252
rect 16715 117249 16727 117283
rect 16776 117280 16804 117320
rect 18601 117283 18659 117289
rect 18601 117280 18613 117283
rect 16776 117252 18613 117280
rect 16669 117243 16727 117249
rect 18601 117249 18613 117252
rect 18647 117249 18659 117283
rect 18708 117280 18736 117320
rect 19058 117308 19064 117360
rect 19116 117348 19122 117360
rect 19886 117348 19892 117360
rect 19116 117320 19892 117348
rect 19116 117308 19122 117320
rect 19886 117308 19892 117320
rect 19944 117308 19950 117360
rect 20533 117283 20591 117289
rect 20533 117280 20545 117283
rect 18708 117252 20545 117280
rect 18601 117243 18659 117249
rect 20533 117249 20545 117252
rect 20579 117249 20591 117283
rect 22066 117280 22094 117388
rect 22370 117376 22376 117428
rect 22428 117416 22434 117428
rect 23845 117419 23903 117425
rect 23845 117416 23857 117419
rect 22428 117388 23857 117416
rect 22428 117376 22434 117388
rect 23845 117385 23857 117388
rect 23891 117385 23903 117419
rect 27246 117416 27252 117428
rect 27207 117388 27252 117416
rect 23845 117379 23903 117385
rect 27246 117376 27252 117388
rect 27304 117376 27310 117428
rect 29822 117376 29828 117428
rect 29880 117416 29886 117428
rect 29917 117419 29975 117425
rect 29917 117416 29929 117419
rect 29880 117388 29929 117416
rect 29880 117376 29886 117388
rect 29917 117385 29929 117388
rect 29963 117385 29975 117419
rect 31110 117416 31116 117428
rect 31071 117388 31116 117416
rect 29917 117379 29975 117385
rect 31110 117376 31116 117388
rect 31168 117376 31174 117428
rect 34146 117376 34152 117428
rect 34204 117416 34210 117428
rect 34333 117419 34391 117425
rect 34333 117416 34345 117419
rect 34204 117388 34345 117416
rect 34204 117376 34210 117388
rect 34333 117385 34345 117388
rect 34379 117385 34391 117419
rect 34333 117379 34391 117385
rect 22922 117308 22928 117360
rect 22980 117348 22986 117360
rect 28537 117351 28595 117357
rect 28537 117348 28549 117351
rect 22980 117320 28549 117348
rect 22980 117308 22986 117320
rect 28537 117317 28549 117320
rect 28583 117317 28595 117351
rect 28537 117311 28595 117317
rect 26605 117283 26663 117289
rect 26605 117280 26617 117283
rect 22066 117252 26617 117280
rect 20533 117243 20591 117249
rect 26605 117249 26617 117252
rect 26651 117249 26663 117283
rect 26605 117243 26663 117249
rect 31941 117283 31999 117289
rect 31941 117249 31953 117283
rect 31987 117280 31999 117283
rect 34330 117280 34336 117292
rect 31987 117252 34336 117280
rect 31987 117249 31999 117252
rect 31941 117243 31999 117249
rect 34330 117240 34336 117252
rect 34388 117240 34394 117292
rect 35345 117283 35403 117289
rect 35345 117249 35357 117283
rect 35391 117280 35403 117283
rect 36262 117280 36268 117292
rect 35391 117252 36268 117280
rect 35391 117249 35403 117252
rect 35345 117243 35403 117249
rect 36262 117240 36268 117252
rect 36320 117240 36326 117292
rect 36538 117280 36544 117292
rect 36499 117252 36544 117280
rect 36538 117240 36544 117252
rect 36596 117240 36602 117292
rect 5261 117215 5319 117221
rect 5261 117212 5273 117215
rect 716 117184 2774 117212
rect 4172 117184 5273 117212
rect 716 117172 722 117184
rect 1854 117144 1860 117156
rect 1815 117116 1860 117144
rect 1854 117104 1860 117116
rect 1912 117104 1918 117156
rect 2593 117147 2651 117153
rect 2593 117113 2605 117147
rect 2639 117144 2651 117147
rect 3602 117144 3608 117156
rect 2639 117116 3608 117144
rect 2639 117113 2651 117116
rect 2593 117107 2651 117113
rect 3602 117104 3608 117116
rect 3660 117104 3666 117156
rect 934 117036 940 117088
rect 992 117076 998 117088
rect 4172 117076 4200 117184
rect 5261 117181 5273 117184
rect 5307 117181 5319 117215
rect 7834 117212 7840 117224
rect 7795 117184 7840 117212
rect 5261 117175 5319 117181
rect 7834 117172 7840 117184
rect 7892 117172 7898 117224
rect 9582 117172 9588 117224
rect 9640 117212 9646 117224
rect 10597 117215 10655 117221
rect 10597 117212 10609 117215
rect 9640 117184 10609 117212
rect 9640 117172 9646 117184
rect 10597 117181 10609 117184
rect 10643 117181 10655 117215
rect 10597 117175 10655 117181
rect 10870 117172 10876 117224
rect 10928 117212 10934 117224
rect 12529 117215 12587 117221
rect 12529 117212 12541 117215
rect 10928 117184 12541 117212
rect 10928 117172 10934 117184
rect 12529 117181 12541 117184
rect 12575 117181 12587 117215
rect 14001 117215 14059 117221
rect 14001 117212 14013 117215
rect 12529 117175 12587 117181
rect 13188 117184 14013 117212
rect 4341 117147 4399 117153
rect 4341 117113 4353 117147
rect 4387 117113 4399 117147
rect 5074 117144 5080 117156
rect 5035 117116 5080 117144
rect 4341 117107 4399 117113
rect 992 117048 4200 117076
rect 4356 117076 4384 117107
rect 5074 117104 5080 117116
rect 5132 117104 5138 117156
rect 5813 117147 5871 117153
rect 5813 117113 5825 117147
rect 5859 117144 5871 117147
rect 6730 117144 6736 117156
rect 5859 117116 6736 117144
rect 5859 117113 5871 117116
rect 5813 117107 5871 117113
rect 6730 117104 6736 117116
rect 6788 117104 6794 117156
rect 7009 117147 7067 117153
rect 7009 117113 7021 117147
rect 7055 117144 7067 117147
rect 8110 117144 8116 117156
rect 7055 117116 8116 117144
rect 7055 117113 7067 117116
rect 7009 117107 7067 117113
rect 8110 117104 8116 117116
rect 8168 117104 8174 117156
rect 8386 117144 8392 117156
rect 8347 117116 8392 117144
rect 8386 117104 8392 117116
rect 8444 117104 8450 117156
rect 9490 117104 9496 117156
rect 9548 117144 9554 117156
rect 9677 117147 9735 117153
rect 9677 117144 9689 117147
rect 9548 117116 9689 117144
rect 9548 117104 9554 117116
rect 9677 117113 9689 117116
rect 9723 117113 9735 117147
rect 9677 117107 9735 117113
rect 9766 117104 9772 117156
rect 9824 117144 9830 117156
rect 10413 117147 10471 117153
rect 10413 117144 10425 117147
rect 9824 117116 10425 117144
rect 9824 117104 9830 117116
rect 10413 117113 10425 117116
rect 10459 117113 10471 117147
rect 11146 117144 11152 117156
rect 11107 117116 11152 117144
rect 10413 117107 10471 117113
rect 11146 117104 11152 117116
rect 11204 117104 11210 117156
rect 11330 117104 11336 117156
rect 11388 117144 11394 117156
rect 12345 117147 12403 117153
rect 12345 117144 12357 117147
rect 11388 117116 12357 117144
rect 11388 117104 11394 117116
rect 12345 117113 12357 117116
rect 12391 117113 12403 117147
rect 13078 117144 13084 117156
rect 13039 117116 13084 117144
rect 12345 117107 12403 117113
rect 13078 117104 13084 117116
rect 13136 117104 13142 117156
rect 5258 117076 5264 117088
rect 4356 117048 5264 117076
rect 992 117036 998 117048
rect 5258 117036 5264 117048
rect 5316 117036 5322 117088
rect 5902 117036 5908 117088
rect 5960 117076 5966 117088
rect 7101 117079 7159 117085
rect 7101 117076 7113 117079
rect 5960 117048 7113 117076
rect 5960 117036 5966 117048
rect 7101 117045 7113 117048
rect 7147 117045 7159 117079
rect 7101 117039 7159 117045
rect 12158 117036 12164 117088
rect 12216 117076 12222 117088
rect 13188 117076 13216 117184
rect 14001 117181 14013 117184
rect 14047 117181 14059 117215
rect 14001 117175 14059 117181
rect 14090 117172 14096 117224
rect 14148 117212 14154 117224
rect 15749 117215 15807 117221
rect 15749 117212 15761 117215
rect 14148 117184 15761 117212
rect 14148 117172 14154 117184
rect 15749 117181 15761 117184
rect 15795 117181 15807 117215
rect 15749 117175 15807 117181
rect 15838 117172 15844 117224
rect 15896 117212 15902 117224
rect 17681 117215 17739 117221
rect 17681 117212 17693 117215
rect 15896 117184 17693 117212
rect 15896 117172 15902 117184
rect 17681 117181 17693 117184
rect 17727 117181 17739 117215
rect 17681 117175 17739 117181
rect 17770 117172 17776 117224
rect 17828 117212 17834 117224
rect 19153 117215 19211 117221
rect 19153 117212 19165 117215
rect 17828 117184 19165 117212
rect 17828 117172 17834 117184
rect 19153 117181 19165 117184
rect 19199 117181 19211 117215
rect 19153 117175 19211 117181
rect 19334 117172 19340 117224
rect 19392 117212 19398 117224
rect 20438 117212 20444 117224
rect 19392 117184 20444 117212
rect 19392 117172 19398 117184
rect 20438 117172 20444 117184
rect 20496 117172 20502 117224
rect 21634 117172 21640 117224
rect 21692 117212 21698 117224
rect 21692 117184 21956 117212
rect 21692 117172 21698 117184
rect 13814 117144 13820 117156
rect 13775 117116 13820 117144
rect 13814 117104 13820 117116
rect 13872 117104 13878 117156
rect 15010 117144 15016 117156
rect 14971 117116 15016 117144
rect 15010 117104 15016 117116
rect 15068 117104 15074 117156
rect 15930 117104 15936 117156
rect 15988 117144 15994 117156
rect 16485 117147 16543 117153
rect 16485 117144 16497 117147
rect 15988 117116 16497 117144
rect 15988 117104 15994 117116
rect 16485 117113 16497 117116
rect 16531 117113 16543 117147
rect 16485 117107 16543 117113
rect 16574 117104 16580 117156
rect 16632 117144 16638 117156
rect 18417 117147 18475 117153
rect 18417 117144 18429 117147
rect 16632 117116 18429 117144
rect 16632 117104 16638 117116
rect 18417 117113 18429 117116
rect 18463 117113 18475 117147
rect 18417 117107 18475 117113
rect 19058 117104 19064 117156
rect 19116 117144 19122 117156
rect 19116 117116 19380 117144
rect 19116 117104 19122 117116
rect 12216 117048 13216 117076
rect 12216 117036 12222 117048
rect 13446 117036 13452 117088
rect 13504 117076 13510 117088
rect 15841 117079 15899 117085
rect 15841 117076 15853 117079
rect 13504 117048 15853 117076
rect 13504 117036 13510 117048
rect 15841 117045 15853 117048
rect 15887 117045 15899 117079
rect 15841 117039 15899 117045
rect 16298 117036 16304 117088
rect 16356 117076 16362 117088
rect 17773 117079 17831 117085
rect 17773 117076 17785 117079
rect 16356 117048 17785 117076
rect 16356 117036 16362 117048
rect 17773 117045 17785 117048
rect 17819 117045 17831 117079
rect 17773 117039 17831 117045
rect 17862 117036 17868 117088
rect 17920 117076 17926 117088
rect 19245 117079 19303 117085
rect 19245 117076 19257 117079
rect 17920 117048 19257 117076
rect 17920 117036 17926 117048
rect 19245 117045 19257 117048
rect 19291 117045 19303 117079
rect 19352 117076 19380 117116
rect 19886 117104 19892 117156
rect 19944 117144 19950 117156
rect 20349 117147 20407 117153
rect 20349 117144 20361 117147
rect 19944 117116 20361 117144
rect 19944 117104 19950 117116
rect 20349 117113 20361 117116
rect 20395 117113 20407 117147
rect 20349 117107 20407 117113
rect 20530 117104 20536 117156
rect 20588 117144 20594 117156
rect 21085 117147 21143 117153
rect 21085 117144 21097 117147
rect 20588 117116 21097 117144
rect 20588 117104 20594 117116
rect 21085 117113 21097 117116
rect 21131 117113 21143 117147
rect 21085 117107 21143 117113
rect 21358 117104 21364 117156
rect 21416 117144 21422 117156
rect 21821 117147 21879 117153
rect 21821 117144 21833 117147
rect 21416 117116 21833 117144
rect 21416 117104 21422 117116
rect 21821 117113 21833 117116
rect 21867 117113 21879 117147
rect 21928 117144 21956 117184
rect 22002 117172 22008 117224
rect 22060 117212 22066 117224
rect 23017 117215 23075 117221
rect 23017 117212 23029 117215
rect 22060 117184 23029 117212
rect 22060 117172 22066 117184
rect 23017 117181 23029 117184
rect 23063 117181 23075 117215
rect 26421 117215 26479 117221
rect 26421 117212 26433 117215
rect 23017 117175 23075 117181
rect 23860 117184 26433 117212
rect 23198 117144 23204 117156
rect 21928 117116 22048 117144
rect 23159 117116 23204 117144
rect 21821 117107 21879 117113
rect 21177 117079 21235 117085
rect 21177 117076 21189 117079
rect 19352 117048 21189 117076
rect 19245 117039 19303 117045
rect 21177 117045 21189 117048
rect 21223 117045 21235 117079
rect 21177 117039 21235 117045
rect 21726 117036 21732 117088
rect 21784 117076 21790 117088
rect 21913 117079 21971 117085
rect 21913 117076 21925 117079
rect 21784 117048 21925 117076
rect 21784 117036 21790 117048
rect 21913 117045 21925 117048
rect 21959 117045 21971 117079
rect 22020 117076 22048 117116
rect 23198 117104 23204 117116
rect 23256 117104 23262 117156
rect 23290 117104 23296 117156
rect 23348 117144 23354 117156
rect 23753 117147 23811 117153
rect 23753 117144 23765 117147
rect 23348 117116 23765 117144
rect 23348 117104 23354 117116
rect 23753 117113 23765 117116
rect 23799 117113 23811 117147
rect 23753 117107 23811 117113
rect 23860 117076 23888 117184
rect 26421 117181 26433 117184
rect 26467 117181 26479 117215
rect 26421 117175 26479 117181
rect 26694 117172 26700 117224
rect 26752 117212 26758 117224
rect 29825 117215 29883 117221
rect 29825 117212 29837 117215
rect 26752 117184 29837 117212
rect 26752 117172 26758 117184
rect 29825 117181 29837 117184
rect 29871 117181 29883 117215
rect 29825 117175 29883 117181
rect 32677 117215 32735 117221
rect 32677 117181 32689 117215
rect 32723 117212 32735 117215
rect 32723 117184 34514 117212
rect 32723 117181 32735 117184
rect 32677 117175 32735 117181
rect 24118 117104 24124 117156
rect 24176 117144 24182 117156
rect 24489 117147 24547 117153
rect 24489 117144 24501 117147
rect 24176 117116 24501 117144
rect 24176 117104 24182 117116
rect 24489 117113 24501 117116
rect 24535 117113 24547 117147
rect 24489 117107 24547 117113
rect 24762 117104 24768 117156
rect 24820 117144 24826 117156
rect 25685 117147 25743 117153
rect 25685 117144 25697 117147
rect 24820 117116 25697 117144
rect 24820 117104 24826 117116
rect 25685 117113 25697 117116
rect 25731 117113 25743 117147
rect 27154 117144 27160 117156
rect 27115 117116 27160 117144
rect 25685 117107 25743 117113
rect 27154 117104 27160 117116
rect 27212 117104 27218 117156
rect 28350 117144 28356 117156
rect 28311 117116 28356 117144
rect 28350 117104 28356 117116
rect 28408 117104 28414 117156
rect 29089 117147 29147 117153
rect 29089 117113 29101 117147
rect 29135 117113 29147 117147
rect 29089 117107 29147 117113
rect 22020 117048 23888 117076
rect 21913 117039 21971 117045
rect 23934 117036 23940 117088
rect 23992 117076 23998 117088
rect 24581 117079 24639 117085
rect 24581 117076 24593 117079
rect 23992 117048 24593 117076
rect 23992 117036 23998 117048
rect 24581 117045 24593 117048
rect 24627 117045 24639 117079
rect 24581 117039 24639 117045
rect 24670 117036 24676 117088
rect 24728 117076 24734 117088
rect 25777 117079 25835 117085
rect 25777 117076 25789 117079
rect 24728 117048 25789 117076
rect 24728 117036 24734 117048
rect 25777 117045 25789 117048
rect 25823 117045 25835 117079
rect 25777 117039 25835 117045
rect 25958 117036 25964 117088
rect 26016 117076 26022 117088
rect 29104 117076 29132 117107
rect 30650 117104 30656 117156
rect 30708 117144 30714 117156
rect 31021 117147 31079 117153
rect 31021 117144 31033 117147
rect 30708 117116 31033 117144
rect 30708 117104 30714 117116
rect 31021 117113 31033 117116
rect 31067 117113 31079 117147
rect 31754 117144 31760 117156
rect 31715 117116 31760 117144
rect 31021 117107 31079 117113
rect 31754 117104 31760 117116
rect 31812 117104 31818 117156
rect 32306 117104 32312 117156
rect 32364 117144 32370 117156
rect 32493 117147 32551 117153
rect 32493 117144 32505 117147
rect 32364 117116 32505 117144
rect 32364 117104 32370 117116
rect 32493 117113 32505 117116
rect 32539 117113 32551 117147
rect 34238 117144 34244 117156
rect 34199 117116 34244 117144
rect 32493 117107 32551 117113
rect 34238 117104 34244 117116
rect 34296 117104 34302 117156
rect 26016 117048 29132 117076
rect 26016 117036 26022 117048
rect 29178 117036 29184 117088
rect 29236 117076 29242 117088
rect 34486 117076 34514 117184
rect 34974 117172 34980 117224
rect 35032 117212 35038 117224
rect 36357 117215 36415 117221
rect 35032 117184 35756 117212
rect 35032 117172 35038 117184
rect 35161 117147 35219 117153
rect 35161 117113 35173 117147
rect 35207 117144 35219 117147
rect 35618 117144 35624 117156
rect 35207 117116 35624 117144
rect 35207 117113 35219 117116
rect 35161 117107 35219 117113
rect 35618 117104 35624 117116
rect 35676 117104 35682 117156
rect 35728 117144 35756 117184
rect 36357 117181 36369 117215
rect 36403 117212 36415 117215
rect 37090 117212 37096 117224
rect 36403 117184 37096 117212
rect 36403 117181 36415 117184
rect 36357 117175 36415 117181
rect 37090 117172 37096 117184
rect 37148 117172 37154 117224
rect 37369 117215 37427 117221
rect 37369 117181 37381 117215
rect 37415 117212 37427 117215
rect 37734 117212 37740 117224
rect 37415 117184 37740 117212
rect 37415 117181 37427 117184
rect 37369 117175 37427 117181
rect 37734 117172 37740 117184
rect 37792 117172 37798 117224
rect 37918 117144 37924 117156
rect 35728 117116 36584 117144
rect 37879 117116 37924 117144
rect 36446 117076 36452 117088
rect 29236 117048 29281 117076
rect 34486 117048 36452 117076
rect 29236 117036 29242 117048
rect 36446 117036 36452 117048
rect 36504 117036 36510 117088
rect 36556 117076 36584 117116
rect 37918 117104 37924 117116
rect 37976 117104 37982 117156
rect 39022 117076 39028 117088
rect 36556 117048 39028 117076
rect 39022 117036 39028 117048
rect 39080 117036 39086 117088
rect 1104 116986 38824 117008
rect 1104 116934 19606 116986
rect 19658 116934 19670 116986
rect 19722 116934 19734 116986
rect 19786 116934 19798 116986
rect 19850 116934 38824 116986
rect 1104 116912 38824 116934
rect 1302 116832 1308 116884
rect 1360 116872 1366 116884
rect 1949 116875 2007 116881
rect 1949 116872 1961 116875
rect 1360 116844 1961 116872
rect 1360 116832 1366 116844
rect 1949 116841 1961 116844
rect 1995 116841 2007 116875
rect 1949 116835 2007 116841
rect 2590 116832 2596 116884
rect 2648 116872 2654 116884
rect 4157 116875 4215 116881
rect 4157 116872 4169 116875
rect 2648 116844 4169 116872
rect 2648 116832 2654 116844
rect 4157 116841 4169 116844
rect 4203 116841 4215 116875
rect 4157 116835 4215 116841
rect 6454 116832 6460 116884
rect 6512 116872 6518 116884
rect 7009 116875 7067 116881
rect 7009 116872 7021 116875
rect 6512 116844 7021 116872
rect 6512 116832 6518 116844
rect 7009 116841 7021 116844
rect 7055 116841 7067 116875
rect 7009 116835 7067 116841
rect 7098 116832 7104 116884
rect 7156 116872 7162 116884
rect 7745 116875 7803 116881
rect 7745 116872 7757 116875
rect 7156 116844 7757 116872
rect 7156 116832 7162 116844
rect 7745 116841 7757 116844
rect 7791 116841 7803 116875
rect 7745 116835 7803 116841
rect 8570 116832 8576 116884
rect 8628 116872 8634 116884
rect 9217 116875 9275 116881
rect 9217 116872 9229 116875
rect 8628 116844 9229 116872
rect 8628 116832 8634 116844
rect 9217 116841 9229 116844
rect 9263 116841 9275 116875
rect 9217 116835 9275 116841
rect 9306 116832 9312 116884
rect 9364 116872 9370 116884
rect 9953 116875 10011 116881
rect 9953 116872 9965 116875
rect 9364 116844 9965 116872
rect 9364 116832 9370 116844
rect 9953 116841 9965 116844
rect 9999 116841 10011 116875
rect 9953 116835 10011 116841
rect 11698 116832 11704 116884
rect 11756 116872 11762 116884
rect 12253 116875 12311 116881
rect 12253 116872 12265 116875
rect 11756 116844 12265 116872
rect 11756 116832 11762 116844
rect 12253 116841 12265 116844
rect 12299 116841 12311 116875
rect 12253 116835 12311 116841
rect 12434 116832 12440 116884
rect 12492 116872 12498 116884
rect 12989 116875 13047 116881
rect 12989 116872 13001 116875
rect 12492 116844 13001 116872
rect 12492 116832 12498 116844
rect 12989 116841 13001 116844
rect 13035 116841 13047 116875
rect 12989 116835 13047 116841
rect 13630 116832 13636 116884
rect 13688 116872 13694 116884
rect 14461 116875 14519 116881
rect 14461 116872 14473 116875
rect 13688 116844 14473 116872
rect 13688 116832 13694 116844
rect 14461 116841 14473 116844
rect 14507 116841 14519 116875
rect 14461 116835 14519 116841
rect 14734 116832 14740 116884
rect 14792 116872 14798 116884
rect 15933 116875 15991 116881
rect 15933 116872 15945 116875
rect 14792 116844 15945 116872
rect 14792 116832 14798 116844
rect 15933 116841 15945 116844
rect 15979 116841 15991 116875
rect 15933 116835 15991 116841
rect 16758 116832 16764 116884
rect 16816 116872 16822 116884
rect 17497 116875 17555 116881
rect 17497 116872 17509 116875
rect 16816 116844 17509 116872
rect 16816 116832 16822 116844
rect 17497 116841 17509 116844
rect 17543 116841 17555 116875
rect 17497 116835 17555 116841
rect 17586 116832 17592 116884
rect 17644 116872 17650 116884
rect 18233 116875 18291 116881
rect 18233 116872 18245 116875
rect 17644 116844 18245 116872
rect 17644 116832 17650 116844
rect 18233 116841 18245 116844
rect 18279 116841 18291 116875
rect 18233 116835 18291 116841
rect 18690 116832 18696 116884
rect 18748 116872 18754 116884
rect 19705 116875 19763 116881
rect 19705 116872 19717 116875
rect 18748 116844 19717 116872
rect 18748 116832 18754 116844
rect 19705 116841 19717 116844
rect 19751 116841 19763 116875
rect 20438 116872 20444 116884
rect 20399 116844 20444 116872
rect 19705 116835 19763 116841
rect 20438 116832 20444 116844
rect 20496 116832 20502 116884
rect 20714 116832 20720 116884
rect 20772 116872 20778 116884
rect 21177 116875 21235 116881
rect 21177 116872 21189 116875
rect 20772 116844 21189 116872
rect 20772 116832 20778 116844
rect 21177 116841 21189 116844
rect 21223 116841 21235 116875
rect 21177 116835 21235 116841
rect 22278 116832 22284 116884
rect 22336 116872 22342 116884
rect 22741 116875 22799 116881
rect 22741 116872 22753 116875
rect 22336 116844 22753 116872
rect 22336 116832 22342 116844
rect 22741 116841 22753 116844
rect 22787 116841 22799 116875
rect 23658 116872 23664 116884
rect 22741 116835 22799 116841
rect 23308 116844 23664 116872
rect 2130 116764 2136 116816
rect 2188 116804 2194 116816
rect 2777 116807 2835 116813
rect 2777 116804 2789 116807
rect 2188 116776 2789 116804
rect 2188 116764 2194 116776
rect 2777 116773 2789 116776
rect 2823 116773 2835 116807
rect 2777 116767 2835 116773
rect 3234 116764 3240 116816
rect 3292 116804 3298 116816
rect 4985 116807 5043 116813
rect 4985 116804 4997 116807
rect 3292 116776 4997 116804
rect 3292 116764 3298 116776
rect 4985 116773 4997 116776
rect 5031 116773 5043 116807
rect 4985 116767 5043 116773
rect 7834 116764 7840 116816
rect 7892 116804 7898 116816
rect 8389 116807 8447 116813
rect 8389 116804 8401 116807
rect 7892 116776 8401 116804
rect 7892 116764 7898 116776
rect 8389 116773 8401 116776
rect 8435 116773 8447 116807
rect 8389 116767 8447 116773
rect 9674 116764 9680 116816
rect 9732 116804 9738 116816
rect 10781 116807 10839 116813
rect 10781 116804 10793 116807
rect 9732 116776 10793 116804
rect 9732 116764 9738 116776
rect 10781 116773 10793 116776
rect 10827 116773 10839 116807
rect 10781 116767 10839 116773
rect 13170 116764 13176 116816
rect 13228 116804 13234 116816
rect 13817 116807 13875 116813
rect 13817 116804 13829 116807
rect 13228 116776 13829 116804
rect 13228 116764 13234 116776
rect 13817 116773 13829 116776
rect 13863 116773 13875 116807
rect 13817 116767 13875 116773
rect 14274 116764 14280 116816
rect 14332 116804 14338 116816
rect 15289 116807 15347 116813
rect 15289 116804 15301 116807
rect 14332 116776 15301 116804
rect 14332 116764 14338 116776
rect 15289 116773 15301 116776
rect 15335 116773 15347 116807
rect 15289 116767 15347 116773
rect 16022 116764 16028 116816
rect 16080 116804 16086 116816
rect 17862 116804 17868 116816
rect 16080 116776 17868 116804
rect 16080 116764 16086 116776
rect 17862 116764 17868 116776
rect 17920 116764 17926 116816
rect 18046 116764 18052 116816
rect 18104 116804 18110 116816
rect 19061 116807 19119 116813
rect 19061 116804 19073 116807
rect 18104 116776 19073 116804
rect 18104 116764 18110 116776
rect 19061 116773 19073 116776
rect 19107 116773 19119 116807
rect 19061 116767 19119 116773
rect 19150 116764 19156 116816
rect 19208 116804 19214 116816
rect 22370 116804 22376 116816
rect 19208 116776 22376 116804
rect 19208 116764 19214 116776
rect 22370 116764 22376 116776
rect 22428 116764 22434 116816
rect 22646 116813 22652 116816
rect 22632 116807 22652 116813
rect 22632 116773 22644 116807
rect 22632 116767 22652 116773
rect 22646 116764 22652 116767
rect 22704 116764 22710 116816
rect 1857 116739 1915 116745
rect 1857 116705 1869 116739
rect 1903 116705 1915 116739
rect 2590 116736 2596 116748
rect 2551 116708 2596 116736
rect 1857 116699 1915 116705
rect 1872 116600 1900 116699
rect 2590 116696 2596 116708
rect 2648 116696 2654 116748
rect 3329 116739 3387 116745
rect 3329 116705 3341 116739
rect 3375 116736 3387 116739
rect 3786 116736 3792 116748
rect 3375 116708 3792 116736
rect 3375 116705 3387 116708
rect 3329 116699 3387 116705
rect 3786 116696 3792 116708
rect 3844 116696 3850 116748
rect 4062 116736 4068 116748
rect 4023 116708 4068 116736
rect 4062 116696 4068 116708
rect 4120 116696 4126 116748
rect 4798 116736 4804 116748
rect 4759 116708 4804 116736
rect 4798 116696 4804 116708
rect 4856 116696 4862 116748
rect 5534 116736 5540 116748
rect 5495 116708 5540 116736
rect 5534 116696 5540 116708
rect 5592 116696 5598 116748
rect 6914 116736 6920 116748
rect 6875 116708 6920 116736
rect 6914 116696 6920 116708
rect 6972 116696 6978 116748
rect 7006 116696 7012 116748
rect 7064 116736 7070 116748
rect 7653 116739 7711 116745
rect 7653 116736 7665 116739
rect 7064 116708 7665 116736
rect 7064 116696 7070 116708
rect 7653 116705 7665 116708
rect 7699 116705 7711 116739
rect 7653 116699 7711 116705
rect 8570 116696 8576 116748
rect 8628 116736 8634 116748
rect 9125 116739 9183 116745
rect 9125 116736 9137 116739
rect 8628 116708 9137 116736
rect 8628 116696 8634 116708
rect 9125 116705 9137 116708
rect 9171 116705 9183 116739
rect 9858 116736 9864 116748
rect 9819 116708 9864 116736
rect 9125 116699 9183 116705
rect 9858 116696 9864 116708
rect 9916 116696 9922 116748
rect 10594 116736 10600 116748
rect 10555 116708 10600 116736
rect 10594 116696 10600 116708
rect 10652 116696 10658 116748
rect 12158 116736 12164 116748
rect 12119 116708 12164 116736
rect 12158 116696 12164 116708
rect 12216 116696 12222 116748
rect 12894 116736 12900 116748
rect 12855 116708 12900 116736
rect 12894 116696 12900 116708
rect 12952 116696 12958 116748
rect 12986 116696 12992 116748
rect 13044 116736 13050 116748
rect 13633 116739 13691 116745
rect 13633 116736 13645 116739
rect 13044 116708 13645 116736
rect 13044 116696 13050 116708
rect 13633 116705 13645 116708
rect 13679 116705 13691 116739
rect 14366 116736 14372 116748
rect 14327 116708 14372 116736
rect 13633 116699 13691 116705
rect 14366 116696 14372 116708
rect 14424 116696 14430 116748
rect 15102 116736 15108 116748
rect 15063 116708 15108 116736
rect 15102 116696 15108 116708
rect 15160 116696 15166 116748
rect 15562 116696 15568 116748
rect 15620 116736 15626 116748
rect 15841 116739 15899 116745
rect 15841 116736 15853 116739
rect 15620 116708 15853 116736
rect 15620 116696 15626 116708
rect 15841 116705 15853 116708
rect 15887 116705 15899 116739
rect 17402 116736 17408 116748
rect 17363 116708 17408 116736
rect 15841 116699 15899 116705
rect 17402 116696 17408 116708
rect 17460 116696 17466 116748
rect 18138 116736 18144 116748
rect 18099 116708 18144 116736
rect 18138 116696 18144 116708
rect 18196 116696 18202 116748
rect 18874 116736 18880 116748
rect 18835 116708 18880 116736
rect 18874 116696 18880 116708
rect 18932 116696 18938 116748
rect 19334 116696 19340 116748
rect 19392 116736 19398 116748
rect 19613 116739 19671 116745
rect 19613 116736 19625 116739
rect 19392 116708 19625 116736
rect 19392 116696 19398 116708
rect 19613 116705 19625 116708
rect 19659 116705 19671 116739
rect 20346 116736 20352 116748
rect 20307 116708 20352 116736
rect 19613 116699 19671 116705
rect 20346 116696 20352 116708
rect 20404 116696 20410 116748
rect 21085 116739 21143 116745
rect 21085 116705 21097 116739
rect 21131 116736 21143 116739
rect 23308 116736 23336 116844
rect 23658 116832 23664 116844
rect 23716 116832 23722 116884
rect 24210 116832 24216 116884
rect 24268 116872 24274 116884
rect 24397 116875 24455 116881
rect 24397 116872 24409 116875
rect 24268 116844 24409 116872
rect 24268 116832 24274 116844
rect 24397 116841 24409 116844
rect 24443 116841 24455 116875
rect 24397 116835 24455 116841
rect 24486 116832 24492 116884
rect 24544 116872 24550 116884
rect 25133 116875 25191 116881
rect 25133 116872 25145 116875
rect 24544 116844 25145 116872
rect 24544 116832 24550 116844
rect 25133 116841 25145 116844
rect 25179 116841 25191 116875
rect 25133 116835 25191 116841
rect 25682 116832 25688 116884
rect 25740 116872 25746 116884
rect 26605 116875 26663 116881
rect 26605 116872 26617 116875
rect 25740 116844 26617 116872
rect 25740 116832 25746 116844
rect 26605 116841 26617 116844
rect 26651 116841 26663 116875
rect 26605 116835 26663 116841
rect 26786 116832 26792 116884
rect 26844 116872 26850 116884
rect 28721 116875 28779 116881
rect 28721 116872 28733 116875
rect 26844 116844 28733 116872
rect 26844 116832 26850 116844
rect 28721 116841 28733 116844
rect 28767 116841 28779 116875
rect 28721 116835 28779 116841
rect 29086 116832 29092 116884
rect 29144 116872 29150 116884
rect 30006 116872 30012 116884
rect 29144 116844 30012 116872
rect 29144 116832 29150 116844
rect 30006 116832 30012 116844
rect 30064 116832 30070 116884
rect 31573 116875 31631 116881
rect 31573 116872 31585 116875
rect 30116 116844 31585 116872
rect 26050 116804 26056 116816
rect 24136 116776 26056 116804
rect 21131 116708 23336 116736
rect 23385 116739 23443 116745
rect 21131 116705 21143 116708
rect 21085 116699 21143 116705
rect 23385 116705 23397 116739
rect 23431 116736 23443 116739
rect 24136 116736 24164 116776
rect 26050 116764 26056 116776
rect 26108 116764 26114 116816
rect 26142 116764 26148 116816
rect 26200 116804 26206 116816
rect 28077 116807 28135 116813
rect 28077 116804 28089 116807
rect 26200 116776 28089 116804
rect 26200 116764 26206 116776
rect 28077 116773 28089 116776
rect 28123 116773 28135 116807
rect 28077 116767 28135 116773
rect 28534 116764 28540 116816
rect 28592 116804 28598 116816
rect 30116 116804 30144 116844
rect 31573 116841 31585 116844
rect 31619 116841 31631 116875
rect 31573 116835 31631 116841
rect 34606 116832 34612 116884
rect 34664 116872 34670 116884
rect 34793 116875 34851 116881
rect 34793 116872 34805 116875
rect 34664 116844 34805 116872
rect 34664 116832 34670 116844
rect 34793 116841 34805 116844
rect 34839 116841 34851 116875
rect 34793 116835 34851 116841
rect 34882 116832 34888 116884
rect 34940 116872 34946 116884
rect 35529 116875 35587 116881
rect 35529 116872 35541 116875
rect 34940 116844 35541 116872
rect 34940 116832 34946 116844
rect 35529 116841 35541 116844
rect 35575 116841 35587 116875
rect 35529 116835 35587 116841
rect 28592 116776 30144 116804
rect 28592 116764 28598 116776
rect 31018 116764 31024 116816
rect 31076 116804 31082 116816
rect 33042 116804 33048 116816
rect 31076 116776 33048 116804
rect 31076 116764 31082 116776
rect 33042 116764 33048 116776
rect 33100 116764 33106 116816
rect 33413 116807 33471 116813
rect 33413 116773 33425 116807
rect 33459 116804 33471 116807
rect 34974 116804 34980 116816
rect 33459 116776 34980 116804
rect 33459 116773 33471 116776
rect 33413 116767 33471 116773
rect 34974 116764 34980 116776
rect 35032 116764 35038 116816
rect 35342 116764 35348 116816
rect 35400 116804 35406 116816
rect 36357 116807 36415 116813
rect 36357 116804 36369 116807
rect 35400 116776 36369 116804
rect 35400 116764 35406 116776
rect 36357 116773 36369 116776
rect 36403 116773 36415 116807
rect 36357 116767 36415 116773
rect 24302 116736 24308 116748
rect 23431 116708 24164 116736
rect 24263 116708 24308 116736
rect 23431 116705 23443 116708
rect 23385 116699 23443 116705
rect 24302 116696 24308 116708
rect 24360 116696 24366 116748
rect 25041 116739 25099 116745
rect 25041 116705 25053 116739
rect 25087 116736 25099 116739
rect 25590 116736 25596 116748
rect 25087 116708 25596 116736
rect 25087 116705 25099 116708
rect 25041 116699 25099 116705
rect 25590 116696 25596 116708
rect 25648 116696 25654 116748
rect 25774 116736 25780 116748
rect 25735 116708 25780 116736
rect 25774 116696 25780 116708
rect 25832 116696 25838 116748
rect 26510 116736 26516 116748
rect 26471 116708 26516 116736
rect 26510 116696 26516 116708
rect 26568 116696 26574 116748
rect 27893 116739 27951 116745
rect 27893 116705 27905 116739
rect 27939 116705 27951 116739
rect 27893 116699 27951 116705
rect 28629 116739 28687 116745
rect 28629 116705 28641 116739
rect 28675 116705 28687 116739
rect 28629 116699 28687 116705
rect 29273 116739 29331 116745
rect 29273 116705 29285 116739
rect 29319 116736 29331 116739
rect 30190 116736 30196 116748
rect 29319 116708 30196 116736
rect 29319 116705 29331 116708
rect 29273 116699 29331 116705
rect 3878 116628 3884 116680
rect 3936 116668 3942 116680
rect 5721 116671 5779 116677
rect 5721 116668 5733 116671
rect 3936 116640 5733 116668
rect 3936 116628 3942 116640
rect 5721 116637 5733 116640
rect 5767 116637 5779 116671
rect 5721 116631 5779 116637
rect 14642 116628 14648 116680
rect 14700 116668 14706 116680
rect 16298 116668 16304 116680
rect 14700 116640 16304 116668
rect 14700 116628 14706 116640
rect 16298 116628 16304 116640
rect 16356 116628 16362 116680
rect 17218 116628 17224 116680
rect 17276 116668 17282 116680
rect 19058 116668 19064 116680
rect 17276 116640 19064 116668
rect 17276 116628 17282 116640
rect 19058 116628 19064 116640
rect 19116 116628 19122 116680
rect 20070 116628 20076 116680
rect 20128 116668 20134 116680
rect 22002 116668 22008 116680
rect 20128 116640 22008 116668
rect 20128 116628 20134 116640
rect 22002 116628 22008 116640
rect 22060 116628 22066 116680
rect 22094 116628 22100 116680
rect 22152 116668 22158 116680
rect 27908 116668 27936 116699
rect 22152 116640 27936 116668
rect 22152 116628 22158 116640
rect 6546 116600 6552 116612
rect 1872 116572 6552 116600
rect 6546 116560 6552 116572
rect 6604 116560 6610 116612
rect 17954 116560 17960 116612
rect 18012 116600 18018 116612
rect 21726 116600 21732 116612
rect 18012 116572 21732 116600
rect 18012 116560 18018 116572
rect 21726 116560 21732 116572
rect 21784 116560 21790 116612
rect 21818 116560 21824 116612
rect 21876 116600 21882 116612
rect 28644 116600 28672 116699
rect 30190 116696 30196 116708
rect 30248 116696 30254 116748
rect 30929 116739 30987 116745
rect 30929 116705 30941 116739
rect 30975 116736 30987 116739
rect 31662 116736 31668 116748
rect 30975 116708 31668 116736
rect 30975 116705 30987 116708
rect 30929 116699 30987 116705
rect 31662 116696 31668 116708
rect 31720 116696 31726 116748
rect 32766 116696 32772 116748
rect 32824 116736 32830 116748
rect 33229 116739 33287 116745
rect 33229 116736 33241 116739
rect 32824 116708 33241 116736
rect 32824 116696 32830 116708
rect 33229 116705 33241 116708
rect 33275 116705 33287 116739
rect 33229 116699 33287 116705
rect 33965 116739 34023 116745
rect 33965 116705 33977 116739
rect 34011 116705 34023 116739
rect 34698 116736 34704 116748
rect 34659 116708 34704 116736
rect 33965 116699 34023 116705
rect 29638 116668 29644 116680
rect 29599 116640 29644 116668
rect 29638 116628 29644 116640
rect 29696 116628 29702 116680
rect 31018 116628 31024 116680
rect 31076 116668 31082 116680
rect 31297 116671 31355 116677
rect 31297 116668 31309 116671
rect 31076 116640 31309 116668
rect 31076 116628 31082 116640
rect 31297 116637 31309 116640
rect 31343 116637 31355 116671
rect 31297 116631 31355 116637
rect 33410 116628 33416 116680
rect 33468 116668 33474 116680
rect 33980 116668 34008 116699
rect 34698 116696 34704 116708
rect 34756 116696 34762 116748
rect 35437 116739 35495 116745
rect 35437 116705 35449 116739
rect 35483 116705 35495 116739
rect 35437 116699 35495 116705
rect 33468 116640 34008 116668
rect 33468 116628 33474 116640
rect 34606 116628 34612 116680
rect 34664 116668 34670 116680
rect 35452 116668 35480 116699
rect 35894 116696 35900 116748
rect 35952 116736 35958 116748
rect 36173 116739 36231 116745
rect 36173 116736 36185 116739
rect 35952 116708 36185 116736
rect 35952 116696 35958 116708
rect 36173 116705 36185 116708
rect 36219 116705 36231 116739
rect 36173 116699 36231 116705
rect 36909 116739 36967 116745
rect 36909 116705 36921 116739
rect 36955 116705 36967 116739
rect 36909 116699 36967 116705
rect 34664 116640 35480 116668
rect 34664 116628 34670 116640
rect 35526 116628 35532 116680
rect 35584 116668 35590 116680
rect 36924 116668 36952 116699
rect 35584 116640 36952 116668
rect 35584 116628 35590 116640
rect 21876 116572 28672 116600
rect 21876 116560 21882 116572
rect 28810 116560 28816 116612
rect 28868 116600 28874 116612
rect 29733 116603 29791 116609
rect 29733 116600 29745 116603
rect 28868 116572 29745 116600
rect 28868 116560 28874 116572
rect 29733 116569 29745 116572
rect 29779 116569 29791 116603
rect 29733 116563 29791 116569
rect 34149 116603 34207 116609
rect 34149 116569 34161 116603
rect 34195 116600 34207 116603
rect 38838 116600 38844 116612
rect 34195 116572 38844 116600
rect 34195 116569 34207 116572
rect 34149 116563 34207 116569
rect 38838 116560 38844 116572
rect 38896 116560 38902 116612
rect 3418 116532 3424 116544
rect 3379 116504 3424 116532
rect 3418 116492 3424 116504
rect 3476 116492 3482 116544
rect 7650 116492 7656 116544
rect 7708 116532 7714 116544
rect 8481 116535 8539 116541
rect 8481 116532 8493 116535
rect 7708 116504 8493 116532
rect 7708 116492 7714 116504
rect 8481 116501 8493 116504
rect 8527 116501 8539 116535
rect 8481 116495 8539 116501
rect 21082 116492 21088 116544
rect 21140 116532 21146 116544
rect 22370 116532 22376 116544
rect 21140 116504 22376 116532
rect 21140 116492 21146 116504
rect 22370 116492 22376 116504
rect 22428 116492 22434 116544
rect 22462 116492 22468 116544
rect 22520 116532 22526 116544
rect 23477 116535 23535 116541
rect 23477 116532 23489 116535
rect 22520 116504 23489 116532
rect 22520 116492 22526 116504
rect 23477 116501 23489 116504
rect 23523 116501 23535 116535
rect 23477 116495 23535 116501
rect 25038 116492 25044 116544
rect 25096 116532 25102 116544
rect 25869 116535 25927 116541
rect 25869 116532 25881 116535
rect 25096 116504 25881 116532
rect 25096 116492 25102 116504
rect 25869 116501 25881 116504
rect 25915 116501 25927 116535
rect 25869 116495 25927 116501
rect 29362 116492 29368 116544
rect 29420 116541 29426 116544
rect 29420 116535 29469 116541
rect 29420 116501 29423 116535
rect 29457 116501 29469 116535
rect 29546 116532 29552 116544
rect 29507 116504 29552 116532
rect 29420 116495 29469 116501
rect 29420 116492 29426 116495
rect 29546 116492 29552 116504
rect 29604 116492 29610 116544
rect 30926 116492 30932 116544
rect 30984 116532 30990 116544
rect 31067 116535 31125 116541
rect 31067 116532 31079 116535
rect 30984 116504 31079 116532
rect 30984 116492 30990 116504
rect 31067 116501 31079 116504
rect 31113 116501 31125 116535
rect 31202 116532 31208 116544
rect 31163 116504 31208 116532
rect 31067 116495 31125 116501
rect 31202 116492 31208 116504
rect 31260 116492 31266 116544
rect 33134 116492 33140 116544
rect 33192 116532 33198 116544
rect 33594 116532 33600 116544
rect 33192 116504 33600 116532
rect 33192 116492 33198 116504
rect 33594 116492 33600 116504
rect 33652 116492 33658 116544
rect 35434 116492 35440 116544
rect 35492 116532 35498 116544
rect 37001 116535 37059 116541
rect 37001 116532 37013 116535
rect 35492 116504 37013 116532
rect 35492 116492 35498 116504
rect 37001 116501 37013 116504
rect 37047 116501 37059 116535
rect 37001 116495 37059 116501
rect 1104 116442 38824 116464
rect 1104 116390 4246 116442
rect 4298 116390 4310 116442
rect 4362 116390 4374 116442
rect 4426 116390 4438 116442
rect 4490 116390 34966 116442
rect 35018 116390 35030 116442
rect 35082 116390 35094 116442
rect 35146 116390 35158 116442
rect 35210 116390 38824 116442
rect 1104 116368 38824 116390
rect 2222 116288 2228 116340
rect 2280 116328 2286 116340
rect 2409 116331 2467 116337
rect 2409 116328 2421 116331
rect 2280 116300 2421 116328
rect 2280 116288 2286 116300
rect 2409 116297 2421 116300
rect 2455 116297 2467 116331
rect 2409 116291 2467 116297
rect 2774 116288 2780 116340
rect 2832 116328 2838 116340
rect 3145 116331 3203 116337
rect 3145 116328 3157 116331
rect 2832 116300 3157 116328
rect 2832 116288 2838 116300
rect 3145 116297 3157 116300
rect 3191 116297 3203 116331
rect 3145 116291 3203 116297
rect 4614 116288 4620 116340
rect 4672 116328 4678 116340
rect 5629 116331 5687 116337
rect 5629 116328 5641 116331
rect 4672 116300 5641 116328
rect 4672 116288 4678 116300
rect 5629 116297 5641 116300
rect 5675 116297 5687 116331
rect 5629 116291 5687 116297
rect 5810 116288 5816 116340
rect 5868 116328 5874 116340
rect 6365 116331 6423 116337
rect 6365 116328 6377 116331
rect 5868 116300 6377 116328
rect 5868 116288 5874 116300
rect 6365 116297 6377 116300
rect 6411 116297 6423 116331
rect 6365 116291 6423 116297
rect 6638 116288 6644 116340
rect 6696 116328 6702 116340
rect 7837 116331 7895 116337
rect 7837 116328 7849 116331
rect 6696 116300 7849 116328
rect 6696 116288 6702 116300
rect 7837 116297 7849 116300
rect 7883 116297 7895 116331
rect 7837 116291 7895 116297
rect 10410 116288 10416 116340
rect 10468 116328 10474 116340
rect 10597 116331 10655 116337
rect 10597 116328 10609 116331
rect 10468 116300 10609 116328
rect 10468 116288 10474 116300
rect 10597 116297 10609 116300
rect 10643 116297 10655 116331
rect 10597 116291 10655 116297
rect 11054 116288 11060 116340
rect 11112 116328 11118 116340
rect 11333 116331 11391 116337
rect 11333 116328 11345 116331
rect 11112 116300 11345 116328
rect 11112 116288 11118 116300
rect 11333 116297 11345 116300
rect 11379 116297 11391 116331
rect 11333 116291 11391 116297
rect 15654 116288 15660 116340
rect 15712 116328 15718 116340
rect 15749 116331 15807 116337
rect 15749 116328 15761 116331
rect 15712 116300 15761 116328
rect 15712 116288 15718 116300
rect 15749 116297 15761 116300
rect 15795 116297 15807 116331
rect 15749 116291 15807 116297
rect 19978 116288 19984 116340
rect 20036 116328 20042 116340
rect 20165 116331 20223 116337
rect 20165 116328 20177 116331
rect 20036 116300 20177 116328
rect 20036 116288 20042 116300
rect 20165 116297 20177 116300
rect 20211 116297 20223 116331
rect 20165 116291 20223 116297
rect 21266 116288 21272 116340
rect 21324 116328 21330 116340
rect 21453 116331 21511 116337
rect 21453 116328 21465 116331
rect 21324 116300 21465 116328
rect 21324 116288 21330 116300
rect 21453 116297 21465 116300
rect 21499 116297 21511 116331
rect 21453 116291 21511 116297
rect 22094 116288 22100 116340
rect 22152 116328 22158 116340
rect 22189 116331 22247 116337
rect 22189 116328 22201 116331
rect 22152 116300 22201 116328
rect 22152 116288 22158 116300
rect 22189 116297 22201 116300
rect 22235 116297 22247 116331
rect 22189 116291 22247 116297
rect 22646 116288 22652 116340
rect 22704 116328 22710 116340
rect 22922 116328 22928 116340
rect 22704 116300 22928 116328
rect 22704 116288 22710 116300
rect 22922 116288 22928 116300
rect 22980 116288 22986 116340
rect 23106 116288 23112 116340
rect 23164 116328 23170 116340
rect 23293 116331 23351 116337
rect 23293 116328 23305 116331
rect 23164 116300 23305 116328
rect 23164 116288 23170 116300
rect 23293 116297 23305 116300
rect 23339 116297 23351 116331
rect 23293 116291 23351 116297
rect 23750 116288 23756 116340
rect 23808 116328 23814 116340
rect 24029 116331 24087 116337
rect 24029 116328 24041 116331
rect 23808 116300 24041 116328
rect 23808 116288 23814 116300
rect 24029 116297 24041 116300
rect 24075 116297 24087 116331
rect 24029 116291 24087 116297
rect 25866 116288 25872 116340
rect 25924 116328 25930 116340
rect 26053 116331 26111 116337
rect 26053 116328 26065 116331
rect 25924 116300 26065 116328
rect 25924 116288 25930 116300
rect 26053 116297 26065 116300
rect 26099 116297 26111 116331
rect 26053 116291 26111 116297
rect 26602 116288 26608 116340
rect 26660 116328 26666 116340
rect 27617 116331 27675 116337
rect 27617 116328 27629 116331
rect 26660 116300 27629 116328
rect 26660 116288 26666 116300
rect 27617 116297 27629 116300
rect 27663 116297 27675 116331
rect 27617 116291 27675 116297
rect 28166 116288 28172 116340
rect 28224 116328 28230 116340
rect 33321 116331 33379 116337
rect 33321 116328 33333 116331
rect 28224 116300 33333 116328
rect 28224 116288 28230 116300
rect 33321 116297 33333 116300
rect 33367 116297 33379 116331
rect 33321 116291 33379 116297
rect 35250 116288 35256 116340
rect 35308 116328 35314 116340
rect 35897 116331 35955 116337
rect 35897 116328 35909 116331
rect 35308 116300 35909 116328
rect 35308 116288 35314 116300
rect 35897 116297 35909 116300
rect 35943 116297 35955 116331
rect 35897 116291 35955 116297
rect 1854 116220 1860 116272
rect 1912 116260 1918 116272
rect 4985 116263 5043 116269
rect 1912 116232 4936 116260
rect 1912 116220 1918 116232
rect 3602 116152 3608 116204
rect 3660 116192 3666 116204
rect 4522 116192 4528 116204
rect 3660 116164 4528 116192
rect 3660 116152 3666 116164
rect 4522 116152 4528 116164
rect 4580 116152 4586 116204
rect 4908 116124 4936 116232
rect 4985 116229 4997 116263
rect 5031 116260 5043 116263
rect 5166 116260 5172 116272
rect 5031 116232 5172 116260
rect 5031 116229 5043 116232
rect 4985 116223 5043 116229
rect 5166 116220 5172 116232
rect 5224 116220 5230 116272
rect 5994 116220 6000 116272
rect 6052 116260 6058 116272
rect 7193 116263 7251 116269
rect 7193 116260 7205 116263
rect 6052 116232 7205 116260
rect 6052 116220 6058 116232
rect 7193 116229 7205 116232
rect 7239 116229 7251 116263
rect 7193 116223 7251 116229
rect 16114 116220 16120 116272
rect 16172 116260 16178 116272
rect 16577 116263 16635 116269
rect 16577 116260 16589 116263
rect 16172 116232 16589 116260
rect 16172 116220 16178 116232
rect 16577 116229 16589 116232
rect 16623 116229 16635 116263
rect 21358 116260 21364 116272
rect 16577 116223 16635 116229
rect 19996 116232 21364 116260
rect 9490 116192 9496 116204
rect 9451 116164 9496 116192
rect 9490 116152 9496 116164
rect 9548 116152 9554 116204
rect 11885 116195 11943 116201
rect 11885 116161 11897 116195
rect 11931 116192 11943 116195
rect 13078 116192 13084 116204
rect 11931 116164 13084 116192
rect 11931 116161 11943 116164
rect 11885 116155 11943 116161
rect 13078 116152 13084 116164
rect 13136 116152 13142 116204
rect 13173 116195 13231 116201
rect 13173 116161 13185 116195
rect 13219 116192 13231 116195
rect 15010 116192 15016 116204
rect 13219 116164 15016 116192
rect 13219 116161 13231 116164
rect 13173 116155 13231 116161
rect 15010 116152 15016 116164
rect 15068 116152 15074 116204
rect 17037 116195 17095 116201
rect 17037 116161 17049 116195
rect 17083 116192 17095 116195
rect 19886 116192 19892 116204
rect 17083 116164 19892 116192
rect 17083 116161 17095 116164
rect 17037 116155 17095 116161
rect 19886 116152 19892 116164
rect 19944 116152 19950 116204
rect 5166 116124 5172 116136
rect 4908 116096 5172 116124
rect 5166 116084 5172 116096
rect 5224 116084 5230 116136
rect 12529 116127 12587 116133
rect 12529 116093 12541 116127
rect 12575 116124 12587 116127
rect 13814 116124 13820 116136
rect 12575 116096 13820 116124
rect 12575 116093 12587 116096
rect 12529 116087 12587 116093
rect 13814 116084 13820 116096
rect 13872 116084 13878 116136
rect 14737 116127 14795 116133
rect 14737 116093 14749 116127
rect 14783 116124 14795 116127
rect 15930 116124 15936 116136
rect 14783 116096 15936 116124
rect 14783 116093 14795 116096
rect 14737 116087 14795 116093
rect 15930 116084 15936 116096
rect 15988 116084 15994 116136
rect 18325 116127 18383 116133
rect 18325 116093 18337 116127
rect 18371 116124 18383 116127
rect 19996 116124 20024 116232
rect 21358 116220 21364 116232
rect 21416 116220 21422 116272
rect 22370 116220 22376 116272
rect 22428 116260 22434 116272
rect 24762 116260 24768 116272
rect 22428 116232 24768 116260
rect 22428 116220 22434 116232
rect 24762 116220 24768 116232
rect 24820 116220 24826 116272
rect 25409 116263 25467 116269
rect 25409 116229 25421 116263
rect 25455 116260 25467 116263
rect 26694 116260 26700 116272
rect 25455 116232 26700 116260
rect 25455 116229 25467 116232
rect 25409 116223 25467 116229
rect 26694 116220 26700 116232
rect 26752 116220 26758 116272
rect 26970 116220 26976 116272
rect 27028 116260 27034 116272
rect 28445 116263 28503 116269
rect 28445 116260 28457 116263
rect 27028 116232 28457 116260
rect 27028 116220 27034 116232
rect 28445 116229 28457 116232
rect 28491 116229 28503 116263
rect 30742 116260 30748 116272
rect 30703 116232 30748 116260
rect 28445 116223 28503 116229
rect 30742 116220 30748 116232
rect 30800 116220 30806 116272
rect 31478 116260 31484 116272
rect 30852 116232 31484 116260
rect 23106 116192 23112 116204
rect 20088 116164 23112 116192
rect 20088 116133 20116 116164
rect 23106 116152 23112 116164
rect 23164 116152 23170 116204
rect 26234 116192 26240 116204
rect 23216 116164 26240 116192
rect 23216 116133 23244 116164
rect 26234 116152 26240 116164
rect 26292 116152 26298 116204
rect 28810 116192 28816 116204
rect 26620 116164 28816 116192
rect 18371 116096 20024 116124
rect 20073 116127 20131 116133
rect 18371 116093 18383 116096
rect 18325 116087 18383 116093
rect 20073 116093 20085 116127
rect 20119 116093 20131 116127
rect 20073 116087 20131 116093
rect 22097 116127 22155 116133
rect 22097 116093 22109 116127
rect 22143 116124 22155 116127
rect 23201 116127 23259 116133
rect 22143 116096 23152 116124
rect 22143 116093 22155 116096
rect 22097 116087 22155 116093
rect 2314 116056 2320 116068
rect 2275 116028 2320 116056
rect 2314 116016 2320 116028
rect 2372 116016 2378 116068
rect 3050 116056 3056 116068
rect 3011 116028 3056 116056
rect 3050 116016 3056 116028
rect 3108 116016 3114 116068
rect 4801 116059 4859 116065
rect 4801 116025 4813 116059
rect 4847 116056 4859 116059
rect 5442 116056 5448 116068
rect 4847 116028 5448 116056
rect 4847 116025 4859 116028
rect 4801 116019 4859 116025
rect 5442 116016 5448 116028
rect 5500 116016 5506 116068
rect 5537 116059 5595 116065
rect 5537 116025 5549 116059
rect 5583 116056 5595 116059
rect 5718 116056 5724 116068
rect 5583 116028 5724 116056
rect 5583 116025 5595 116028
rect 5537 116019 5595 116025
rect 5718 116016 5724 116028
rect 5776 116016 5782 116068
rect 6270 116056 6276 116068
rect 6231 116028 6276 116056
rect 6270 116016 6276 116028
rect 6328 116016 6334 116068
rect 7009 116059 7067 116065
rect 7009 116025 7021 116059
rect 7055 116056 7067 116059
rect 7558 116056 7564 116068
rect 7055 116028 7564 116056
rect 7055 116025 7067 116028
rect 7009 116019 7067 116025
rect 7558 116016 7564 116028
rect 7616 116016 7622 116068
rect 7742 116056 7748 116068
rect 7703 116028 7748 116056
rect 7742 116016 7748 116028
rect 7800 116016 7806 116068
rect 10505 116059 10563 116065
rect 10505 116025 10517 116059
rect 10551 116056 10563 116059
rect 10962 116056 10968 116068
rect 10551 116028 10968 116056
rect 10551 116025 10563 116028
rect 10505 116019 10563 116025
rect 10962 116016 10968 116028
rect 11020 116016 11026 116068
rect 11238 116056 11244 116068
rect 11199 116028 11244 116056
rect 11238 116016 11244 116028
rect 11296 116016 11302 116068
rect 15654 116056 15660 116068
rect 15615 116028 15660 116056
rect 15654 116016 15660 116028
rect 15712 116016 15718 116068
rect 16390 116056 16396 116068
rect 16351 116028 16396 116056
rect 16390 116016 16396 116028
rect 16448 116016 16454 116068
rect 17681 116059 17739 116065
rect 17681 116025 17693 116059
rect 17727 116056 17739 116059
rect 20530 116056 20536 116068
rect 17727 116028 20536 116056
rect 17727 116025 17739 116028
rect 17681 116019 17739 116025
rect 20530 116016 20536 116028
rect 20588 116016 20594 116068
rect 21361 116059 21419 116065
rect 21361 116025 21373 116059
rect 21407 116056 21419 116059
rect 23014 116056 23020 116068
rect 21407 116028 23020 116056
rect 21407 116025 21419 116028
rect 21361 116019 21419 116025
rect 23014 116016 23020 116028
rect 23072 116016 23078 116068
rect 23124 116056 23152 116096
rect 23201 116093 23213 116127
rect 23247 116093 23259 116127
rect 25314 116124 25320 116136
rect 23201 116087 23259 116093
rect 23860 116096 25320 116124
rect 23860 116056 23888 116096
rect 25314 116084 25320 116096
rect 25372 116084 25378 116136
rect 26620 116133 26648 116164
rect 28810 116152 28816 116164
rect 28868 116152 28874 116204
rect 30558 116152 30564 116204
rect 30616 116201 30622 116204
rect 30852 116201 30880 116232
rect 31478 116220 31484 116232
rect 31536 116220 31542 116272
rect 31938 116260 31944 116272
rect 31899 116232 31944 116260
rect 31938 116220 31944 116232
rect 31996 116220 32002 116272
rect 33134 116260 33140 116272
rect 33095 116232 33140 116260
rect 33134 116220 33140 116232
rect 33192 116220 33198 116272
rect 35710 116220 35716 116272
rect 35768 116260 35774 116272
rect 36725 116263 36783 116269
rect 36725 116260 36737 116263
rect 35768 116232 36737 116260
rect 35768 116220 35774 116232
rect 36725 116229 36737 116232
rect 36771 116229 36783 116263
rect 38194 116260 38200 116272
rect 36725 116223 36783 116229
rect 36832 116232 38200 116260
rect 30616 116195 30674 116201
rect 30616 116161 30628 116195
rect 30662 116161 30674 116195
rect 30616 116155 30674 116161
rect 30837 116195 30895 116201
rect 30837 116161 30849 116195
rect 30883 116161 30895 116195
rect 30837 116155 30895 116161
rect 30929 116195 30987 116201
rect 30929 116161 30941 116195
rect 30975 116161 30987 116195
rect 30929 116155 30987 116161
rect 30616 116152 30622 116155
rect 26605 116127 26663 116133
rect 26605 116093 26617 116127
rect 26651 116093 26663 116127
rect 26605 116087 26663 116093
rect 26789 116127 26847 116133
rect 26789 116093 26801 116127
rect 26835 116124 26847 116127
rect 30944 116124 30972 116155
rect 31110 116152 31116 116204
rect 31168 116192 31174 116204
rect 32033 116195 32091 116201
rect 32033 116192 32045 116195
rect 31168 116164 32045 116192
rect 31168 116152 31174 116164
rect 32033 116161 32045 116164
rect 32079 116161 32091 116195
rect 32033 116155 32091 116161
rect 33229 116195 33287 116201
rect 33229 116161 33241 116195
rect 33275 116192 33287 116195
rect 33870 116192 33876 116204
rect 33275 116164 33876 116192
rect 33275 116161 33287 116164
rect 33229 116155 33287 116161
rect 33870 116152 33876 116164
rect 33928 116152 33934 116204
rect 34793 116195 34851 116201
rect 34793 116161 34805 116195
rect 34839 116192 34851 116195
rect 36832 116192 36860 116232
rect 38194 116220 38200 116232
rect 38252 116220 38258 116272
rect 37826 116192 37832 116204
rect 34839 116164 36860 116192
rect 37787 116164 37832 116192
rect 34839 116161 34851 116164
rect 34793 116155 34851 116161
rect 37826 116152 37832 116164
rect 37884 116152 37890 116204
rect 26835 116096 30972 116124
rect 31812 116127 31870 116133
rect 26835 116093 26847 116096
rect 26789 116087 26847 116093
rect 31812 116093 31824 116127
rect 31858 116124 31870 116127
rect 32122 116124 32128 116136
rect 31858 116096 32128 116124
rect 31858 116093 31870 116096
rect 31812 116087 31870 116093
rect 32122 116084 32128 116096
rect 32180 116084 32186 116136
rect 32398 116084 32404 116136
rect 32456 116124 32462 116136
rect 33008 116127 33066 116133
rect 33008 116124 33020 116127
rect 32456 116096 33020 116124
rect 32456 116084 32462 116096
rect 33008 116093 33020 116096
rect 33054 116093 33066 116127
rect 33008 116087 33066 116093
rect 35710 116084 35716 116136
rect 35768 116124 35774 116136
rect 36541 116127 36599 116133
rect 36541 116124 36553 116127
rect 35768 116096 36553 116124
rect 35768 116084 35774 116096
rect 36541 116093 36553 116096
rect 36587 116093 36599 116127
rect 37642 116124 37648 116136
rect 37603 116096 37648 116124
rect 36541 116087 36599 116093
rect 37642 116084 37648 116096
rect 37700 116084 37706 116136
rect 23124 116028 23888 116056
rect 23937 116059 23995 116065
rect 23937 116025 23949 116059
rect 23983 116056 23995 116059
rect 25866 116056 25872 116068
rect 23983 116028 25872 116056
rect 23983 116025 23995 116028
rect 23937 116019 23995 116025
rect 25866 116016 25872 116028
rect 25924 116016 25930 116068
rect 25961 116059 26019 116065
rect 25961 116025 25973 116059
rect 26007 116025 26019 116059
rect 25961 116019 26019 116025
rect 5074 115948 5080 116000
rect 5132 115988 5138 116000
rect 5626 115988 5632 116000
rect 5132 115960 5632 115988
rect 5132 115948 5138 115960
rect 5626 115948 5632 115960
rect 5684 115948 5690 116000
rect 20714 115948 20720 116000
rect 20772 115988 20778 116000
rect 25976 115988 26004 116019
rect 26142 116016 26148 116068
rect 26200 116056 26206 116068
rect 26973 116059 27031 116065
rect 26973 116056 26985 116059
rect 26200 116028 26985 116056
rect 26200 116016 26206 116028
rect 26973 116025 26985 116028
rect 27019 116025 27031 116059
rect 27522 116056 27528 116068
rect 27483 116028 27528 116056
rect 26973 116019 27031 116025
rect 27522 116016 27528 116028
rect 27580 116016 27586 116068
rect 28258 116056 28264 116068
rect 28219 116028 28264 116056
rect 28258 116016 28264 116028
rect 28316 116016 28322 116068
rect 28994 116056 29000 116068
rect 28955 116028 29000 116056
rect 28994 116016 29000 116028
rect 29052 116016 29058 116068
rect 30469 116059 30527 116065
rect 30469 116025 30481 116059
rect 30515 116056 30527 116059
rect 30650 116056 30656 116068
rect 30515 116028 30656 116056
rect 30515 116025 30527 116028
rect 30469 116019 30527 116025
rect 30650 116016 30656 116028
rect 30708 116016 30714 116068
rect 31665 116059 31723 116065
rect 31665 116025 31677 116059
rect 31711 116056 31723 116059
rect 32674 116056 32680 116068
rect 31711 116028 32680 116056
rect 31711 116025 31723 116028
rect 31665 116019 31723 116025
rect 32674 116016 32680 116028
rect 32732 116016 32738 116068
rect 32858 116056 32864 116068
rect 32819 116028 32864 116056
rect 32858 116016 32864 116028
rect 32916 116016 32922 116068
rect 34054 116016 34060 116068
rect 34112 116056 34118 116068
rect 34609 116059 34667 116065
rect 34609 116056 34621 116059
rect 34112 116028 34621 116056
rect 34112 116016 34118 116028
rect 34609 116025 34621 116028
rect 34655 116025 34667 116059
rect 34609 116019 34667 116025
rect 35250 116016 35256 116068
rect 35308 116056 35314 116068
rect 35805 116059 35863 116065
rect 35805 116056 35817 116059
rect 35308 116028 35817 116056
rect 35308 116016 35314 116028
rect 35805 116025 35817 116028
rect 35851 116025 35863 116059
rect 35805 116019 35863 116025
rect 20772 115960 26004 115988
rect 20772 115948 20778 115960
rect 27338 115948 27344 116000
rect 27396 115988 27402 116000
rect 29089 115991 29147 115997
rect 29089 115988 29101 115991
rect 27396 115960 29101 115988
rect 27396 115948 27402 115960
rect 29089 115957 29101 115960
rect 29135 115957 29147 115991
rect 29089 115951 29147 115957
rect 29822 115948 29828 116000
rect 29880 115988 29886 116000
rect 32309 115991 32367 115997
rect 32309 115988 32321 115991
rect 29880 115960 32321 115988
rect 29880 115948 29886 115960
rect 32309 115957 32321 115960
rect 32355 115957 32367 115991
rect 32309 115951 32367 115957
rect 1104 115898 38824 115920
rect 1104 115846 19606 115898
rect 19658 115846 19670 115898
rect 19722 115846 19734 115898
rect 19786 115846 19798 115898
rect 19850 115846 38824 115898
rect 1104 115824 38824 115846
rect 1670 115744 1676 115796
rect 1728 115784 1734 115796
rect 2406 115784 2412 115796
rect 1728 115756 2412 115784
rect 1728 115744 1734 115756
rect 2406 115744 2412 115756
rect 2464 115744 2470 115796
rect 3418 115784 3424 115796
rect 2700 115756 3424 115784
rect 474 115676 480 115728
rect 532 115716 538 115728
rect 2700 115716 2728 115756
rect 3418 115744 3424 115756
rect 3476 115744 3482 115796
rect 3510 115744 3516 115796
rect 3568 115784 3574 115796
rect 4433 115787 4491 115793
rect 4433 115784 4445 115787
rect 3568 115756 4445 115784
rect 3568 115744 3574 115756
rect 4433 115753 4445 115756
rect 4479 115753 4491 115787
rect 4433 115747 4491 115753
rect 4706 115744 4712 115796
rect 4764 115784 4770 115796
rect 5169 115787 5227 115793
rect 5169 115784 5181 115787
rect 4764 115756 5181 115784
rect 4764 115744 4770 115756
rect 5169 115753 5181 115756
rect 5215 115753 5227 115787
rect 5169 115747 5227 115753
rect 7282 115744 7288 115796
rect 7340 115784 7346 115796
rect 8297 115787 8355 115793
rect 8297 115784 8309 115787
rect 7340 115756 8309 115784
rect 7340 115744 7346 115756
rect 8297 115753 8309 115756
rect 8343 115753 8355 115787
rect 8297 115747 8355 115753
rect 8386 115744 8392 115796
rect 8444 115784 8450 115796
rect 8849 115787 8907 115793
rect 8849 115784 8861 115787
rect 8444 115756 8861 115784
rect 8444 115744 8450 115756
rect 8849 115753 8861 115756
rect 8895 115753 8907 115787
rect 8849 115747 8907 115753
rect 9493 115787 9551 115793
rect 9493 115753 9505 115787
rect 9539 115784 9551 115787
rect 9766 115784 9772 115796
rect 9539 115756 9772 115784
rect 9539 115753 9551 115756
rect 9493 115747 9551 115753
rect 9766 115744 9772 115756
rect 9824 115744 9830 115796
rect 10137 115787 10195 115793
rect 10137 115753 10149 115787
rect 10183 115784 10195 115787
rect 11146 115784 11152 115796
rect 10183 115756 11152 115784
rect 10183 115753 10195 115756
rect 10137 115747 10195 115753
rect 11146 115744 11152 115756
rect 11204 115744 11210 115796
rect 13357 115787 13415 115793
rect 13357 115753 13369 115787
rect 13403 115784 13415 115787
rect 14090 115784 14096 115796
rect 13403 115756 14096 115784
rect 13403 115753 13415 115756
rect 13357 115747 13415 115753
rect 14090 115744 14096 115756
rect 14148 115744 14154 115796
rect 14553 115787 14611 115793
rect 14553 115753 14565 115787
rect 14599 115784 14611 115787
rect 15838 115784 15844 115796
rect 14599 115756 15844 115784
rect 14599 115753 14611 115756
rect 14553 115747 14611 115753
rect 15838 115744 15844 115756
rect 15896 115744 15902 115796
rect 18417 115787 18475 115793
rect 18417 115753 18429 115787
rect 18463 115784 18475 115787
rect 20070 115784 20076 115796
rect 18463 115756 20076 115784
rect 18463 115753 18475 115756
rect 18417 115747 18475 115753
rect 20070 115744 20076 115756
rect 20128 115744 20134 115796
rect 23290 115784 23296 115796
rect 21284 115756 23296 115784
rect 532 115688 2728 115716
rect 2777 115719 2835 115725
rect 532 115676 538 115688
rect 2777 115685 2789 115719
rect 2823 115716 2835 115719
rect 2958 115716 2964 115728
rect 2823 115688 2964 115716
rect 2823 115685 2835 115688
rect 2777 115679 2835 115685
rect 2958 115676 2964 115688
rect 3016 115676 3022 115728
rect 3789 115719 3847 115725
rect 3436 115688 3740 115716
rect 1857 115651 1915 115657
rect 1857 115617 1869 115651
rect 1903 115648 1915 115651
rect 2498 115648 2504 115660
rect 1903 115620 2504 115648
rect 1903 115617 1915 115620
rect 1857 115611 1915 115617
rect 2498 115608 2504 115620
rect 2556 115608 2562 115660
rect 2593 115651 2651 115657
rect 2593 115617 2605 115651
rect 2639 115648 2651 115651
rect 3436 115648 3464 115688
rect 3602 115648 3608 115660
rect 2639 115620 3464 115648
rect 3563 115620 3608 115648
rect 2639 115617 2651 115620
rect 2593 115611 2651 115617
rect 3602 115608 3608 115620
rect 3660 115608 3666 115660
rect 3712 115648 3740 115688
rect 3789 115685 3801 115719
rect 3835 115716 3847 115719
rect 3970 115716 3976 115728
rect 3835 115688 3976 115716
rect 3835 115685 3847 115688
rect 3789 115679 3847 115685
rect 3970 115676 3976 115688
rect 4028 115676 4034 115728
rect 8662 115716 8668 115728
rect 4264 115688 8668 115716
rect 4264 115648 4292 115688
rect 8662 115676 8668 115688
rect 8720 115676 8726 115728
rect 10781 115719 10839 115725
rect 10781 115685 10793 115719
rect 10827 115716 10839 115719
rect 11330 115716 11336 115728
rect 10827 115688 11336 115716
rect 10827 115685 10839 115688
rect 10781 115679 10839 115685
rect 11330 115676 11336 115688
rect 11388 115676 11394 115728
rect 15197 115719 15255 115725
rect 15197 115685 15209 115719
rect 15243 115716 15255 115719
rect 16574 115716 16580 115728
rect 15243 115688 16580 115716
rect 15243 115685 15255 115688
rect 15197 115679 15255 115685
rect 16574 115676 16580 115688
rect 16632 115676 16638 115728
rect 19061 115719 19119 115725
rect 19061 115685 19073 115719
rect 19107 115716 19119 115719
rect 21284 115716 21312 115756
rect 23290 115744 23296 115756
rect 23348 115744 23354 115796
rect 23566 115744 23572 115796
rect 23624 115784 23630 115796
rect 24670 115784 24676 115796
rect 23624 115756 24676 115784
rect 23624 115744 23630 115756
rect 24670 115744 24676 115756
rect 24728 115744 24734 115796
rect 25958 115784 25964 115796
rect 24780 115756 25964 115784
rect 24780 115716 24808 115756
rect 25958 115744 25964 115756
rect 26016 115744 26022 115796
rect 26326 115744 26332 115796
rect 26384 115784 26390 115796
rect 26513 115787 26571 115793
rect 26513 115784 26525 115787
rect 26384 115756 26525 115784
rect 26384 115744 26390 115756
rect 26513 115753 26525 115756
rect 26559 115753 26571 115787
rect 26513 115747 26571 115753
rect 27246 115744 27252 115796
rect 27304 115784 27310 115796
rect 27985 115787 28043 115793
rect 27985 115784 27997 115787
rect 27304 115756 27997 115784
rect 27304 115744 27310 115756
rect 27985 115753 27997 115756
rect 28031 115753 28043 115787
rect 27985 115747 28043 115753
rect 29454 115744 29460 115796
rect 29512 115784 29518 115796
rect 29641 115787 29699 115793
rect 29641 115784 29653 115787
rect 29512 115756 29653 115784
rect 29512 115744 29518 115756
rect 29641 115753 29653 115756
rect 29687 115753 29699 115787
rect 29641 115747 29699 115753
rect 29730 115744 29736 115796
rect 29788 115784 29794 115796
rect 30377 115787 30435 115793
rect 30377 115784 30389 115787
rect 29788 115756 30389 115784
rect 29788 115744 29794 115756
rect 30377 115753 30389 115756
rect 30423 115753 30435 115787
rect 30377 115747 30435 115753
rect 30929 115787 30987 115793
rect 30929 115753 30941 115787
rect 30975 115784 30987 115787
rect 31018 115784 31024 115796
rect 30975 115756 31024 115784
rect 30975 115753 30987 115756
rect 30929 115747 30987 115753
rect 31018 115744 31024 115756
rect 31076 115744 31082 115796
rect 31202 115744 31208 115796
rect 31260 115784 31266 115796
rect 31573 115787 31631 115793
rect 31573 115784 31585 115787
rect 31260 115756 31585 115784
rect 31260 115744 31266 115756
rect 31573 115753 31585 115756
rect 31619 115753 31631 115787
rect 31573 115747 31631 115753
rect 35802 115744 35808 115796
rect 35860 115784 35866 115796
rect 35989 115787 36047 115793
rect 35989 115784 36001 115787
rect 35860 115756 36001 115784
rect 35860 115744 35866 115756
rect 35989 115753 36001 115756
rect 36035 115753 36047 115787
rect 35989 115747 36047 115753
rect 36078 115744 36084 115796
rect 36136 115784 36142 115796
rect 36725 115787 36783 115793
rect 36725 115784 36737 115787
rect 36136 115756 36737 115784
rect 36136 115744 36142 115756
rect 36725 115753 36737 115756
rect 36771 115753 36783 115787
rect 36725 115747 36783 115753
rect 19107 115688 21312 115716
rect 24044 115688 24808 115716
rect 19107 115685 19119 115688
rect 19061 115679 19119 115685
rect 3712 115620 4292 115648
rect 4341 115651 4399 115657
rect 4341 115617 4353 115651
rect 4387 115648 4399 115651
rect 4614 115648 4620 115660
rect 4387 115620 4620 115648
rect 4387 115617 4399 115620
rect 4341 115611 4399 115617
rect 4614 115608 4620 115620
rect 4672 115608 4678 115660
rect 5074 115648 5080 115660
rect 5035 115620 5080 115648
rect 5074 115608 5080 115620
rect 5132 115608 5138 115660
rect 6914 115608 6920 115660
rect 6972 115648 6978 115660
rect 7009 115651 7067 115657
rect 7009 115648 7021 115651
rect 6972 115620 7021 115648
rect 6972 115608 6978 115620
rect 7009 115617 7021 115620
rect 7055 115617 7067 115651
rect 7009 115611 7067 115617
rect 8205 115651 8263 115657
rect 8205 115617 8217 115651
rect 8251 115617 8263 115651
rect 8205 115611 8263 115617
rect 1578 115540 1584 115592
rect 1636 115580 1642 115592
rect 5902 115580 5908 115592
rect 1636 115552 5908 115580
rect 1636 115540 1642 115552
rect 5902 115540 5908 115552
rect 5960 115540 5966 115592
rect 4522 115472 4528 115524
rect 4580 115512 4586 115524
rect 4706 115512 4712 115524
rect 4580 115484 4712 115512
rect 4580 115472 4586 115484
rect 4706 115472 4712 115484
rect 4764 115472 4770 115524
rect 8220 115512 8248 115611
rect 12158 115608 12164 115660
rect 12216 115648 12222 115660
rect 12253 115651 12311 115657
rect 12253 115648 12265 115651
rect 12216 115620 12265 115648
rect 12216 115608 12222 115620
rect 12253 115617 12265 115620
rect 12299 115617 12311 115651
rect 12894 115648 12900 115660
rect 12855 115620 12900 115648
rect 12253 115611 12311 115617
rect 12894 115608 12900 115620
rect 12952 115608 12958 115660
rect 17402 115608 17408 115660
rect 17460 115648 17466 115660
rect 17497 115651 17555 115657
rect 17497 115648 17509 115651
rect 17460 115620 17509 115648
rect 17460 115608 17466 115620
rect 17497 115617 17509 115620
rect 17543 115617 17555 115651
rect 17497 115611 17555 115617
rect 20533 115651 20591 115657
rect 20533 115617 20545 115651
rect 20579 115648 20591 115651
rect 21082 115648 21088 115660
rect 20579 115620 21088 115648
rect 20579 115617 20591 115620
rect 20533 115611 20591 115617
rect 21082 115608 21088 115620
rect 21140 115608 21146 115660
rect 21177 115651 21235 115657
rect 21177 115617 21189 115651
rect 21223 115648 21235 115651
rect 21634 115648 21640 115660
rect 21223 115620 21640 115648
rect 21223 115617 21235 115620
rect 21177 115611 21235 115617
rect 21634 115608 21640 115620
rect 21692 115608 21698 115660
rect 22741 115651 22799 115657
rect 22741 115617 22753 115651
rect 22787 115648 22799 115651
rect 22922 115648 22928 115660
rect 22787 115620 22928 115648
rect 22787 115617 22799 115620
rect 22741 115611 22799 115617
rect 22922 115608 22928 115620
rect 22980 115608 22986 115660
rect 23014 115608 23020 115660
rect 23072 115648 23078 115660
rect 23842 115648 23848 115660
rect 23072 115620 23848 115648
rect 23072 115608 23078 115620
rect 23842 115608 23848 115620
rect 23900 115608 23906 115660
rect 24044 115657 24072 115688
rect 25406 115676 25412 115728
rect 25464 115716 25470 115728
rect 30285 115719 30343 115725
rect 30285 115716 30297 115719
rect 25464 115688 30297 115716
rect 25464 115676 25470 115688
rect 30285 115685 30297 115688
rect 30331 115685 30343 115719
rect 31846 115716 31852 115728
rect 30285 115679 30343 115685
rect 31128 115688 31852 115716
rect 24029 115651 24087 115657
rect 24029 115617 24041 115651
rect 24075 115617 24087 115651
rect 24029 115611 24087 115617
rect 24302 115608 24308 115660
rect 24360 115648 24366 115660
rect 24673 115651 24731 115657
rect 24673 115648 24685 115651
rect 24360 115620 24685 115648
rect 24360 115608 24366 115620
rect 24673 115617 24685 115620
rect 24719 115617 24731 115651
rect 25498 115648 25504 115660
rect 25459 115620 25504 115648
rect 24673 115611 24731 115617
rect 25498 115608 25504 115620
rect 25556 115608 25562 115660
rect 26418 115648 26424 115660
rect 26379 115620 26424 115648
rect 26418 115608 26424 115620
rect 26476 115608 26482 115660
rect 27893 115651 27951 115657
rect 27893 115617 27905 115651
rect 27939 115617 27951 115651
rect 28718 115648 28724 115660
rect 28679 115620 28724 115648
rect 27893 115611 27951 115617
rect 15841 115583 15899 115589
rect 15841 115549 15853 115583
rect 15887 115580 15899 115583
rect 17770 115580 17776 115592
rect 15887 115552 17776 115580
rect 15887 115549 15899 115552
rect 15841 115543 15899 115549
rect 17770 115540 17776 115552
rect 17828 115540 17834 115592
rect 22002 115580 22008 115592
rect 18524 115552 22008 115580
rect 18524 115512 18552 115552
rect 22002 115540 22008 115552
rect 22060 115540 22066 115592
rect 22554 115540 22560 115592
rect 22612 115580 22618 115592
rect 27908 115580 27936 115611
rect 28718 115608 28724 115620
rect 28776 115608 28782 115660
rect 28810 115608 28816 115660
rect 28868 115648 28874 115660
rect 31128 115657 31156 115688
rect 31846 115676 31852 115688
rect 31904 115676 31910 115728
rect 33873 115719 33931 115725
rect 33873 115685 33885 115719
rect 33919 115716 33931 115719
rect 34514 115716 34520 115728
rect 33919 115688 34520 115716
rect 33919 115685 33931 115688
rect 33873 115679 33931 115685
rect 34514 115676 34520 115688
rect 34572 115676 34578 115728
rect 35342 115716 35348 115728
rect 35303 115688 35348 115716
rect 35342 115676 35348 115688
rect 35400 115676 35406 115728
rect 29549 115651 29607 115657
rect 29549 115648 29561 115651
rect 28868 115620 29561 115648
rect 28868 115608 28874 115620
rect 29549 115617 29561 115620
rect 29595 115617 29607 115651
rect 29549 115611 29607 115617
rect 31113 115651 31171 115657
rect 31113 115617 31125 115651
rect 31159 115617 31171 115651
rect 31113 115611 31171 115617
rect 31570 115608 31576 115660
rect 31628 115648 31634 115660
rect 31757 115651 31815 115657
rect 31757 115648 31769 115651
rect 31628 115620 31769 115648
rect 31628 115608 31634 115620
rect 31757 115617 31769 115620
rect 31803 115617 31815 115651
rect 31757 115611 31815 115617
rect 33689 115651 33747 115657
rect 33689 115617 33701 115651
rect 33735 115648 33747 115651
rect 33778 115648 33784 115660
rect 33735 115620 33784 115648
rect 33735 115617 33747 115620
rect 33689 115611 33747 115617
rect 33778 115608 33784 115620
rect 33836 115608 33842 115660
rect 34330 115608 34336 115660
rect 34388 115648 34394 115660
rect 34425 115651 34483 115657
rect 34425 115648 34437 115651
rect 34388 115620 34437 115648
rect 34388 115608 34394 115620
rect 34425 115617 34437 115620
rect 34471 115617 34483 115651
rect 34425 115611 34483 115617
rect 35161 115651 35219 115657
rect 35161 115617 35173 115651
rect 35207 115617 35219 115651
rect 35161 115611 35219 115617
rect 35897 115651 35955 115657
rect 35897 115617 35909 115651
rect 35943 115648 35955 115651
rect 36262 115648 36268 115660
rect 35943 115620 36268 115648
rect 35943 115617 35955 115620
rect 35897 115611 35955 115617
rect 22612 115552 27936 115580
rect 22612 115540 22618 115552
rect 34514 115540 34520 115592
rect 34572 115580 34578 115592
rect 34882 115580 34888 115592
rect 34572 115552 34888 115580
rect 34572 115540 34578 115552
rect 34882 115540 34888 115552
rect 34940 115540 34946 115592
rect 35176 115580 35204 115611
rect 36262 115608 36268 115620
rect 36320 115608 36326 115660
rect 36630 115648 36636 115660
rect 36591 115620 36636 115648
rect 36630 115608 36636 115620
rect 36688 115608 36694 115660
rect 35342 115580 35348 115592
rect 35176 115552 35348 115580
rect 35342 115540 35348 115552
rect 35400 115540 35406 115592
rect 8220 115484 18552 115512
rect 19889 115515 19947 115521
rect 19889 115481 19901 115515
rect 19935 115512 19947 115515
rect 19935 115484 21312 115512
rect 19935 115481 19947 115484
rect 19889 115475 19947 115481
rect 1946 115444 1952 115456
rect 1907 115416 1952 115444
rect 1946 115404 1952 115416
rect 2004 115404 2010 115456
rect 10042 115404 10048 115456
rect 10100 115444 10106 115456
rect 10870 115444 10876 115456
rect 10100 115416 10876 115444
rect 10100 115404 10106 115416
rect 10870 115404 10876 115416
rect 10928 115404 10934 115456
rect 21284 115444 21312 115484
rect 21634 115472 21640 115524
rect 21692 115512 21698 115524
rect 23198 115512 23204 115524
rect 21692 115484 23204 115512
rect 21692 115472 21698 115484
rect 23198 115472 23204 115484
rect 23256 115472 23262 115524
rect 24118 115512 24124 115524
rect 23308 115484 24124 115512
rect 23308 115444 23336 115484
rect 24118 115472 24124 115484
rect 24176 115472 24182 115524
rect 24670 115472 24676 115524
rect 24728 115512 24734 115524
rect 24728 115484 25820 115512
rect 24728 115472 24734 115484
rect 21284 115416 23336 115444
rect 23385 115447 23443 115453
rect 23385 115413 23397 115447
rect 23431 115444 23443 115447
rect 25130 115444 25136 115456
rect 23431 115416 25136 115444
rect 23431 115413 23443 115416
rect 23385 115407 23443 115413
rect 25130 115404 25136 115416
rect 25188 115404 25194 115456
rect 25792 115444 25820 115484
rect 25866 115472 25872 115524
rect 25924 115512 25930 115524
rect 28537 115515 28595 115521
rect 28537 115512 28549 115515
rect 25924 115484 28549 115512
rect 25924 115472 25930 115484
rect 28537 115481 28549 115484
rect 28583 115481 28595 115515
rect 28537 115475 28595 115481
rect 34609 115515 34667 115521
rect 34609 115481 34621 115515
rect 34655 115512 34667 115515
rect 39482 115512 39488 115524
rect 34655 115484 39488 115512
rect 34655 115481 34667 115484
rect 34609 115475 34667 115481
rect 39482 115472 39488 115484
rect 39540 115472 39546 115524
rect 29178 115444 29184 115456
rect 25792 115416 29184 115444
rect 29178 115404 29184 115416
rect 29236 115404 29242 115456
rect 29730 115404 29736 115456
rect 29788 115444 29794 115456
rect 33410 115444 33416 115456
rect 29788 115416 33416 115444
rect 29788 115404 29794 115416
rect 33410 115404 33416 115416
rect 33468 115404 33474 115456
rect 1104 115354 38824 115376
rect 1104 115302 4246 115354
rect 4298 115302 4310 115354
rect 4362 115302 4374 115354
rect 4426 115302 4438 115354
rect 4490 115302 34966 115354
rect 35018 115302 35030 115354
rect 35082 115302 35094 115354
rect 35146 115302 35158 115354
rect 35210 115302 38824 115354
rect 1104 115280 38824 115302
rect 1394 115200 1400 115252
rect 1452 115240 1458 115252
rect 1949 115243 2007 115249
rect 1949 115240 1961 115243
rect 1452 115212 1961 115240
rect 1452 115200 1458 115212
rect 1949 115209 1961 115212
rect 1995 115209 2007 115243
rect 1949 115203 2007 115209
rect 4062 115200 4068 115252
rect 4120 115240 4126 115252
rect 4433 115243 4491 115249
rect 4433 115240 4445 115243
rect 4120 115212 4445 115240
rect 4120 115200 4126 115212
rect 4433 115209 4445 115212
rect 4479 115209 4491 115243
rect 4433 115203 4491 115209
rect 5077 115243 5135 115249
rect 5077 115209 5089 115243
rect 5123 115240 5135 115243
rect 5534 115240 5540 115252
rect 5123 115212 5540 115240
rect 5123 115209 5135 115212
rect 5077 115203 5135 115209
rect 5534 115200 5540 115212
rect 5592 115200 5598 115252
rect 6270 115200 6276 115252
rect 6328 115240 6334 115252
rect 7101 115243 7159 115249
rect 7101 115240 7113 115243
rect 6328 115212 7113 115240
rect 6328 115200 6334 115212
rect 7101 115209 7113 115212
rect 7147 115209 7159 115243
rect 7101 115203 7159 115209
rect 7926 115200 7932 115252
rect 7984 115240 7990 115252
rect 8113 115243 8171 115249
rect 8113 115240 8125 115243
rect 7984 115212 8125 115240
rect 7984 115200 7990 115212
rect 8113 115209 8125 115212
rect 8159 115209 8171 115243
rect 8113 115203 8171 115209
rect 9677 115243 9735 115249
rect 9677 115209 9689 115243
rect 9723 115240 9735 115243
rect 9858 115240 9864 115252
rect 9723 115212 9864 115240
rect 9723 115209 9735 115212
rect 9677 115203 9735 115209
rect 9858 115200 9864 115212
rect 9916 115200 9922 115252
rect 10321 115243 10379 115249
rect 10321 115209 10333 115243
rect 10367 115240 10379 115243
rect 10594 115240 10600 115252
rect 10367 115212 10600 115240
rect 10367 115209 10379 115212
rect 10321 115203 10379 115209
rect 10594 115200 10600 115212
rect 10652 115200 10658 115252
rect 10962 115240 10968 115252
rect 10923 115212 10968 115240
rect 10962 115200 10968 115212
rect 11020 115200 11026 115252
rect 11238 115200 11244 115252
rect 11296 115240 11302 115252
rect 11609 115243 11667 115249
rect 11609 115240 11621 115243
rect 11296 115212 11621 115240
rect 11296 115200 11302 115212
rect 11609 115209 11621 115212
rect 11655 115209 11667 115243
rect 12986 115240 12992 115252
rect 12947 115212 12992 115240
rect 11609 115203 11667 115209
rect 12986 115200 12992 115212
rect 13044 115200 13050 115252
rect 13633 115243 13691 115249
rect 13633 115209 13645 115243
rect 13679 115240 13691 115243
rect 14366 115240 14372 115252
rect 13679 115212 14372 115240
rect 13679 115209 13691 115212
rect 13633 115203 13691 115209
rect 14366 115200 14372 115212
rect 14424 115200 14430 115252
rect 14921 115243 14979 115249
rect 14921 115209 14933 115243
rect 14967 115240 14979 115243
rect 15102 115240 15108 115252
rect 14967 115212 15108 115240
rect 14967 115209 14979 115212
rect 14921 115203 14979 115209
rect 15102 115200 15108 115212
rect 15160 115200 15166 115252
rect 15562 115240 15568 115252
rect 15523 115212 15568 115240
rect 15562 115200 15568 115212
rect 15620 115200 15626 115252
rect 15654 115200 15660 115252
rect 15712 115240 15718 115252
rect 16209 115243 16267 115249
rect 16209 115240 16221 115243
rect 15712 115212 16221 115240
rect 15712 115200 15718 115212
rect 16209 115209 16221 115212
rect 16255 115209 16267 115243
rect 16209 115203 16267 115209
rect 16390 115200 16396 115252
rect 16448 115240 16454 115252
rect 16853 115243 16911 115249
rect 16853 115240 16865 115243
rect 16448 115212 16865 115240
rect 16448 115200 16454 115212
rect 16853 115209 16865 115212
rect 16899 115209 16911 115243
rect 16853 115203 16911 115209
rect 17497 115243 17555 115249
rect 17497 115209 17509 115243
rect 17543 115240 17555 115243
rect 18138 115240 18144 115252
rect 17543 115212 18144 115240
rect 17543 115209 17555 115212
rect 17497 115203 17555 115209
rect 18138 115200 18144 115212
rect 18196 115200 18202 115252
rect 18785 115243 18843 115249
rect 18785 115209 18797 115243
rect 18831 115240 18843 115243
rect 19334 115240 19340 115252
rect 18831 115212 19340 115240
rect 18831 115209 18843 115212
rect 18785 115203 18843 115209
rect 19334 115200 19340 115212
rect 19392 115200 19398 115252
rect 20165 115243 20223 115249
rect 20165 115209 20177 115243
rect 20211 115240 20223 115243
rect 20346 115240 20352 115252
rect 20211 115212 20352 115240
rect 20211 115209 20223 115212
rect 20165 115203 20223 115209
rect 20346 115200 20352 115212
rect 20404 115200 20410 115252
rect 20625 115243 20683 115249
rect 20625 115209 20637 115243
rect 20671 115240 20683 115243
rect 20714 115240 20720 115252
rect 20671 115212 20720 115240
rect 20671 115209 20683 115212
rect 20625 115203 20683 115209
rect 20714 115200 20720 115212
rect 20772 115200 20778 115252
rect 21634 115240 21640 115252
rect 21595 115212 21640 115240
rect 21634 115200 21640 115212
rect 21692 115200 21698 115252
rect 22094 115240 22100 115252
rect 22055 115212 22100 115240
rect 22094 115200 22100 115212
rect 22152 115200 22158 115252
rect 25409 115243 25467 115249
rect 25409 115209 25421 115243
rect 25455 115240 25467 115243
rect 25774 115240 25780 115252
rect 25455 115212 25780 115240
rect 25455 115209 25467 115212
rect 25409 115203 25467 115209
rect 25774 115200 25780 115212
rect 25832 115200 25838 115252
rect 26053 115243 26111 115249
rect 26053 115209 26065 115243
rect 26099 115240 26111 115243
rect 26510 115240 26516 115252
rect 26099 115212 26516 115240
rect 26099 115209 26111 115212
rect 26053 115203 26111 115209
rect 26510 115200 26516 115212
rect 26568 115200 26574 115252
rect 27614 115200 27620 115252
rect 27672 115240 27678 115252
rect 27801 115243 27859 115249
rect 27801 115240 27813 115243
rect 27672 115212 27813 115240
rect 27672 115200 27678 115212
rect 27801 115209 27813 115212
rect 27847 115209 27859 115243
rect 27801 115203 27859 115209
rect 28902 115200 28908 115252
rect 28960 115240 28966 115252
rect 31110 115240 31116 115252
rect 28960 115212 30052 115240
rect 31071 115212 31116 115240
rect 28960 115200 28966 115212
rect 2777 115175 2835 115181
rect 2777 115141 2789 115175
rect 2823 115172 2835 115175
rect 2866 115172 2872 115184
rect 2823 115144 2872 115172
rect 2823 115141 2835 115144
rect 2777 115135 2835 115141
rect 2866 115132 2872 115144
rect 2924 115132 2930 115184
rect 5350 115132 5356 115184
rect 5408 115172 5414 115184
rect 5813 115175 5871 115181
rect 5813 115172 5825 115175
rect 5408 115144 5825 115172
rect 5408 115132 5414 115144
rect 5813 115141 5825 115144
rect 5859 115141 5871 115175
rect 18690 115172 18696 115184
rect 5813 115135 5871 115141
rect 9968 115144 18696 115172
rect 5442 115064 5448 115116
rect 5500 115104 5506 115116
rect 6457 115107 6515 115113
rect 6457 115104 6469 115107
rect 5500 115076 6469 115104
rect 5500 115064 5506 115076
rect 6457 115073 6469 115076
rect 6503 115073 6515 115107
rect 6457 115067 6515 115073
rect 9858 115064 9864 115116
rect 9916 115104 9922 115116
rect 9968 115104 9996 115144
rect 18690 115132 18696 115144
rect 18748 115132 18754 115184
rect 22741 115175 22799 115181
rect 22741 115141 22753 115175
rect 22787 115172 22799 115175
rect 22787 115144 24440 115172
rect 22787 115141 22799 115144
rect 22741 115135 22799 115141
rect 9916 115076 9996 115104
rect 9916 115064 9922 115076
rect 10686 115064 10692 115116
rect 10744 115104 10750 115116
rect 18141 115107 18199 115113
rect 10744 115076 12296 115104
rect 10744 115064 10750 115076
rect 2593 115039 2651 115045
rect 2593 115005 2605 115039
rect 2639 115036 2651 115039
rect 2682 115036 2688 115048
rect 2639 115008 2688 115036
rect 2639 115005 2651 115008
rect 2593 114999 2651 115005
rect 2682 114996 2688 115008
rect 2740 114996 2746 115048
rect 6270 114996 6276 115048
rect 6328 115036 6334 115048
rect 10962 115036 10968 115048
rect 6328 115008 10968 115036
rect 6328 114996 6334 115008
rect 10962 114996 10968 115008
rect 11020 114996 11026 115048
rect 12268 115045 12296 115076
rect 18141 115073 18153 115107
rect 18187 115104 18199 115107
rect 18874 115104 18880 115116
rect 18187 115076 18880 115104
rect 18187 115073 18199 115076
rect 18141 115067 18199 115073
rect 18874 115064 18880 115076
rect 18932 115064 18938 115116
rect 19334 115064 19340 115116
rect 19392 115104 19398 115116
rect 24412 115104 24440 115144
rect 26418 115132 26424 115184
rect 26476 115172 26482 115184
rect 28997 115175 29055 115181
rect 28997 115172 29009 115175
rect 26476 115144 29009 115172
rect 26476 115132 26482 115144
rect 28997 115141 29009 115144
rect 29043 115141 29055 115175
rect 28997 115135 29055 115141
rect 27522 115104 27528 115116
rect 19392 115076 23612 115104
rect 24412 115076 27528 115104
rect 19392 115064 19398 115076
rect 12253 115039 12311 115045
rect 12253 115005 12265 115039
rect 12299 115005 12311 115039
rect 12253 114999 12311 115005
rect 15286 114996 15292 115048
rect 15344 115036 15350 115048
rect 23584 115045 23612 115076
rect 27522 115064 27528 115076
rect 27580 115064 27586 115116
rect 28350 115064 28356 115116
rect 28408 115104 28414 115116
rect 28408 115076 29224 115104
rect 28408 115064 28414 115076
rect 20809 115039 20867 115045
rect 20809 115036 20821 115039
rect 15344 115008 20821 115036
rect 15344 114996 15350 115008
rect 20809 115005 20821 115008
rect 20855 115005 20867 115039
rect 22281 115039 22339 115045
rect 22281 115036 22293 115039
rect 20809 114999 20867 115005
rect 22066 115008 22293 115036
rect 1854 114968 1860 114980
rect 1815 114940 1860 114968
rect 1854 114928 1860 114940
rect 1912 114928 1918 114980
rect 5626 114968 5632 114980
rect 5587 114940 5632 114968
rect 5626 114928 5632 114940
rect 5684 114928 5690 114980
rect 8018 114968 8024 114980
rect 7979 114940 8024 114968
rect 8018 114928 8024 114940
rect 8076 114928 8082 114980
rect 9398 114928 9404 114980
rect 9456 114968 9462 114980
rect 10502 114968 10508 114980
rect 9456 114940 10508 114968
rect 9456 114928 9462 114940
rect 10502 114928 10508 114940
rect 10560 114928 10566 114980
rect 11882 114928 11888 114980
rect 11940 114968 11946 114980
rect 12894 114968 12900 114980
rect 11940 114940 12900 114968
rect 11940 114928 11946 114940
rect 12894 114928 12900 114940
rect 12952 114928 12958 114980
rect 17310 114928 17316 114980
rect 17368 114968 17374 114980
rect 22066 114968 22094 115008
rect 22281 115005 22293 115008
rect 22327 115005 22339 115039
rect 22281 114999 22339 115005
rect 22925 115039 22983 115045
rect 22925 115005 22937 115039
rect 22971 115005 22983 115039
rect 22925 114999 22983 115005
rect 23569 115039 23627 115045
rect 23569 115005 23581 115039
rect 23615 115005 23627 115039
rect 23569 114999 23627 115005
rect 24305 115039 24363 115045
rect 24305 115005 24317 115039
rect 24351 115005 24363 115039
rect 26694 115036 26700 115048
rect 26655 115008 26700 115036
rect 24305 114999 24363 115005
rect 22940 114968 22968 114999
rect 17368 114940 22094 114968
rect 22480 114940 22968 114968
rect 17368 114928 17374 114940
rect 8386 114860 8392 114912
rect 8444 114900 8450 114912
rect 12069 114903 12127 114909
rect 12069 114900 12081 114903
rect 8444 114872 12081 114900
rect 8444 114860 8450 114872
rect 12069 114869 12081 114872
rect 12115 114869 12127 114903
rect 12069 114863 12127 114869
rect 12526 114860 12532 114912
rect 12584 114900 12590 114912
rect 13538 114900 13544 114912
rect 12584 114872 13544 114900
rect 12584 114860 12590 114872
rect 13538 114860 13544 114872
rect 13596 114860 13602 114912
rect 18874 114860 18880 114912
rect 18932 114900 18938 114912
rect 20898 114900 20904 114912
rect 18932 114872 20904 114900
rect 18932 114860 18938 114872
rect 20898 114860 20904 114872
rect 20956 114860 20962 114912
rect 20990 114860 20996 114912
rect 21048 114900 21054 114912
rect 22480 114900 22508 114940
rect 23106 114928 23112 114980
rect 23164 114968 23170 114980
rect 24320 114968 24348 114999
rect 26694 114996 26700 115008
rect 26752 114996 26758 115048
rect 27798 114996 27804 115048
rect 27856 115036 27862 115048
rect 29196 115045 29224 115076
rect 28537 115039 28595 115045
rect 28537 115036 28549 115039
rect 27856 115008 28549 115036
rect 27856 114996 27862 115008
rect 28537 115005 28549 115008
rect 28583 115005 28595 115039
rect 28537 114999 28595 115005
rect 29181 115039 29239 115045
rect 29181 115005 29193 115039
rect 29227 115005 29239 115039
rect 30024 115036 30052 115212
rect 31110 115200 31116 115212
rect 31168 115200 31174 115252
rect 31662 115200 31668 115252
rect 31720 115240 31726 115252
rect 31757 115243 31815 115249
rect 31757 115240 31769 115243
rect 31720 115212 31769 115240
rect 31720 115200 31726 115212
rect 31757 115209 31769 115212
rect 31803 115209 31815 115243
rect 32398 115240 32404 115252
rect 32359 115212 32404 115240
rect 31757 115203 31815 115209
rect 32398 115200 32404 115212
rect 32456 115200 32462 115252
rect 34701 115243 34759 115249
rect 34701 115209 34713 115243
rect 34747 115240 34759 115243
rect 36906 115240 36912 115252
rect 34747 115212 36912 115240
rect 34747 115209 34759 115212
rect 34701 115203 34759 115209
rect 36906 115200 36912 115212
rect 36964 115200 36970 115252
rect 37090 115240 37096 115252
rect 37051 115212 37096 115240
rect 37090 115200 37096 115212
rect 37148 115200 37154 115252
rect 32582 115132 32588 115184
rect 32640 115132 32646 115184
rect 34057 115175 34115 115181
rect 34057 115141 34069 115175
rect 34103 115172 34115 115175
rect 34514 115172 34520 115184
rect 34103 115144 34520 115172
rect 34103 115141 34115 115144
rect 34057 115135 34115 115141
rect 34514 115132 34520 115144
rect 34572 115132 34578 115184
rect 36449 115175 36507 115181
rect 36449 115141 36461 115175
rect 36495 115172 36507 115175
rect 38010 115172 38016 115184
rect 36495 115144 38016 115172
rect 36495 115141 36507 115144
rect 36449 115135 36507 115141
rect 38010 115132 38016 115144
rect 38068 115132 38074 115184
rect 32600 115104 32628 115132
rect 31312 115076 32628 115104
rect 33321 115107 33379 115113
rect 31312 115045 31340 115076
rect 33321 115073 33333 115107
rect 33367 115104 33379 115107
rect 37550 115104 37556 115116
rect 33367 115076 37556 115104
rect 33367 115073 33379 115076
rect 33321 115067 33379 115073
rect 37550 115064 37556 115076
rect 37608 115064 37614 115116
rect 30653 115039 30711 115045
rect 30653 115036 30665 115039
rect 30024 115008 30665 115036
rect 29181 114999 29239 115005
rect 30653 115005 30665 115008
rect 30699 115005 30711 115039
rect 30653 114999 30711 115005
rect 31297 115039 31355 115045
rect 31297 115005 31309 115039
rect 31343 115005 31355 115039
rect 31297 114999 31355 115005
rect 31941 115039 31999 115045
rect 31941 115005 31953 115039
rect 31987 115036 31999 115039
rect 32030 115036 32036 115048
rect 31987 115008 32036 115036
rect 31987 115005 31999 115008
rect 31941 114999 31999 115005
rect 32030 114996 32036 115008
rect 32088 114996 32094 115048
rect 32585 115039 32643 115045
rect 32585 115005 32597 115039
rect 32631 115036 32643 115039
rect 33962 115036 33968 115048
rect 32631 115008 33968 115036
rect 32631 115005 32643 115008
rect 32585 114999 32643 115005
rect 33962 114996 33968 115008
rect 34020 114996 34026 115048
rect 35066 114996 35072 115048
rect 35124 115036 35130 115048
rect 36722 115036 36728 115048
rect 35124 115008 36728 115036
rect 35124 114996 35130 115008
rect 36722 114996 36728 115008
rect 36780 114996 36786 115048
rect 37642 115036 37648 115048
rect 37603 115008 37648 115036
rect 37642 114996 37648 115008
rect 37700 114996 37706 115048
rect 27706 114968 27712 114980
rect 23164 114940 24164 114968
rect 24320 114940 27568 114968
rect 27667 114940 27712 114968
rect 23164 114928 23170 114940
rect 21048 114872 22508 114900
rect 21048 114860 21054 114872
rect 23290 114860 23296 114912
rect 23348 114900 23354 114912
rect 24136 114909 24164 114940
rect 23385 114903 23443 114909
rect 23385 114900 23397 114903
rect 23348 114872 23397 114900
rect 23348 114860 23354 114872
rect 23385 114869 23397 114872
rect 23431 114869 23443 114903
rect 23385 114863 23443 114869
rect 24121 114903 24179 114909
rect 24121 114869 24133 114903
rect 24167 114869 24179 114903
rect 24121 114863 24179 114869
rect 26050 114860 26056 114912
rect 26108 114900 26114 114912
rect 26513 114903 26571 114909
rect 26513 114900 26525 114903
rect 26108 114872 26525 114900
rect 26108 114860 26114 114872
rect 26513 114869 26525 114872
rect 26559 114869 26571 114903
rect 27540 114900 27568 114940
rect 27706 114928 27712 114940
rect 27764 114928 27770 114980
rect 29086 114968 29092 114980
rect 27816 114940 29092 114968
rect 27816 114900 27844 114940
rect 29086 114928 29092 114940
rect 29144 114928 29150 114980
rect 32398 114928 32404 114980
rect 32456 114968 32462 114980
rect 33137 114971 33195 114977
rect 33137 114968 33149 114971
rect 32456 114940 33149 114968
rect 32456 114928 32462 114940
rect 33137 114937 33149 114940
rect 33183 114937 33195 114971
rect 33137 114931 33195 114937
rect 33410 114928 33416 114980
rect 33468 114968 33474 114980
rect 33873 114971 33931 114977
rect 33873 114968 33885 114971
rect 33468 114940 33885 114968
rect 33468 114928 33474 114940
rect 33873 114937 33885 114940
rect 33919 114937 33931 114971
rect 33873 114931 33931 114937
rect 34514 114928 34520 114980
rect 34572 114968 34578 114980
rect 34609 114971 34667 114977
rect 34609 114968 34621 114971
rect 34572 114940 34621 114968
rect 34572 114928 34578 114940
rect 34609 114937 34621 114940
rect 34655 114937 34667 114971
rect 34609 114931 34667 114937
rect 35986 114928 35992 114980
rect 36044 114968 36050 114980
rect 36265 114971 36323 114977
rect 36265 114968 36277 114971
rect 36044 114940 36277 114968
rect 36044 114928 36050 114940
rect 36265 114937 36277 114940
rect 36311 114937 36323 114971
rect 36265 114931 36323 114937
rect 36906 114928 36912 114980
rect 36964 114968 36970 114980
rect 37001 114971 37059 114977
rect 37001 114968 37013 114971
rect 36964 114940 37013 114968
rect 36964 114928 36970 114940
rect 37001 114937 37013 114940
rect 37047 114937 37059 114971
rect 37001 114931 37059 114937
rect 37921 114971 37979 114977
rect 37921 114937 37933 114971
rect 37967 114968 37979 114971
rect 38286 114968 38292 114980
rect 37967 114940 38292 114968
rect 37967 114937 37979 114940
rect 37921 114931 37979 114937
rect 38286 114928 38292 114940
rect 38344 114928 38350 114980
rect 27540 114872 27844 114900
rect 26513 114863 26571 114869
rect 27890 114860 27896 114912
rect 27948 114900 27954 114912
rect 28353 114903 28411 114909
rect 28353 114900 28365 114903
rect 27948 114872 28365 114900
rect 27948 114860 27954 114872
rect 28353 114869 28365 114872
rect 28399 114869 28411 114903
rect 30466 114900 30472 114912
rect 30427 114872 30472 114900
rect 28353 114863 28411 114869
rect 30466 114860 30472 114872
rect 30524 114860 30530 114912
rect 1104 114810 38824 114832
rect 1104 114758 19606 114810
rect 19658 114758 19670 114810
rect 19722 114758 19734 114810
rect 19786 114758 19798 114810
rect 19850 114758 38824 114810
rect 1104 114736 38824 114758
rect 6638 114656 6644 114708
rect 6696 114696 6702 114708
rect 10321 114699 10379 114705
rect 10321 114696 10333 114699
rect 6696 114668 10333 114696
rect 6696 114656 6702 114668
rect 10321 114665 10333 114668
rect 10367 114665 10379 114699
rect 10321 114659 10379 114665
rect 10410 114656 10416 114708
rect 10468 114696 10474 114708
rect 12713 114699 12771 114705
rect 12713 114696 12725 114699
rect 10468 114668 12725 114696
rect 10468 114656 10474 114668
rect 12713 114665 12725 114668
rect 12759 114665 12771 114699
rect 12713 114659 12771 114665
rect 14001 114699 14059 114705
rect 14001 114665 14013 114699
rect 14047 114665 14059 114699
rect 14001 114659 14059 114665
rect 1857 114631 1915 114637
rect 1857 114597 1869 114631
rect 1903 114628 1915 114631
rect 3510 114628 3516 114640
rect 1903 114600 3516 114628
rect 1903 114597 1915 114600
rect 1857 114591 1915 114597
rect 3510 114588 3516 114600
rect 3568 114588 3574 114640
rect 14016 114628 14044 114659
rect 14458 114656 14464 114708
rect 14516 114696 14522 114708
rect 15933 114699 15991 114705
rect 14516 114668 15516 114696
rect 14516 114656 14522 114668
rect 9232 114600 14044 114628
rect 14108 114600 14872 114628
rect 2406 114520 2412 114572
rect 2464 114560 2470 114572
rect 2593 114563 2651 114569
rect 2593 114560 2605 114563
rect 2464 114532 2605 114560
rect 2464 114520 2470 114532
rect 2593 114529 2605 114532
rect 2639 114529 2651 114563
rect 2593 114523 2651 114529
rect 3329 114563 3387 114569
rect 3329 114529 3341 114563
rect 3375 114560 3387 114563
rect 3694 114560 3700 114572
rect 3375 114532 3700 114560
rect 3375 114529 3387 114532
rect 3329 114523 3387 114529
rect 3694 114520 3700 114532
rect 3752 114520 3758 114572
rect 4982 114520 4988 114572
rect 5040 114560 5046 114572
rect 5534 114560 5540 114572
rect 5040 114532 5540 114560
rect 5040 114520 5046 114532
rect 5534 114520 5540 114532
rect 5592 114520 5598 114572
rect 6546 114520 6552 114572
rect 6604 114560 6610 114572
rect 6604 114532 8156 114560
rect 6604 114520 6610 114532
rect 2038 114492 2044 114504
rect 1999 114464 2044 114492
rect 2038 114452 2044 114464
rect 2096 114452 2102 114504
rect 2777 114495 2835 114501
rect 2777 114461 2789 114495
rect 2823 114492 2835 114495
rect 3234 114492 3240 114504
rect 2823 114464 3240 114492
rect 2823 114461 2835 114464
rect 2777 114455 2835 114461
rect 3234 114452 3240 114464
rect 3292 114452 3298 114504
rect 4157 114495 4215 114501
rect 4157 114461 4169 114495
rect 4203 114492 4215 114495
rect 4798 114492 4804 114504
rect 4203 114464 4804 114492
rect 4203 114461 4215 114464
rect 4157 114455 4215 114461
rect 4798 114452 4804 114464
rect 4856 114452 4862 114504
rect 5077 114495 5135 114501
rect 5077 114461 5089 114495
rect 5123 114492 5135 114495
rect 5718 114492 5724 114504
rect 5123 114464 5724 114492
rect 5123 114461 5135 114464
rect 5077 114455 5135 114461
rect 5718 114452 5724 114464
rect 5776 114452 5782 114504
rect 7006 114492 7012 114504
rect 6967 114464 7012 114492
rect 7006 114452 7012 114464
rect 7064 114452 7070 114504
rect 7558 114452 7564 114504
rect 7616 114492 7622 114504
rect 7653 114495 7711 114501
rect 7653 114492 7665 114495
rect 7616 114464 7665 114492
rect 7616 114452 7622 114464
rect 7653 114461 7665 114464
rect 7699 114461 7711 114495
rect 7653 114455 7711 114461
rect 3326 114316 3332 114368
rect 3384 114356 3390 114368
rect 3421 114359 3479 114365
rect 3421 114356 3433 114359
rect 3384 114328 3433 114356
rect 3384 114316 3390 114328
rect 3421 114325 3433 114328
rect 3467 114325 3479 114359
rect 3421 114319 3479 114325
rect 5074 114316 5080 114368
rect 5132 114356 5138 114368
rect 5721 114359 5779 114365
rect 5721 114356 5733 114359
rect 5132 114328 5733 114356
rect 5132 114316 5138 114328
rect 5721 114325 5733 114328
rect 5767 114325 5779 114359
rect 8128 114356 8156 114532
rect 8202 114520 8208 114572
rect 8260 114560 8266 114572
rect 9232 114569 9260 114600
rect 9217 114563 9275 114569
rect 8260 114532 9168 114560
rect 8260 114520 8266 114532
rect 8570 114492 8576 114504
rect 8531 114464 8576 114492
rect 8570 114452 8576 114464
rect 8628 114452 8634 114504
rect 9140 114492 9168 114532
rect 9217 114529 9229 114563
rect 9263 114529 9275 114563
rect 9677 114563 9735 114569
rect 9677 114560 9689 114563
rect 9217 114523 9275 114529
rect 9324 114532 9689 114560
rect 9324 114492 9352 114532
rect 9677 114529 9689 114532
rect 9723 114529 9735 114563
rect 10502 114560 10508 114572
rect 10463 114532 10508 114560
rect 9677 114523 9735 114529
rect 10502 114520 10508 114532
rect 10560 114520 10566 114572
rect 10870 114520 10876 114572
rect 10928 114560 10934 114572
rect 11149 114563 11207 114569
rect 11149 114560 11161 114563
rect 10928 114532 11161 114560
rect 10928 114520 10934 114532
rect 11149 114529 11161 114532
rect 11195 114529 11207 114563
rect 11149 114523 11207 114529
rect 11422 114520 11428 114572
rect 11480 114560 11486 114572
rect 12253 114563 12311 114569
rect 12253 114560 12265 114563
rect 11480 114532 12265 114560
rect 11480 114520 11486 114532
rect 12253 114529 12265 114532
rect 12299 114529 12311 114563
rect 12894 114560 12900 114572
rect 12855 114532 12900 114560
rect 12253 114523 12311 114529
rect 12894 114520 12900 114532
rect 12952 114520 12958 114572
rect 13262 114520 13268 114572
rect 13320 114560 13326 114572
rect 13320 114532 13492 114560
rect 13320 114520 13326 114532
rect 9140 114464 9352 114492
rect 13464 114492 13492 114532
rect 13538 114520 13544 114572
rect 13596 114560 13602 114572
rect 13596 114532 13641 114560
rect 13596 114520 13602 114532
rect 13906 114520 13912 114572
rect 13964 114560 13970 114572
rect 14108 114560 14136 114600
rect 14844 114569 14872 114600
rect 13964 114532 14136 114560
rect 14185 114563 14243 114569
rect 13964 114520 13970 114532
rect 14185 114529 14197 114563
rect 14231 114529 14243 114563
rect 14185 114523 14243 114529
rect 14829 114563 14887 114569
rect 14829 114529 14841 114563
rect 14875 114529 14887 114563
rect 14829 114523 14887 114529
rect 14200 114492 14228 114523
rect 14918 114520 14924 114572
rect 14976 114560 14982 114572
rect 15488 114569 15516 114668
rect 15933 114665 15945 114699
rect 15979 114665 15991 114699
rect 17310 114696 17316 114708
rect 17271 114668 17316 114696
rect 15933 114659 15991 114665
rect 15948 114628 15976 114659
rect 17310 114656 17316 114668
rect 17368 114656 17374 114708
rect 18233 114699 18291 114705
rect 18233 114665 18245 114699
rect 18279 114696 18291 114699
rect 20714 114696 20720 114708
rect 18279 114668 20720 114696
rect 18279 114665 18291 114668
rect 18233 114659 18291 114665
rect 20714 114656 20720 114668
rect 20772 114656 20778 114708
rect 20809 114699 20867 114705
rect 20809 114665 20821 114699
rect 20855 114696 20867 114699
rect 21358 114696 21364 114708
rect 20855 114668 21364 114696
rect 20855 114665 20867 114668
rect 20809 114659 20867 114665
rect 21358 114656 21364 114668
rect 21416 114656 21422 114708
rect 21453 114699 21511 114705
rect 21453 114665 21465 114699
rect 21499 114696 21511 114699
rect 21726 114696 21732 114708
rect 21499 114668 21732 114696
rect 21499 114665 21511 114668
rect 21453 114659 21511 114665
rect 21726 114656 21732 114668
rect 21784 114656 21790 114708
rect 22554 114696 22560 114708
rect 22515 114668 22560 114696
rect 22554 114656 22560 114668
rect 22612 114656 22618 114708
rect 23658 114656 23664 114708
rect 23716 114696 23722 114708
rect 24029 114699 24087 114705
rect 24029 114696 24041 114699
rect 23716 114668 24041 114696
rect 23716 114656 23722 114668
rect 24029 114665 24041 114668
rect 24075 114665 24087 114699
rect 27890 114696 27896 114708
rect 24029 114659 24087 114665
rect 24228 114668 27896 114696
rect 15948 114600 18920 114628
rect 15473 114563 15531 114569
rect 14976 114532 15424 114560
rect 14976 114520 14982 114532
rect 13464 114464 14228 114492
rect 15396 114492 15424 114532
rect 15473 114529 15485 114563
rect 15519 114529 15531 114563
rect 16117 114563 16175 114569
rect 16117 114560 16129 114563
rect 15473 114523 15531 114529
rect 15580 114532 16129 114560
rect 15580 114492 15608 114532
rect 16117 114529 16129 114532
rect 16163 114529 16175 114563
rect 16117 114523 16175 114529
rect 17034 114520 17040 114572
rect 17092 114560 17098 114572
rect 17497 114563 17555 114569
rect 17497 114560 17509 114563
rect 17092 114532 17509 114560
rect 17092 114520 17098 114532
rect 17497 114529 17509 114532
rect 17543 114529 17555 114563
rect 18046 114560 18052 114572
rect 18007 114532 18052 114560
rect 17497 114523 17555 114529
rect 18046 114520 18052 114532
rect 18104 114520 18110 114572
rect 18690 114560 18696 114572
rect 18651 114532 18696 114560
rect 18690 114520 18696 114532
rect 18748 114520 18754 114572
rect 15396 114464 15608 114492
rect 18892 114492 18920 114600
rect 19426 114588 19432 114640
rect 19484 114628 19490 114640
rect 19484 114600 20024 114628
rect 19484 114588 19490 114600
rect 18966 114520 18972 114572
rect 19024 114560 19030 114572
rect 19996 114569 20024 114600
rect 20088 114600 21680 114628
rect 19521 114563 19579 114569
rect 19521 114560 19533 114563
rect 19024 114532 19533 114560
rect 19024 114520 19030 114532
rect 19521 114529 19533 114532
rect 19567 114529 19579 114563
rect 19521 114523 19579 114529
rect 19981 114563 20039 114569
rect 19981 114529 19993 114563
rect 20027 114529 20039 114563
rect 19981 114523 20039 114529
rect 20088 114492 20116 114600
rect 20254 114520 20260 114572
rect 20312 114560 20318 114572
rect 20898 114560 20904 114572
rect 20312 114532 20904 114560
rect 20312 114520 20318 114532
rect 20898 114520 20904 114532
rect 20956 114520 20962 114572
rect 21652 114569 21680 114600
rect 21818 114588 21824 114640
rect 21876 114628 21882 114640
rect 22186 114628 22192 114640
rect 21876 114600 22192 114628
rect 21876 114588 21882 114600
rect 22186 114588 22192 114600
rect 22244 114588 22250 114640
rect 22278 114588 22284 114640
rect 22336 114628 22342 114640
rect 22336 114600 23244 114628
rect 22336 114588 22342 114600
rect 20993 114563 21051 114569
rect 20993 114529 21005 114563
rect 21039 114529 21051 114563
rect 20993 114523 21051 114529
rect 21637 114563 21695 114569
rect 21637 114529 21649 114563
rect 21683 114529 21695 114563
rect 22738 114560 22744 114572
rect 22699 114532 22744 114560
rect 21637 114523 21695 114529
rect 18892 114464 20116 114492
rect 20714 114452 20720 114504
rect 20772 114492 20778 114504
rect 21008 114492 21036 114523
rect 22738 114520 22744 114532
rect 22796 114520 22802 114572
rect 23216 114569 23244 114600
rect 23201 114563 23259 114569
rect 23201 114529 23213 114563
rect 23247 114529 23259 114563
rect 23201 114523 23259 114529
rect 23842 114520 23848 114572
rect 23900 114560 23906 114572
rect 24228 114569 24256 114668
rect 27890 114656 27896 114668
rect 27948 114656 27954 114708
rect 27985 114699 28043 114705
rect 27985 114665 27997 114699
rect 28031 114665 28043 114699
rect 27985 114659 28043 114665
rect 28000 114628 28028 114659
rect 29086 114656 29092 114708
rect 29144 114696 29150 114708
rect 29273 114699 29331 114705
rect 29273 114696 29285 114699
rect 29144 114668 29285 114696
rect 29144 114656 29150 114668
rect 29273 114665 29285 114668
rect 29319 114665 29331 114699
rect 29273 114659 29331 114665
rect 29546 114656 29552 114708
rect 29604 114696 29610 114708
rect 30561 114699 30619 114705
rect 30561 114696 30573 114699
rect 29604 114668 30573 114696
rect 29604 114656 29610 114668
rect 30561 114665 30573 114668
rect 30607 114665 30619 114699
rect 30561 114659 30619 114665
rect 30926 114656 30932 114708
rect 30984 114696 30990 114708
rect 31941 114699 31999 114705
rect 31941 114696 31953 114699
rect 30984 114668 31953 114696
rect 30984 114656 30990 114668
rect 31941 114665 31953 114668
rect 31987 114665 31999 114699
rect 31941 114659 31999 114665
rect 25792 114600 28028 114628
rect 25792 114569 25820 114600
rect 28626 114588 28632 114640
rect 28684 114628 28690 114640
rect 28684 114600 29500 114628
rect 28684 114588 28690 114600
rect 24213 114563 24271 114569
rect 23900 114532 24164 114560
rect 23900 114520 23906 114532
rect 20772 114464 21036 114492
rect 24136 114492 24164 114532
rect 24213 114529 24225 114563
rect 24259 114529 24271 114563
rect 25133 114563 25191 114569
rect 24213 114523 24271 114529
rect 24320 114532 24854 114560
rect 24320 114492 24348 114532
rect 24136 114464 24348 114492
rect 20772 114452 20778 114464
rect 8294 114384 8300 114436
rect 8352 114424 8358 114436
rect 12069 114427 12127 114433
rect 12069 114424 12081 114427
rect 8352 114396 12081 114424
rect 8352 114384 8358 114396
rect 12069 114393 12081 114396
rect 12115 114393 12127 114427
rect 15286 114424 15292 114436
rect 15247 114396 15292 114424
rect 12069 114387 12127 114393
rect 15286 114384 15292 114396
rect 15344 114384 15350 114436
rect 18874 114424 18880 114436
rect 18835 114396 18880 114424
rect 18874 114384 18880 114396
rect 18932 114384 18938 114436
rect 19334 114424 19340 114436
rect 19295 114396 19340 114424
rect 19334 114384 19340 114396
rect 19392 114384 19398 114436
rect 24826 114424 24854 114532
rect 25133 114529 25145 114563
rect 25179 114529 25191 114563
rect 25133 114523 25191 114529
rect 25777 114563 25835 114569
rect 25777 114529 25789 114563
rect 25823 114529 25835 114563
rect 26418 114560 26424 114572
rect 26379 114532 26424 114560
rect 25777 114523 25835 114529
rect 25148 114492 25176 114523
rect 26418 114520 26424 114532
rect 26476 114520 26482 114572
rect 27982 114520 27988 114572
rect 28040 114560 28046 114572
rect 28169 114563 28227 114569
rect 28169 114560 28181 114563
rect 28040 114532 28181 114560
rect 28040 114520 28046 114532
rect 28169 114529 28181 114532
rect 28215 114529 28227 114563
rect 28169 114523 28227 114529
rect 28442 114520 28448 114572
rect 28500 114560 28506 114572
rect 29472 114569 29500 114600
rect 29914 114588 29920 114640
rect 29972 114628 29978 114640
rect 32766 114628 32772 114640
rect 29972 114600 30788 114628
rect 29972 114588 29978 114600
rect 28813 114563 28871 114569
rect 28813 114560 28825 114563
rect 28500 114532 28825 114560
rect 28500 114520 28506 114532
rect 28813 114529 28825 114532
rect 28859 114529 28871 114563
rect 28813 114523 28871 114529
rect 29457 114563 29515 114569
rect 29457 114529 29469 114563
rect 29503 114529 29515 114563
rect 29457 114523 29515 114529
rect 30006 114520 30012 114572
rect 30064 114560 30070 114572
rect 30101 114563 30159 114569
rect 30101 114560 30113 114563
rect 30064 114532 30113 114560
rect 30064 114520 30070 114532
rect 30101 114529 30113 114532
rect 30147 114529 30159 114563
rect 30101 114523 30159 114529
rect 30282 114520 30288 114572
rect 30340 114560 30346 114572
rect 30760 114569 30788 114600
rect 31496 114600 32772 114628
rect 30745 114563 30803 114569
rect 30340 114532 30696 114560
rect 30340 114520 30346 114532
rect 30466 114492 30472 114504
rect 25148 114464 30472 114492
rect 30466 114452 30472 114464
rect 30524 114452 30530 114504
rect 30668 114492 30696 114532
rect 30745 114529 30757 114563
rect 30791 114529 30803 114563
rect 30745 114523 30803 114529
rect 31389 114563 31447 114569
rect 31389 114529 31401 114563
rect 31435 114529 31447 114563
rect 31389 114523 31447 114529
rect 31404 114492 31432 114523
rect 30668 114464 31432 114492
rect 24949 114427 25007 114433
rect 24949 114424 24961 114427
rect 24826 114396 24961 114424
rect 24949 114393 24961 114396
rect 24995 114393 25007 114427
rect 24949 114387 25007 114393
rect 25314 114384 25320 114436
rect 25372 114424 25378 114436
rect 25593 114427 25651 114433
rect 25593 114424 25605 114427
rect 25372 114396 25605 114424
rect 25372 114384 25378 114396
rect 25593 114393 25605 114396
rect 25639 114393 25651 114427
rect 26234 114424 26240 114436
rect 26195 114396 26240 114424
rect 25593 114387 25651 114393
rect 26234 114384 26240 114396
rect 26292 114384 26298 114436
rect 26694 114384 26700 114436
rect 26752 114424 26758 114436
rect 29917 114427 29975 114433
rect 29917 114424 29929 114427
rect 26752 114396 29929 114424
rect 26752 114384 26758 114396
rect 29917 114393 29929 114396
rect 29963 114393 29975 114427
rect 29917 114387 29975 114393
rect 30190 114384 30196 114436
rect 30248 114424 30254 114436
rect 31205 114427 31263 114433
rect 31205 114424 31217 114427
rect 30248 114396 31217 114424
rect 30248 114384 30254 114396
rect 31205 114393 31217 114396
rect 31251 114393 31263 114427
rect 31205 114387 31263 114393
rect 9033 114359 9091 114365
rect 9033 114356 9045 114359
rect 8128 114328 9045 114356
rect 5721 114319 5779 114325
rect 9033 114325 9045 114328
rect 9079 114325 9091 114359
rect 9858 114356 9864 114368
rect 9819 114328 9864 114356
rect 9033 114319 9091 114325
rect 9858 114316 9864 114328
rect 9916 114316 9922 114368
rect 10962 114356 10968 114368
rect 10923 114328 10968 114356
rect 10962 114316 10968 114328
rect 11020 114316 11026 114368
rect 13354 114356 13360 114368
rect 13315 114328 13360 114356
rect 13354 114316 13360 114328
rect 13412 114316 13418 114368
rect 14642 114356 14648 114368
rect 14603 114328 14648 114356
rect 14642 114316 14648 114328
rect 14700 114316 14706 114368
rect 28626 114356 28632 114368
rect 28587 114328 28632 114356
rect 28626 114316 28632 114328
rect 28684 114316 28690 114368
rect 30282 114316 30288 114368
rect 30340 114356 30346 114368
rect 31496 114356 31524 114600
rect 32766 114588 32772 114600
rect 32824 114588 32830 114640
rect 34146 114588 34152 114640
rect 34204 114628 34210 114640
rect 35713 114631 35771 114637
rect 35713 114628 35725 114631
rect 34204 114600 35725 114628
rect 34204 114588 34210 114600
rect 35713 114597 35725 114600
rect 35759 114597 35771 114631
rect 35713 114591 35771 114597
rect 35897 114631 35955 114637
rect 35897 114597 35909 114631
rect 35943 114628 35955 114631
rect 39206 114628 39212 114640
rect 35943 114600 39212 114628
rect 35943 114597 35955 114600
rect 35897 114591 35955 114597
rect 39206 114588 39212 114600
rect 39264 114588 39270 114640
rect 32125 114563 32183 114569
rect 32125 114529 32137 114563
rect 32171 114560 32183 114563
rect 32214 114560 32220 114572
rect 32171 114532 32220 114560
rect 32171 114529 32183 114532
rect 32125 114523 32183 114529
rect 32214 114520 32220 114532
rect 32272 114520 32278 114572
rect 33226 114520 33232 114572
rect 33284 114560 33290 114572
rect 33505 114563 33563 114569
rect 33505 114560 33517 114563
rect 33284 114532 33517 114560
rect 33284 114520 33290 114532
rect 33505 114529 33517 114532
rect 33551 114529 33563 114563
rect 34241 114563 34299 114569
rect 34241 114560 34253 114563
rect 33505 114523 33563 114529
rect 33612 114532 34253 114560
rect 32766 114452 32772 114504
rect 32824 114492 32830 114504
rect 33612 114492 33640 114532
rect 34241 114529 34253 114532
rect 34287 114529 34299 114563
rect 34241 114523 34299 114529
rect 34790 114520 34796 114572
rect 34848 114560 34854 114572
rect 34977 114563 35035 114569
rect 34977 114560 34989 114563
rect 34848 114532 34989 114560
rect 34848 114520 34854 114532
rect 34977 114529 34989 114532
rect 35023 114529 35035 114563
rect 34977 114523 35035 114529
rect 36170 114520 36176 114572
rect 36228 114560 36234 114572
rect 36449 114563 36507 114569
rect 36449 114560 36461 114563
rect 36228 114532 36461 114560
rect 36228 114520 36234 114532
rect 36449 114529 36461 114532
rect 36495 114529 36507 114563
rect 37090 114560 37096 114572
rect 36449 114523 36507 114529
rect 36556 114532 36860 114560
rect 37051 114532 37096 114560
rect 32824 114464 33640 114492
rect 33689 114495 33747 114501
rect 32824 114452 32830 114464
rect 33689 114461 33701 114495
rect 33735 114492 33747 114495
rect 35066 114492 35072 114504
rect 33735 114464 35072 114492
rect 33735 114461 33747 114464
rect 33689 114455 33747 114461
rect 35066 114452 35072 114464
rect 35124 114452 35130 114504
rect 35161 114495 35219 114501
rect 35161 114461 35173 114495
rect 35207 114492 35219 114495
rect 36556 114492 36584 114532
rect 35207 114464 36584 114492
rect 36633 114495 36691 114501
rect 35207 114461 35219 114464
rect 35161 114455 35219 114461
rect 36633 114461 36645 114495
rect 36679 114492 36691 114495
rect 36722 114492 36728 114504
rect 36679 114464 36728 114492
rect 36679 114461 36691 114464
rect 36633 114455 36691 114461
rect 36722 114452 36728 114464
rect 36780 114452 36786 114504
rect 36832 114492 36860 114532
rect 37090 114520 37096 114532
rect 37148 114520 37154 114572
rect 39666 114492 39672 114504
rect 36832 114464 39672 114492
rect 39666 114452 39672 114464
rect 39724 114452 39730 114504
rect 34425 114427 34483 114433
rect 34425 114393 34437 114427
rect 34471 114424 34483 114427
rect 37366 114424 37372 114436
rect 34471 114396 37372 114424
rect 34471 114393 34483 114396
rect 34425 114387 34483 114393
rect 37366 114384 37372 114396
rect 37424 114384 37430 114436
rect 37274 114356 37280 114368
rect 30340 114328 31524 114356
rect 37235 114328 37280 114356
rect 30340 114316 30346 114328
rect 37274 114316 37280 114328
rect 37332 114316 37338 114368
rect 1104 114266 38824 114288
rect 1104 114214 4246 114266
rect 4298 114214 4310 114266
rect 4362 114214 4374 114266
rect 4426 114214 4438 114266
rect 4490 114214 34966 114266
rect 35018 114214 35030 114266
rect 35082 114214 35094 114266
rect 35146 114214 35158 114266
rect 35210 114214 38824 114266
rect 1104 114192 38824 114214
rect 2590 114112 2596 114164
rect 2648 114152 2654 114164
rect 3053 114155 3111 114161
rect 3053 114152 3065 114155
rect 2648 114124 3065 114152
rect 2648 114112 2654 114124
rect 3053 114121 3065 114124
rect 3099 114121 3111 114155
rect 3053 114115 3111 114121
rect 4433 114155 4491 114161
rect 4433 114121 4445 114155
rect 4479 114152 4491 114155
rect 4614 114152 4620 114164
rect 4479 114124 4620 114152
rect 4479 114121 4491 114124
rect 4433 114115 4491 114121
rect 4614 114112 4620 114124
rect 4672 114112 4678 114164
rect 5626 114112 5632 114164
rect 5684 114152 5690 114164
rect 5813 114155 5871 114161
rect 5813 114152 5825 114155
rect 5684 114124 5825 114152
rect 5684 114112 5690 114124
rect 5813 114121 5825 114124
rect 5859 114121 5871 114155
rect 5813 114115 5871 114121
rect 7009 114155 7067 114161
rect 7009 114121 7021 114155
rect 7055 114152 7067 114155
rect 7742 114152 7748 114164
rect 7055 114124 7748 114152
rect 7055 114121 7067 114124
rect 7009 114115 7067 114121
rect 7742 114112 7748 114124
rect 7800 114112 7806 114164
rect 9493 114155 9551 114161
rect 9493 114121 9505 114155
rect 9539 114152 9551 114155
rect 18046 114152 18052 114164
rect 9539 114124 18052 114152
rect 9539 114121 9551 114124
rect 9493 114115 9551 114121
rect 18046 114112 18052 114124
rect 18104 114112 18110 114164
rect 18325 114155 18383 114161
rect 18325 114121 18337 114155
rect 18371 114152 18383 114155
rect 20254 114152 20260 114164
rect 18371 114124 20260 114152
rect 18371 114121 18383 114124
rect 18325 114115 18383 114121
rect 20254 114112 20260 114124
rect 20312 114112 20318 114164
rect 21545 114155 21603 114161
rect 21545 114121 21557 114155
rect 21591 114152 21603 114155
rect 24486 114152 24492 114164
rect 21591 114124 24492 114152
rect 21591 114121 21603 114124
rect 21545 114115 21603 114121
rect 24486 114112 24492 114124
rect 24544 114112 24550 114164
rect 25225 114155 25283 114161
rect 25225 114121 25237 114155
rect 25271 114152 25283 114155
rect 25406 114152 25412 114164
rect 25271 114124 25412 114152
rect 25271 114121 25283 114124
rect 25225 114115 25283 114121
rect 25406 114112 25412 114124
rect 25464 114112 25470 114164
rect 25590 114112 25596 114164
rect 25648 114152 25654 114164
rect 26237 114155 26295 114161
rect 26237 114152 26249 114155
rect 25648 114124 26249 114152
rect 25648 114112 25654 114124
rect 26237 114121 26249 114124
rect 26283 114121 26295 114155
rect 26237 114115 26295 114121
rect 28718 114112 28724 114164
rect 28776 114152 28782 114164
rect 29273 114155 29331 114161
rect 29273 114152 29285 114155
rect 28776 114124 29285 114152
rect 28776 114112 28782 114124
rect 29273 114121 29285 114124
rect 29319 114121 29331 114155
rect 29273 114115 29331 114121
rect 29638 114112 29644 114164
rect 29696 114152 29702 114164
rect 30469 114155 30527 114161
rect 30469 114152 30481 114155
rect 29696 114124 30481 114152
rect 29696 114112 29702 114124
rect 30469 114121 30481 114124
rect 30515 114121 30527 114155
rect 30469 114115 30527 114121
rect 31478 114112 31484 114164
rect 31536 114152 31542 114164
rect 31757 114155 31815 114161
rect 31757 114152 31769 114155
rect 31536 114124 31769 114152
rect 31536 114112 31542 114124
rect 31757 114121 31769 114124
rect 31803 114121 31815 114155
rect 31757 114115 31815 114121
rect 31938 114112 31944 114164
rect 31996 114152 32002 114164
rect 32493 114155 32551 114161
rect 32493 114152 32505 114155
rect 31996 114124 32505 114152
rect 31996 114112 32002 114124
rect 32493 114121 32505 114124
rect 32539 114121 32551 114155
rect 32493 114115 32551 114121
rect 32858 114112 32864 114164
rect 32916 114152 32922 114164
rect 33689 114155 33747 114161
rect 33689 114152 33701 114155
rect 32916 114124 33701 114152
rect 32916 114112 32922 114124
rect 33689 114121 33701 114124
rect 33735 114121 33747 114155
rect 33689 114115 33747 114121
rect 34701 114155 34759 114161
rect 34701 114121 34713 114155
rect 34747 114152 34759 114155
rect 34747 114124 36952 114152
rect 34747 114121 34759 114124
rect 34701 114115 34759 114121
rect 3602 114044 3608 114096
rect 3660 114084 3666 114096
rect 5077 114087 5135 114093
rect 5077 114084 5089 114087
rect 3660 114056 5089 114084
rect 3660 114044 3666 114056
rect 5077 114053 5089 114056
rect 5123 114053 5135 114087
rect 5077 114047 5135 114053
rect 5442 114044 5448 114096
rect 5500 114084 5506 114096
rect 8113 114087 8171 114093
rect 8113 114084 8125 114087
rect 5500 114056 8125 114084
rect 5500 114044 5506 114056
rect 8113 114053 8125 114056
rect 8159 114053 8171 114087
rect 8113 114047 8171 114053
rect 15749 114087 15807 114093
rect 15749 114053 15761 114087
rect 15795 114053 15807 114087
rect 15749 114047 15807 114053
rect 17681 114087 17739 114093
rect 17681 114053 17693 114087
rect 17727 114084 17739 114087
rect 22738 114084 22744 114096
rect 17727 114056 22744 114084
rect 17727 114053 17739 114056
rect 17681 114047 17739 114053
rect 10410 114016 10416 114028
rect 8312 113988 10416 114016
rect 8312 113957 8340 113988
rect 10410 113976 10416 113988
rect 10468 113976 10474 114028
rect 15764 114016 15792 114047
rect 22738 114044 22744 114056
rect 22796 114044 22802 114096
rect 29362 114044 29368 114096
rect 29420 114084 29426 114096
rect 31113 114087 31171 114093
rect 31113 114084 31125 114087
rect 29420 114056 31125 114084
rect 29420 114044 29426 114056
rect 31113 114053 31125 114056
rect 31159 114053 31171 114087
rect 31113 114047 31171 114053
rect 36633 114087 36691 114093
rect 36633 114053 36645 114087
rect 36679 114084 36691 114087
rect 36814 114084 36820 114096
rect 36679 114056 36820 114084
rect 36679 114053 36691 114056
rect 36633 114047 36691 114053
rect 36814 114044 36820 114056
rect 36872 114044 36878 114096
rect 36924 114084 36952 114124
rect 37182 114112 37188 114164
rect 37240 114152 37246 114164
rect 38013 114155 38071 114161
rect 38013 114152 38025 114155
rect 37240 114124 38025 114152
rect 37240 114112 37246 114124
rect 38013 114121 38025 114124
rect 38059 114121 38071 114155
rect 38013 114115 38071 114121
rect 38378 114084 38384 114096
rect 36924 114056 38384 114084
rect 38378 114044 38384 114056
rect 38436 114044 38442 114096
rect 20714 114016 20720 114028
rect 15764 113988 20720 114016
rect 20714 113976 20720 113988
rect 20772 113976 20778 114028
rect 30374 113976 30380 114028
rect 30432 114016 30438 114028
rect 33042 114016 33048 114028
rect 30432 113988 31340 114016
rect 30432 113976 30438 113988
rect 7653 113951 7711 113957
rect 7653 113917 7665 113951
rect 7699 113917 7711 113951
rect 7653 113911 7711 113917
rect 8297 113951 8355 113957
rect 8297 113917 8309 113951
rect 8343 113917 8355 113951
rect 8297 113911 8355 113917
rect 1857 113883 1915 113889
rect 1857 113849 1869 113883
rect 1903 113880 1915 113883
rect 2130 113880 2136 113892
rect 1903 113852 2136 113880
rect 1903 113849 1915 113852
rect 1857 113843 1915 113849
rect 2130 113840 2136 113852
rect 2188 113840 2194 113892
rect 7668 113880 7696 113911
rect 8754 113908 8760 113960
rect 8812 113948 8818 113960
rect 9677 113951 9735 113957
rect 9677 113948 9689 113951
rect 8812 113920 9689 113948
rect 8812 113908 8818 113920
rect 9677 113917 9689 113920
rect 9723 113917 9735 113951
rect 9677 113911 9735 113917
rect 15746 113908 15752 113960
rect 15804 113948 15810 113960
rect 15933 113951 15991 113957
rect 15933 113948 15945 113951
rect 15804 113920 15945 113948
rect 15804 113908 15810 113920
rect 15933 113917 15945 113920
rect 15979 113917 15991 113951
rect 15933 113911 15991 113917
rect 16482 113908 16488 113960
rect 16540 113948 16546 113960
rect 16577 113951 16635 113957
rect 16577 113948 16589 113951
rect 16540 113920 16589 113948
rect 16540 113908 16546 113920
rect 16577 113917 16589 113920
rect 16623 113917 16635 113951
rect 16577 113911 16635 113917
rect 17678 113908 17684 113960
rect 17736 113948 17742 113960
rect 17865 113951 17923 113957
rect 17865 113948 17877 113951
rect 17736 113920 17877 113948
rect 17736 113908 17742 113920
rect 17865 113917 17877 113920
rect 17911 113917 17923 113951
rect 17865 113911 17923 113917
rect 18230 113908 18236 113960
rect 18288 113948 18294 113960
rect 18509 113951 18567 113957
rect 18509 113948 18521 113951
rect 18288 113920 18521 113948
rect 18288 113908 18294 113920
rect 18509 113917 18521 113920
rect 18555 113917 18567 113951
rect 20162 113948 20168 113960
rect 20123 113920 20168 113948
rect 18509 113911 18567 113917
rect 20162 113908 20168 113920
rect 20220 113908 20226 113960
rect 20806 113948 20812 113960
rect 20767 113920 20812 113948
rect 20806 113908 20812 113920
rect 20864 113908 20870 113960
rect 21729 113951 21787 113957
rect 21729 113917 21741 113951
rect 21775 113917 21787 113951
rect 22186 113948 22192 113960
rect 22147 113920 22192 113948
rect 21729 113911 21787 113917
rect 8386 113880 8392 113892
rect 7668 113852 8392 113880
rect 8386 113840 8392 113852
rect 8444 113840 8450 113892
rect 21744 113880 21772 113911
rect 22186 113908 22192 113920
rect 22244 113908 22250 113960
rect 22830 113948 22836 113960
rect 22791 113920 22836 113948
rect 22830 113908 22836 113920
rect 22888 113908 22894 113960
rect 23382 113908 23388 113960
rect 23440 113948 23446 113960
rect 23477 113951 23535 113957
rect 23477 113948 23489 113951
rect 23440 113920 23489 113948
rect 23440 113908 23446 113920
rect 23477 113917 23489 113920
rect 23523 113917 23535 113951
rect 23477 113911 23535 113917
rect 24026 113908 24032 113960
rect 24084 113948 24090 113960
rect 24121 113951 24179 113957
rect 24121 113948 24133 113951
rect 24084 113920 24133 113948
rect 24084 113908 24090 113920
rect 24121 113917 24133 113920
rect 24167 113917 24179 113951
rect 24121 113911 24179 113917
rect 25409 113951 25467 113957
rect 25409 113917 25421 113951
rect 25455 113948 25467 113951
rect 26142 113948 26148 113960
rect 25455 113920 26148 113948
rect 25455 113917 25467 113920
rect 25409 113911 25467 113917
rect 26142 113908 26148 113920
rect 26200 113908 26206 113960
rect 26421 113951 26479 113957
rect 26421 113917 26433 113951
rect 26467 113948 26479 113951
rect 28626 113948 28632 113960
rect 26467 113920 28632 113948
rect 26467 113917 26479 113920
rect 26421 113911 26479 113917
rect 28626 113908 28632 113920
rect 28684 113908 28690 113960
rect 29270 113908 29276 113960
rect 29328 113948 29334 113960
rect 29457 113951 29515 113957
rect 29457 113948 29469 113951
rect 29328 113920 29469 113948
rect 29328 113908 29334 113920
rect 29457 113917 29469 113920
rect 29503 113917 29515 113951
rect 29457 113911 29515 113917
rect 30098 113908 30104 113960
rect 30156 113948 30162 113960
rect 31312 113957 31340 113988
rect 31956 113988 33048 114016
rect 31956 113957 31984 113988
rect 33042 113976 33048 113988
rect 33100 113976 33106 114028
rect 33962 113976 33968 114028
rect 34020 114016 34026 114028
rect 35802 114016 35808 114028
rect 34020 113988 35808 114016
rect 34020 113976 34026 113988
rect 35802 113976 35808 113988
rect 35860 113976 35866 114028
rect 37366 114016 37372 114028
rect 37327 113988 37372 114016
rect 37366 113976 37372 113988
rect 37424 113976 37430 114028
rect 30653 113951 30711 113957
rect 30653 113948 30665 113951
rect 30156 113920 30665 113948
rect 30156 113908 30162 113920
rect 30653 113917 30665 113920
rect 30699 113917 30711 113951
rect 30653 113911 30711 113917
rect 31297 113951 31355 113957
rect 31297 113917 31309 113951
rect 31343 113917 31355 113951
rect 31297 113911 31355 113917
rect 31941 113951 31999 113957
rect 31941 113917 31953 113951
rect 31987 113917 31999 113951
rect 31941 113911 31999 113917
rect 32490 113908 32496 113960
rect 32548 113948 32554 113960
rect 32677 113951 32735 113957
rect 32677 113948 32689 113951
rect 32548 113920 32689 113948
rect 32548 113908 32554 113920
rect 32677 113917 32689 113920
rect 32723 113917 32735 113951
rect 32677 113911 32735 113917
rect 33686 113908 33692 113960
rect 33744 113948 33750 113960
rect 33873 113951 33931 113957
rect 33873 113948 33885 113951
rect 33744 113920 33885 113948
rect 33744 113908 33750 113920
rect 33873 113917 33885 113920
rect 33919 113917 33931 113951
rect 33873 113911 33931 113917
rect 35526 113908 35532 113960
rect 35584 113948 35590 113960
rect 37185 113951 37243 113957
rect 37185 113948 37197 113951
rect 35584 113920 37197 113948
rect 35584 113908 35590 113920
rect 37185 113917 37197 113920
rect 37231 113917 37243 113951
rect 37185 113911 37243 113917
rect 16408 113852 21772 113880
rect 1946 113812 1952 113824
rect 1907 113784 1952 113812
rect 1946 113772 1952 113784
rect 2004 113772 2010 113824
rect 3878 113772 3884 113824
rect 3936 113812 3942 113824
rect 16408 113821 16436 113852
rect 31570 113840 31576 113892
rect 31628 113880 31634 113892
rect 34609 113883 34667 113889
rect 34609 113880 34621 113883
rect 31628 113852 34621 113880
rect 31628 113840 31634 113852
rect 34609 113849 34621 113852
rect 34655 113849 34667 113883
rect 34609 113843 34667 113849
rect 35342 113840 35348 113892
rect 35400 113880 35406 113892
rect 36449 113883 36507 113889
rect 36449 113880 36461 113883
rect 35400 113852 36461 113880
rect 35400 113840 35406 113852
rect 36449 113849 36461 113852
rect 36495 113849 36507 113883
rect 36449 113843 36507 113849
rect 37458 113840 37464 113892
rect 37516 113880 37522 113892
rect 37921 113883 37979 113889
rect 37921 113880 37933 113883
rect 37516 113852 37933 113880
rect 37516 113840 37522 113852
rect 37921 113849 37933 113852
rect 37967 113849 37979 113883
rect 37921 113843 37979 113849
rect 7469 113815 7527 113821
rect 7469 113812 7481 113815
rect 3936 113784 7481 113812
rect 3936 113772 3942 113784
rect 7469 113781 7481 113784
rect 7515 113781 7527 113815
rect 7469 113775 7527 113781
rect 16393 113815 16451 113821
rect 16393 113781 16405 113815
rect 16439 113781 16451 113815
rect 16393 113775 16451 113781
rect 25406 113772 25412 113824
rect 25464 113812 25470 113824
rect 34054 113812 34060 113824
rect 25464 113784 34060 113812
rect 25464 113772 25470 113784
rect 34054 113772 34060 113784
rect 34112 113772 34118 113824
rect 1104 113722 38824 113744
rect 1104 113670 19606 113722
rect 19658 113670 19670 113722
rect 19722 113670 19734 113722
rect 19786 113670 19798 113722
rect 19850 113670 38824 113722
rect 1104 113648 38824 113670
rect 4617 113611 4675 113617
rect 4617 113577 4629 113611
rect 4663 113608 4675 113611
rect 5166 113608 5172 113620
rect 4663 113580 5172 113608
rect 4663 113577 4675 113580
rect 4617 113571 4675 113577
rect 5166 113568 5172 113580
rect 5224 113568 5230 113620
rect 5258 113568 5264 113620
rect 5316 113608 5322 113620
rect 6825 113611 6883 113617
rect 6825 113608 6837 113611
rect 5316 113580 6837 113608
rect 5316 113568 5322 113580
rect 6825 113577 6837 113580
rect 6871 113577 6883 113611
rect 8294 113608 8300 113620
rect 6825 113571 6883 113577
rect 7024 113580 8300 113608
rect 6638 113540 6644 113552
rect 4816 113512 6644 113540
rect 1489 113475 1547 113481
rect 1489 113441 1501 113475
rect 1535 113472 1547 113475
rect 1762 113472 1768 113484
rect 1535 113444 1768 113472
rect 1535 113441 1547 113444
rect 1489 113435 1547 113441
rect 1762 113432 1768 113444
rect 1820 113432 1826 113484
rect 2314 113472 2320 113484
rect 2275 113444 2320 113472
rect 2314 113432 2320 113444
rect 2372 113432 2378 113484
rect 2961 113475 3019 113481
rect 2961 113441 2973 113475
rect 3007 113472 3019 113475
rect 3050 113472 3056 113484
rect 3007 113444 3056 113472
rect 3007 113441 3019 113444
rect 2961 113435 3019 113441
rect 3050 113432 3056 113444
rect 3108 113432 3114 113484
rect 3142 113432 3148 113484
rect 3200 113472 3206 113484
rect 4816 113481 4844 113512
rect 6638 113500 6644 113512
rect 6696 113500 6702 113552
rect 3421 113475 3479 113481
rect 3421 113472 3433 113475
rect 3200 113444 3433 113472
rect 3200 113432 3206 113444
rect 3421 113441 3433 113444
rect 3467 113441 3479 113475
rect 3421 113435 3479 113441
rect 4801 113475 4859 113481
rect 4801 113441 4813 113475
rect 4847 113441 4859 113475
rect 4801 113435 4859 113441
rect 5445 113475 5503 113481
rect 5445 113441 5457 113475
rect 5491 113472 5503 113475
rect 6270 113472 6276 113484
rect 5491 113444 6276 113472
rect 5491 113441 5503 113444
rect 5445 113435 5503 113441
rect 6270 113432 6276 113444
rect 6328 113432 6334 113484
rect 7024 113481 7052 113580
rect 8294 113568 8300 113580
rect 8352 113568 8358 113620
rect 30742 113608 30748 113620
rect 30703 113580 30748 113608
rect 30742 113568 30748 113580
rect 30800 113568 30806 113620
rect 32674 113568 32680 113620
rect 32732 113608 32738 113620
rect 33045 113611 33103 113617
rect 33045 113608 33057 113611
rect 32732 113580 33057 113608
rect 32732 113568 32738 113580
rect 33045 113577 33057 113580
rect 33091 113577 33103 113611
rect 33045 113571 33103 113577
rect 35069 113611 35127 113617
rect 35069 113577 35081 113611
rect 35115 113608 35127 113611
rect 38562 113608 38568 113620
rect 35115 113580 38568 113608
rect 35115 113577 35127 113580
rect 35069 113571 35127 113577
rect 38562 113568 38568 113580
rect 38620 113568 38626 113620
rect 7466 113500 7472 113552
rect 7524 113540 7530 113552
rect 8202 113540 8208 113552
rect 7524 113512 8208 113540
rect 7524 113500 7530 113512
rect 8202 113500 8208 113512
rect 8260 113500 8266 113552
rect 14642 113540 14648 113552
rect 8312 113512 14648 113540
rect 8312 113481 8340 113512
rect 14642 113500 14648 113512
rect 14700 113500 14706 113552
rect 35897 113543 35955 113549
rect 35897 113509 35909 113543
rect 35943 113540 35955 113543
rect 36354 113540 36360 113552
rect 35943 113512 36360 113540
rect 35943 113509 35955 113512
rect 35897 113503 35955 113509
rect 36354 113500 36360 113512
rect 36412 113500 36418 113552
rect 36633 113543 36691 113549
rect 36633 113509 36645 113543
rect 36679 113540 36691 113543
rect 36998 113540 37004 113552
rect 36679 113512 37004 113540
rect 36679 113509 36691 113512
rect 36633 113503 36691 113509
rect 36998 113500 37004 113512
rect 37056 113500 37062 113552
rect 7009 113475 7067 113481
rect 7009 113441 7021 113475
rect 7055 113441 7067 113475
rect 7009 113435 7067 113441
rect 7653 113475 7711 113481
rect 7653 113441 7665 113475
rect 7699 113441 7711 113475
rect 7653 113435 7711 113441
rect 8289 113475 8347 113481
rect 8289 113441 8301 113475
rect 8335 113441 8347 113475
rect 8289 113435 8347 113441
rect 7668 113404 7696 113435
rect 8386 113432 8392 113484
rect 8444 113472 8450 113484
rect 8757 113475 8815 113481
rect 8757 113472 8769 113475
rect 8444 113444 8769 113472
rect 8444 113432 8450 113444
rect 8757 113441 8769 113444
rect 8803 113441 8815 113475
rect 24578 113472 24584 113484
rect 24539 113444 24584 113472
rect 8757 113435 8815 113441
rect 24578 113432 24584 113444
rect 24636 113432 24642 113484
rect 25222 113472 25228 113484
rect 25183 113444 25228 113472
rect 25222 113432 25228 113444
rect 25280 113432 25286 113484
rect 30834 113432 30840 113484
rect 30892 113472 30898 113484
rect 30929 113475 30987 113481
rect 30929 113472 30941 113475
rect 30892 113444 30941 113472
rect 30892 113432 30898 113444
rect 30929 113441 30941 113444
rect 30975 113441 30987 113475
rect 30929 113435 30987 113441
rect 31294 113432 31300 113484
rect 31352 113472 31358 113484
rect 31573 113475 31631 113481
rect 31573 113472 31585 113475
rect 31352 113444 31585 113472
rect 31352 113432 31358 113444
rect 31573 113441 31585 113444
rect 31619 113441 31631 113475
rect 31573 113435 31631 113441
rect 32950 113432 32956 113484
rect 33008 113472 33014 113484
rect 33229 113475 33287 113481
rect 33229 113472 33241 113475
rect 33008 113444 33241 113472
rect 33008 113432 33014 113444
rect 33229 113441 33241 113444
rect 33275 113441 33287 113475
rect 33229 113435 33287 113441
rect 33594 113432 33600 113484
rect 33652 113472 33658 113484
rect 33873 113475 33931 113481
rect 33873 113472 33885 113475
rect 33652 113444 33885 113472
rect 33652 113432 33658 113444
rect 33873 113441 33885 113444
rect 33919 113441 33931 113475
rect 33873 113435 33931 113441
rect 34514 113432 34520 113484
rect 34572 113472 34578 113484
rect 34977 113475 35035 113481
rect 34977 113472 34989 113475
rect 34572 113444 34989 113472
rect 34572 113432 34578 113444
rect 34977 113441 34989 113444
rect 35023 113441 35035 113475
rect 35710 113472 35716 113484
rect 35671 113444 35716 113472
rect 34977 113435 35035 113441
rect 35710 113432 35716 113444
rect 35768 113432 35774 113484
rect 36078 113432 36084 113484
rect 36136 113472 36142 113484
rect 36449 113475 36507 113481
rect 36449 113472 36461 113475
rect 36136 113444 36461 113472
rect 36136 113432 36142 113444
rect 36449 113441 36461 113444
rect 36495 113441 36507 113475
rect 36449 113435 36507 113441
rect 37185 113475 37243 113481
rect 37185 113441 37197 113475
rect 37231 113441 37243 113475
rect 37185 113435 37243 113441
rect 13354 113404 13360 113416
rect 7668 113376 13360 113404
rect 13354 113364 13360 113376
rect 13412 113364 13418 113416
rect 21634 113364 21640 113416
rect 21692 113404 21698 113416
rect 37200 113404 37228 113435
rect 21692 113376 37228 113404
rect 21692 113364 21698 113376
rect 4706 113296 4712 113348
rect 4764 113336 4770 113348
rect 5261 113339 5319 113345
rect 5261 113336 5273 113339
rect 4764 113308 5273 113336
rect 4764 113296 4770 113308
rect 5261 113305 5273 113308
rect 5307 113305 5319 113339
rect 5261 113299 5319 113305
rect 6730 113296 6736 113348
rect 6788 113336 6794 113348
rect 7469 113339 7527 113345
rect 7469 113336 7481 113339
rect 6788 113308 7481 113336
rect 6788 113296 6794 113308
rect 7469 113305 7481 113308
rect 7515 113305 7527 113339
rect 8110 113336 8116 113348
rect 8071 113308 8116 113336
rect 7469 113299 7527 113305
rect 8110 113296 8116 113308
rect 8168 113296 8174 113348
rect 30650 113296 30656 113348
rect 30708 113336 30714 113348
rect 31389 113339 31447 113345
rect 31389 113336 31401 113339
rect 30708 113308 31401 113336
rect 30708 113296 30714 113308
rect 31389 113305 31401 113308
rect 31435 113305 31447 113339
rect 31389 113299 31447 113305
rect 32122 113296 32128 113348
rect 32180 113336 32186 113348
rect 33689 113339 33747 113345
rect 33689 113336 33701 113339
rect 32180 113308 33701 113336
rect 32180 113296 32186 113308
rect 33689 113305 33701 113308
rect 33735 113305 33747 113339
rect 37366 113336 37372 113348
rect 37327 113308 37372 113336
rect 33689 113299 33747 113305
rect 37366 113296 37372 113308
rect 37424 113296 37430 113348
rect 1104 113178 38824 113200
rect 1104 113126 4246 113178
rect 4298 113126 4310 113178
rect 4362 113126 4374 113178
rect 4426 113126 4438 113178
rect 4490 113126 34966 113178
rect 35018 113126 35030 113178
rect 35082 113126 35094 113178
rect 35146 113126 35158 113178
rect 35210 113126 38824 113178
rect 1104 113104 38824 113126
rect 30558 113024 30564 113076
rect 30616 113064 30622 113076
rect 31389 113067 31447 113073
rect 31389 113064 31401 113067
rect 30616 113036 31401 113064
rect 30616 113024 30622 113036
rect 31389 113033 31401 113036
rect 31435 113033 31447 113067
rect 31389 113027 31447 113033
rect 33134 113024 33140 113076
rect 33192 113064 33198 113076
rect 33321 113067 33379 113073
rect 33321 113064 33333 113067
rect 33192 113036 33333 113064
rect 33192 113024 33198 113036
rect 33321 113033 33333 113036
rect 33367 113033 33379 113067
rect 33321 113027 33379 113033
rect 33870 113024 33876 113076
rect 33928 113064 33934 113076
rect 33965 113067 34023 113073
rect 33965 113064 33977 113067
rect 33928 113036 33977 113064
rect 33928 113024 33934 113036
rect 33965 113033 33977 113036
rect 34011 113033 34023 113067
rect 36538 113064 36544 113076
rect 36499 113036 36544 113064
rect 33965 113027 34023 113033
rect 36538 113024 36544 113036
rect 36596 113024 36602 113076
rect 6822 112956 6828 113008
rect 6880 112956 6886 113008
rect 28261 112999 28319 113005
rect 28261 112965 28273 112999
rect 28307 112996 28319 112999
rect 28534 112996 28540 113008
rect 28307 112968 28540 112996
rect 28307 112965 28319 112968
rect 28261 112959 28319 112965
rect 28534 112956 28540 112968
rect 28592 112956 28598 113008
rect 1670 112888 1676 112940
rect 1728 112928 1734 112940
rect 6840 112928 6868 112956
rect 1728 112900 2728 112928
rect 6840 112900 7512 112928
rect 1728 112888 1734 112900
rect 1854 112860 1860 112872
rect 1815 112832 1860 112860
rect 1854 112820 1860 112832
rect 1912 112820 1918 112872
rect 2700 112869 2728 112900
rect 2685 112863 2743 112869
rect 2685 112829 2697 112863
rect 2731 112829 2743 112863
rect 2685 112823 2743 112829
rect 3786 112820 3792 112872
rect 3844 112860 3850 112872
rect 4249 112863 4307 112869
rect 4249 112860 4261 112863
rect 3844 112832 4261 112860
rect 3844 112820 3850 112832
rect 4249 112829 4261 112832
rect 4295 112829 4307 112863
rect 4890 112860 4896 112872
rect 4851 112832 4896 112860
rect 4249 112823 4307 112829
rect 4890 112820 4896 112832
rect 4948 112820 4954 112872
rect 5534 112860 5540 112872
rect 5495 112832 5540 112860
rect 5534 112820 5540 112832
rect 5592 112820 5598 112872
rect 5810 112820 5816 112872
rect 5868 112860 5874 112872
rect 6181 112863 6239 112869
rect 6181 112860 6193 112863
rect 5868 112832 6193 112860
rect 5868 112820 5874 112832
rect 6181 112829 6193 112832
rect 6227 112829 6239 112863
rect 6181 112823 6239 112829
rect 6270 112820 6276 112872
rect 6328 112860 6334 112872
rect 7484 112869 7512 112900
rect 31018 112888 31024 112940
rect 31076 112928 31082 112940
rect 31076 112900 37964 112928
rect 31076 112888 31082 112900
rect 6825 112863 6883 112869
rect 6825 112860 6837 112863
rect 6328 112832 6837 112860
rect 6328 112820 6334 112832
rect 6825 112829 6837 112832
rect 6871 112829 6883 112863
rect 6825 112823 6883 112829
rect 7469 112863 7527 112869
rect 7469 112829 7481 112863
rect 7515 112829 7527 112863
rect 28166 112860 28172 112872
rect 28127 112832 28172 112860
rect 7469 112823 7527 112829
rect 28166 112820 28172 112832
rect 28224 112820 28230 112872
rect 28445 112863 28503 112869
rect 28445 112829 28457 112863
rect 28491 112860 28503 112863
rect 29822 112860 29828 112872
rect 28491 112832 29828 112860
rect 28491 112829 28503 112832
rect 28445 112823 28503 112829
rect 29822 112820 29828 112832
rect 29880 112820 29886 112872
rect 31386 112820 31392 112872
rect 31444 112860 31450 112872
rect 31573 112863 31631 112869
rect 31573 112860 31585 112863
rect 31444 112832 31585 112860
rect 31444 112820 31450 112832
rect 31573 112829 31585 112832
rect 31619 112829 31631 112863
rect 31573 112823 31631 112829
rect 33318 112820 33324 112872
rect 33376 112860 33382 112872
rect 33505 112863 33563 112869
rect 33505 112860 33517 112863
rect 33376 112832 33517 112860
rect 33376 112820 33382 112832
rect 33505 112829 33517 112832
rect 33551 112829 33563 112863
rect 33505 112823 33563 112829
rect 33594 112820 33600 112872
rect 33652 112860 33658 112872
rect 37936 112869 37964 112900
rect 34149 112863 34207 112869
rect 34149 112860 34161 112863
rect 33652 112832 34161 112860
rect 33652 112820 33658 112832
rect 34149 112829 34161 112832
rect 34195 112829 34207 112863
rect 37185 112863 37243 112869
rect 37185 112860 37197 112863
rect 34149 112823 34207 112829
rect 34486 112832 37197 112860
rect 31938 112752 31944 112804
rect 31996 112792 32002 112804
rect 34486 112792 34514 112832
rect 37185 112829 37197 112832
rect 37231 112829 37243 112863
rect 37185 112823 37243 112829
rect 37921 112863 37979 112869
rect 37921 112829 37933 112863
rect 37967 112829 37979 112863
rect 37921 112823 37979 112829
rect 31996 112764 34514 112792
rect 31996 112752 32002 112764
rect 36354 112752 36360 112804
rect 36412 112792 36418 112804
rect 36449 112795 36507 112801
rect 36449 112792 36461 112795
rect 36412 112764 36461 112792
rect 36412 112752 36418 112764
rect 36449 112761 36461 112764
rect 36495 112761 36507 112795
rect 37366 112792 37372 112804
rect 37327 112764 37372 112792
rect 36449 112755 36507 112761
rect 37366 112752 37372 112764
rect 37424 112752 37430 112804
rect 38102 112792 38108 112804
rect 38063 112764 38108 112792
rect 38102 112752 38108 112764
rect 38160 112752 38166 112804
rect 2133 112727 2191 112733
rect 2133 112693 2145 112727
rect 2179 112724 2191 112727
rect 16022 112724 16028 112736
rect 2179 112696 16028 112724
rect 2179 112693 2191 112696
rect 2133 112687 2191 112693
rect 16022 112684 16028 112696
rect 16080 112684 16086 112736
rect 26234 112684 26240 112736
rect 26292 112724 26298 112736
rect 28629 112727 28687 112733
rect 28629 112724 28641 112727
rect 26292 112696 28641 112724
rect 26292 112684 26298 112696
rect 28629 112693 28641 112696
rect 28675 112693 28687 112727
rect 28629 112687 28687 112693
rect 33134 112684 33140 112736
rect 33192 112724 33198 112736
rect 34238 112724 34244 112736
rect 33192 112696 34244 112724
rect 33192 112684 33198 112696
rect 34238 112684 34244 112696
rect 34296 112684 34302 112736
rect 1104 112634 38824 112656
rect 1104 112582 19606 112634
rect 19658 112582 19670 112634
rect 19722 112582 19734 112634
rect 19786 112582 19798 112634
rect 19850 112582 38824 112634
rect 1104 112560 38824 112582
rect 35802 112480 35808 112532
rect 35860 112520 35866 112532
rect 36541 112523 36599 112529
rect 36541 112520 36553 112523
rect 35860 112492 36553 112520
rect 35860 112480 35866 112492
rect 36541 112489 36553 112492
rect 36587 112489 36599 112523
rect 36541 112483 36599 112489
rect 20714 112412 20720 112464
rect 20772 112452 20778 112464
rect 20772 112424 22094 112452
rect 20772 112412 20778 112424
rect 1857 112387 1915 112393
rect 1857 112353 1869 112387
rect 1903 112384 1915 112387
rect 12710 112384 12716 112396
rect 1903 112356 12716 112384
rect 1903 112353 1915 112356
rect 1857 112347 1915 112353
rect 12710 112344 12716 112356
rect 12768 112344 12774 112396
rect 22066 112248 22094 112424
rect 23566 112412 23572 112464
rect 23624 112452 23630 112464
rect 35986 112452 35992 112464
rect 23624 112424 35992 112452
rect 23624 112412 23630 112424
rect 35986 112412 35992 112424
rect 36044 112412 36050 112464
rect 37369 112455 37427 112461
rect 37369 112421 37381 112455
rect 37415 112452 37427 112455
rect 39850 112452 39856 112464
rect 37415 112424 39856 112452
rect 37415 112421 37427 112424
rect 37369 112415 37427 112421
rect 39850 112412 39856 112424
rect 39908 112412 39914 112464
rect 36449 112387 36507 112393
rect 36449 112353 36461 112387
rect 36495 112353 36507 112387
rect 36449 112347 36507 112353
rect 34422 112248 34428 112260
rect 22066 112220 34428 112248
rect 34422 112208 34428 112220
rect 34480 112208 34486 112260
rect 1946 112180 1952 112192
rect 1907 112152 1952 112180
rect 1946 112140 1952 112152
rect 2004 112140 2010 112192
rect 23290 112140 23296 112192
rect 23348 112180 23354 112192
rect 36464 112180 36492 112347
rect 36814 112344 36820 112396
rect 36872 112384 36878 112396
rect 37185 112387 37243 112393
rect 37185 112384 37197 112387
rect 36872 112356 37197 112384
rect 36872 112344 36878 112356
rect 37185 112353 37197 112356
rect 37231 112353 37243 112387
rect 37185 112347 37243 112353
rect 23348 112152 36492 112180
rect 23348 112140 23354 112152
rect 1104 112090 38824 112112
rect 1104 112038 4246 112090
rect 4298 112038 4310 112090
rect 4362 112038 4374 112090
rect 4426 112038 4438 112090
rect 4490 112038 34966 112090
rect 35018 112038 35030 112090
rect 35082 112038 35094 112090
rect 35146 112038 35158 112090
rect 35210 112038 38824 112090
rect 1104 112016 38824 112038
rect 35526 111800 35532 111852
rect 35584 111840 35590 111852
rect 35802 111840 35808 111852
rect 35584 111812 35808 111840
rect 35584 111800 35590 111812
rect 35802 111800 35808 111812
rect 35860 111800 35866 111852
rect 37642 111772 37648 111784
rect 37603 111744 37648 111772
rect 37642 111732 37648 111744
rect 37700 111732 37706 111784
rect 35526 111664 35532 111716
rect 35584 111704 35590 111716
rect 37921 111707 37979 111713
rect 37921 111704 37933 111707
rect 35584 111676 37933 111704
rect 35584 111664 35590 111676
rect 37921 111673 37933 111676
rect 37967 111673 37979 111707
rect 37921 111667 37979 111673
rect 1104 111546 38824 111568
rect 1104 111494 19606 111546
rect 19658 111494 19670 111546
rect 19722 111494 19734 111546
rect 19786 111494 19798 111546
rect 19850 111494 38824 111546
rect 1104 111472 38824 111494
rect 31757 111435 31815 111441
rect 31757 111401 31769 111435
rect 31803 111432 31815 111435
rect 33778 111432 33784 111444
rect 31803 111404 33784 111432
rect 31803 111401 31815 111404
rect 31757 111395 31815 111401
rect 33778 111392 33784 111404
rect 33836 111392 33842 111444
rect 36538 111432 36544 111444
rect 36499 111404 36544 111432
rect 36538 111392 36544 111404
rect 36596 111392 36602 111444
rect 25314 111324 25320 111376
rect 25372 111364 25378 111376
rect 34514 111364 34520 111376
rect 25372 111336 34520 111364
rect 25372 111324 25378 111336
rect 34514 111324 34520 111336
rect 34572 111324 34578 111376
rect 1394 111296 1400 111308
rect 1355 111268 1400 111296
rect 1394 111256 1400 111268
rect 1452 111256 1458 111308
rect 31478 111256 31484 111308
rect 31536 111296 31542 111308
rect 31573 111299 31631 111305
rect 31573 111296 31585 111299
rect 31536 111268 31585 111296
rect 31536 111256 31542 111268
rect 31573 111265 31585 111268
rect 31619 111265 31631 111299
rect 36446 111296 36452 111308
rect 36407 111268 36452 111296
rect 31573 111259 31631 111265
rect 36446 111256 36452 111268
rect 36504 111256 36510 111308
rect 37185 111299 37243 111305
rect 37185 111265 37197 111299
rect 37231 111265 37243 111299
rect 37185 111259 37243 111265
rect 1673 111231 1731 111237
rect 1673 111197 1685 111231
rect 1719 111228 1731 111231
rect 7650 111228 7656 111240
rect 1719 111200 7656 111228
rect 1719 111197 1731 111200
rect 1673 111191 1731 111197
rect 7650 111188 7656 111200
rect 7708 111188 7714 111240
rect 31110 111188 31116 111240
rect 31168 111228 31174 111240
rect 37200 111228 37228 111259
rect 31168 111200 37228 111228
rect 31168 111188 31174 111200
rect 26786 111120 26792 111172
rect 26844 111160 26850 111172
rect 37366 111160 37372 111172
rect 26844 111132 36032 111160
rect 37327 111132 37372 111160
rect 26844 111120 26850 111132
rect 34606 111052 34612 111104
rect 34664 111092 34670 111104
rect 35894 111092 35900 111104
rect 34664 111064 35900 111092
rect 34664 111052 34670 111064
rect 35894 111052 35900 111064
rect 35952 111052 35958 111104
rect 36004 111092 36032 111132
rect 37366 111120 37372 111132
rect 37424 111120 37430 111172
rect 37458 111092 37464 111104
rect 36004 111064 37464 111092
rect 37458 111052 37464 111064
rect 37516 111052 37522 111104
rect 1104 111002 38824 111024
rect 1104 110950 4246 111002
rect 4298 110950 4310 111002
rect 4362 110950 4374 111002
rect 4426 110950 4438 111002
rect 4490 110950 34966 111002
rect 35018 110950 35030 111002
rect 35082 110950 35094 111002
rect 35146 110950 35158 111002
rect 35210 110950 38824 111002
rect 1104 110928 38824 110950
rect 28258 110848 28264 110900
rect 28316 110888 28322 110900
rect 36446 110888 36452 110900
rect 28316 110860 36452 110888
rect 28316 110848 28322 110860
rect 36446 110848 36452 110860
rect 36504 110848 36510 110900
rect 36262 110712 36268 110764
rect 36320 110752 36326 110764
rect 36446 110752 36452 110764
rect 36320 110724 36452 110752
rect 36320 110712 36326 110724
rect 36446 110712 36452 110724
rect 36504 110712 36510 110764
rect 37458 110684 37464 110696
rect 37419 110656 37464 110684
rect 37458 110644 37464 110656
rect 37516 110644 37522 110696
rect 1857 110619 1915 110625
rect 1857 110585 1869 110619
rect 1903 110616 1915 110619
rect 2222 110616 2228 110628
rect 1903 110588 2228 110616
rect 1903 110585 1915 110588
rect 1857 110579 1915 110585
rect 2222 110576 2228 110588
rect 2280 110576 2286 110628
rect 37826 110616 37832 110628
rect 37787 110588 37832 110616
rect 37826 110576 37832 110588
rect 37884 110576 37890 110628
rect 1946 110548 1952 110560
rect 1907 110520 1952 110548
rect 1946 110508 1952 110520
rect 2004 110508 2010 110560
rect 1104 110458 38824 110480
rect 1104 110406 19606 110458
rect 19658 110406 19670 110458
rect 19722 110406 19734 110458
rect 19786 110406 19798 110458
rect 19850 110406 38824 110458
rect 1104 110384 38824 110406
rect 37182 110208 37188 110220
rect 37143 110180 37188 110208
rect 37182 110168 37188 110180
rect 37240 110168 37246 110220
rect 22554 110032 22560 110084
rect 22612 110072 22618 110084
rect 32766 110072 32772 110084
rect 22612 110044 32772 110072
rect 22612 110032 22618 110044
rect 32766 110032 32772 110044
rect 32824 110032 32830 110084
rect 37369 110075 37427 110081
rect 37369 110041 37381 110075
rect 37415 110072 37427 110075
rect 38194 110072 38200 110084
rect 37415 110044 38200 110072
rect 37415 110041 37427 110044
rect 37369 110035 37427 110041
rect 38194 110032 38200 110044
rect 38252 110032 38258 110084
rect 26694 109964 26700 110016
rect 26752 110004 26758 110016
rect 36906 110004 36912 110016
rect 26752 109976 36912 110004
rect 26752 109964 26758 109976
rect 36906 109964 36912 109976
rect 36964 109964 36970 110016
rect 1104 109914 38824 109936
rect 1104 109862 4246 109914
rect 4298 109862 4310 109914
rect 4362 109862 4374 109914
rect 4426 109862 4438 109914
rect 4490 109862 34966 109914
rect 35018 109862 35030 109914
rect 35082 109862 35094 109914
rect 35146 109862 35158 109914
rect 35210 109862 38824 109914
rect 1104 109840 38824 109862
rect 24670 109760 24676 109812
rect 24728 109800 24734 109812
rect 37826 109800 37832 109812
rect 24728 109772 37832 109800
rect 24728 109760 24734 109772
rect 37826 109760 37832 109772
rect 37884 109760 37890 109812
rect 5258 109692 5264 109744
rect 5316 109732 5322 109744
rect 26234 109732 26240 109744
rect 5316 109704 26240 109732
rect 5316 109692 5322 109704
rect 26234 109692 26240 109704
rect 26292 109692 26298 109744
rect 27614 109692 27620 109744
rect 27672 109732 27678 109744
rect 36170 109732 36176 109744
rect 27672 109704 36176 109732
rect 27672 109692 27678 109704
rect 36170 109692 36176 109704
rect 36228 109692 36234 109744
rect 2038 109596 2044 109608
rect 1999 109568 2044 109596
rect 2038 109556 2044 109568
rect 2096 109556 2102 109608
rect 37182 109596 37188 109608
rect 37143 109568 37188 109596
rect 37182 109556 37188 109568
rect 37240 109556 37246 109608
rect 1857 109531 1915 109537
rect 1857 109497 1869 109531
rect 1903 109528 1915 109531
rect 11054 109528 11060 109540
rect 1903 109500 11060 109528
rect 1903 109497 1915 109500
rect 1857 109491 1915 109497
rect 11054 109488 11060 109500
rect 11112 109488 11118 109540
rect 37918 109528 37924 109540
rect 37879 109500 37924 109528
rect 37918 109488 37924 109500
rect 37976 109488 37982 109540
rect 38105 109531 38163 109537
rect 38105 109497 38117 109531
rect 38151 109528 38163 109531
rect 38654 109528 38660 109540
rect 38151 109500 38660 109528
rect 38151 109497 38163 109500
rect 38105 109491 38163 109497
rect 38654 109488 38660 109500
rect 38712 109488 38718 109540
rect 37277 109463 37335 109469
rect 37277 109429 37289 109463
rect 37323 109460 37335 109463
rect 38378 109460 38384 109472
rect 37323 109432 38384 109460
rect 37323 109429 37335 109432
rect 37277 109423 37335 109429
rect 38378 109420 38384 109432
rect 38436 109420 38442 109472
rect 1104 109370 38824 109392
rect 1104 109318 19606 109370
rect 19658 109318 19670 109370
rect 19722 109318 19734 109370
rect 19786 109318 19798 109370
rect 19850 109318 38824 109370
rect 1104 109296 38824 109318
rect 8662 109256 8668 109268
rect 8623 109228 8668 109256
rect 8662 109216 8668 109228
rect 8720 109216 8726 109268
rect 8481 109123 8539 109129
rect 8481 109089 8493 109123
rect 8527 109120 8539 109123
rect 13078 109120 13084 109132
rect 8527 109092 13084 109120
rect 8527 109089 8539 109092
rect 8481 109083 8539 109089
rect 13078 109080 13084 109092
rect 13136 109080 13142 109132
rect 37182 109120 37188 109132
rect 37143 109092 37188 109120
rect 37182 109080 37188 109092
rect 37240 109080 37246 109132
rect 2498 109012 2504 109064
rect 2556 109052 2562 109064
rect 3418 109052 3424 109064
rect 2556 109024 3424 109052
rect 2556 109012 2562 109024
rect 3418 109012 3424 109024
rect 3476 109012 3482 109064
rect 32674 109012 32680 109064
rect 32732 109052 32738 109064
rect 37369 109055 37427 109061
rect 37369 109052 37381 109055
rect 32732 109024 37381 109052
rect 32732 109012 32738 109024
rect 37369 109021 37381 109024
rect 37415 109021 37427 109055
rect 37369 109015 37427 109021
rect 1104 108826 38824 108848
rect 1104 108774 4246 108826
rect 4298 108774 4310 108826
rect 4362 108774 4374 108826
rect 4426 108774 4438 108826
rect 4490 108774 34966 108826
rect 35018 108774 35030 108826
rect 35082 108774 35094 108826
rect 35146 108774 35158 108826
rect 35210 108774 38824 108826
rect 1104 108752 38824 108774
rect 1946 108712 1952 108724
rect 1907 108684 1952 108712
rect 1946 108672 1952 108684
rect 2004 108672 2010 108724
rect 32766 108468 32772 108520
rect 32824 108508 32830 108520
rect 38105 108511 38163 108517
rect 38105 108508 38117 108511
rect 32824 108480 38117 108508
rect 32824 108468 32830 108480
rect 38105 108477 38117 108480
rect 38151 108477 38163 108511
rect 38105 108471 38163 108477
rect 1857 108443 1915 108449
rect 1857 108409 1869 108443
rect 1903 108440 1915 108443
rect 7558 108440 7564 108452
rect 1903 108412 7564 108440
rect 1903 108409 1915 108412
rect 1857 108403 1915 108409
rect 7558 108400 7564 108412
rect 7616 108400 7622 108452
rect 21542 108400 21548 108452
rect 21600 108440 21606 108452
rect 33226 108440 33232 108452
rect 21600 108412 33232 108440
rect 21600 108400 21606 108412
rect 33226 108400 33232 108412
rect 33284 108400 33290 108452
rect 37918 108440 37924 108452
rect 37879 108412 37924 108440
rect 37918 108400 37924 108412
rect 37976 108400 37982 108452
rect 23106 108332 23112 108384
rect 23164 108372 23170 108384
rect 31938 108372 31944 108384
rect 23164 108344 31944 108372
rect 23164 108332 23170 108344
rect 31938 108332 31944 108344
rect 31996 108332 32002 108384
rect 1104 108282 38824 108304
rect 1104 108230 19606 108282
rect 19658 108230 19670 108282
rect 19722 108230 19734 108282
rect 19786 108230 19798 108282
rect 19850 108230 38824 108282
rect 1104 108208 38824 108230
rect 1857 108035 1915 108041
rect 1857 108001 1869 108035
rect 1903 108032 1915 108035
rect 13446 108032 13452 108044
rect 1903 108004 13452 108032
rect 1903 108001 1915 108004
rect 1857 107995 1915 108001
rect 13446 107992 13452 108004
rect 13504 107992 13510 108044
rect 37182 108032 37188 108044
rect 37143 108004 37188 108032
rect 37182 107992 37188 108004
rect 37240 107992 37246 108044
rect 2038 107896 2044 107908
rect 1999 107868 2044 107896
rect 2038 107856 2044 107868
rect 2096 107856 2102 107908
rect 33226 107788 33232 107840
rect 33284 107828 33290 107840
rect 37277 107831 37335 107837
rect 37277 107828 37289 107831
rect 33284 107800 37289 107828
rect 33284 107788 33290 107800
rect 37277 107797 37289 107800
rect 37323 107797 37335 107831
rect 37277 107791 37335 107797
rect 1104 107738 38824 107760
rect 1104 107686 4246 107738
rect 4298 107686 4310 107738
rect 4362 107686 4374 107738
rect 4426 107686 4438 107738
rect 4490 107686 34966 107738
rect 35018 107686 35030 107738
rect 35082 107686 35094 107738
rect 35146 107686 35158 107738
rect 35210 107686 38824 107738
rect 1104 107664 38824 107686
rect 32950 107584 32956 107636
rect 33008 107624 33014 107636
rect 37366 107624 37372 107636
rect 33008 107596 37372 107624
rect 33008 107584 33014 107596
rect 37366 107584 37372 107596
rect 37424 107584 37430 107636
rect 37182 107420 37188 107432
rect 37143 107392 37188 107420
rect 37182 107380 37188 107392
rect 37240 107380 37246 107432
rect 37369 107355 37427 107361
rect 37369 107321 37381 107355
rect 37415 107352 37427 107355
rect 37550 107352 37556 107364
rect 37415 107324 37556 107352
rect 37415 107321 37427 107324
rect 37369 107315 37427 107321
rect 37550 107312 37556 107324
rect 37608 107312 37614 107364
rect 37918 107352 37924 107364
rect 37879 107324 37924 107352
rect 37918 107312 37924 107324
rect 37976 107312 37982 107364
rect 36906 107244 36912 107296
rect 36964 107284 36970 107296
rect 38013 107287 38071 107293
rect 38013 107284 38025 107287
rect 36964 107256 38025 107284
rect 36964 107244 36970 107256
rect 38013 107253 38025 107256
rect 38059 107253 38071 107287
rect 38013 107247 38071 107253
rect 1104 107194 38824 107216
rect 1104 107142 19606 107194
rect 19658 107142 19670 107194
rect 19722 107142 19734 107194
rect 19786 107142 19798 107194
rect 19850 107142 38824 107194
rect 1104 107120 38824 107142
rect 1946 107080 1952 107092
rect 1907 107052 1952 107080
rect 1946 107040 1952 107052
rect 2004 107040 2010 107092
rect 24026 106972 24032 107024
rect 24084 107012 24090 107024
rect 37826 107012 37832 107024
rect 24084 106984 37832 107012
rect 24084 106972 24090 106984
rect 37826 106972 37832 106984
rect 37884 106972 37890 107024
rect 1857 106947 1915 106953
rect 1857 106913 1869 106947
rect 1903 106944 1915 106947
rect 7742 106944 7748 106956
rect 1903 106916 7748 106944
rect 1903 106913 1915 106916
rect 1857 106907 1915 106913
rect 7742 106904 7748 106916
rect 7800 106904 7806 106956
rect 22462 106904 22468 106956
rect 22520 106944 22526 106956
rect 32398 106944 32404 106956
rect 22520 106916 32404 106944
rect 22520 106904 22526 106916
rect 32398 106904 32404 106916
rect 32456 106904 32462 106956
rect 37182 106944 37188 106956
rect 37143 106916 37188 106944
rect 37182 106904 37188 106916
rect 37240 106904 37246 106956
rect 37369 106811 37427 106817
rect 37369 106777 37381 106811
rect 37415 106808 37427 106811
rect 38470 106808 38476 106820
rect 37415 106780 38476 106808
rect 37415 106777 37427 106780
rect 37369 106771 37427 106777
rect 38470 106768 38476 106780
rect 38528 106768 38534 106820
rect 1104 106650 38824 106672
rect 1104 106598 4246 106650
rect 4298 106598 4310 106650
rect 4362 106598 4374 106650
rect 4426 106598 4438 106650
rect 4490 106598 34966 106650
rect 35018 106598 35030 106650
rect 35082 106598 35094 106650
rect 35146 106598 35158 106650
rect 35210 106598 38824 106650
rect 1104 106576 38824 106598
rect 1673 106403 1731 106409
rect 1673 106369 1685 106403
rect 1719 106400 1731 106403
rect 29638 106400 29644 106412
rect 1719 106372 29644 106400
rect 1719 106369 1731 106372
rect 1673 106363 1731 106369
rect 1762 106332 1768 106344
rect 1723 106304 1768 106332
rect 1762 106292 1768 106304
rect 1820 106292 1826 106344
rect 1964 106341 1992 106372
rect 29638 106360 29644 106372
rect 29696 106360 29702 106412
rect 36538 106360 36544 106412
rect 36596 106400 36602 106412
rect 37553 106403 37611 106409
rect 37553 106400 37565 106403
rect 36596 106372 37565 106400
rect 36596 106360 36602 106372
rect 37553 106369 37565 106372
rect 37599 106369 37611 106403
rect 37553 106363 37611 106369
rect 1949 106335 2007 106341
rect 1949 106301 1961 106335
rect 1995 106301 2007 106335
rect 1949 106295 2007 106301
rect 32858 106292 32864 106344
rect 32916 106332 32922 106344
rect 33226 106332 33232 106344
rect 32916 106304 33232 106332
rect 32916 106292 32922 106304
rect 33226 106292 33232 106304
rect 33284 106292 33290 106344
rect 37274 106332 37280 106344
rect 37235 106304 37280 106332
rect 37274 106292 37280 106304
rect 37332 106292 37338 106344
rect 1104 106106 38824 106128
rect 1104 106054 19606 106106
rect 19658 106054 19670 106106
rect 19722 106054 19734 106106
rect 19786 106054 19798 106106
rect 19850 106054 38824 106106
rect 1104 106032 38824 106054
rect 37182 105856 37188 105868
rect 37143 105828 37188 105856
rect 37182 105816 37188 105828
rect 37240 105816 37246 105868
rect 25958 105680 25964 105732
rect 26016 105720 26022 105732
rect 35802 105720 35808 105732
rect 26016 105692 35808 105720
rect 26016 105680 26022 105692
rect 35802 105680 35808 105692
rect 35860 105680 35866 105732
rect 33318 105612 33324 105664
rect 33376 105652 33382 105664
rect 37277 105655 37335 105661
rect 37277 105652 37289 105655
rect 33376 105624 37289 105652
rect 33376 105612 33382 105624
rect 37277 105621 37289 105624
rect 37323 105621 37335 105655
rect 37277 105615 37335 105621
rect 1104 105562 38824 105584
rect 1104 105510 4246 105562
rect 4298 105510 4310 105562
rect 4362 105510 4374 105562
rect 4426 105510 4438 105562
rect 4490 105510 34966 105562
rect 35018 105510 35030 105562
rect 35082 105510 35094 105562
rect 35146 105510 35158 105562
rect 35210 105510 38824 105562
rect 1104 105488 38824 105510
rect 26329 105451 26387 105457
rect 26329 105417 26341 105451
rect 26375 105448 26387 105451
rect 27614 105448 27620 105460
rect 26375 105420 27620 105448
rect 26375 105417 26387 105420
rect 26329 105411 26387 105417
rect 27614 105408 27620 105420
rect 27672 105408 27678 105460
rect 32217 105451 32275 105457
rect 32217 105417 32229 105451
rect 32263 105448 32275 105451
rect 36078 105448 36084 105460
rect 32263 105420 36084 105448
rect 32263 105417 32275 105420
rect 32217 105411 32275 105417
rect 36078 105408 36084 105420
rect 36136 105408 36142 105460
rect 1394 105244 1400 105256
rect 1355 105216 1400 105244
rect 1394 105204 1400 105216
rect 1452 105204 1458 105256
rect 24854 105204 24860 105256
rect 24912 105244 24918 105256
rect 25225 105247 25283 105253
rect 25225 105244 25237 105247
rect 24912 105216 25237 105244
rect 24912 105204 24918 105216
rect 25225 105213 25237 105216
rect 25271 105213 25283 105247
rect 25225 105207 25283 105213
rect 25685 105247 25743 105253
rect 25685 105213 25697 105247
rect 25731 105213 25743 105247
rect 26050 105244 26056 105256
rect 26011 105216 26056 105244
rect 25685 105207 25743 105213
rect 20622 105136 20628 105188
rect 20680 105176 20686 105188
rect 25700 105176 25728 105207
rect 26050 105204 26056 105216
rect 26108 105204 26114 105256
rect 32030 105244 32036 105256
rect 31991 105216 32036 105244
rect 32030 105204 32036 105216
rect 32088 105204 32094 105256
rect 37182 105244 37188 105256
rect 37143 105216 37188 105244
rect 37182 105204 37188 105216
rect 37240 105204 37246 105256
rect 37918 105176 37924 105188
rect 20680 105148 25728 105176
rect 37879 105148 37924 105176
rect 20680 105136 20686 105148
rect 37918 105136 37924 105148
rect 37976 105136 37982 105188
rect 1581 105111 1639 105117
rect 1581 105077 1593 105111
rect 1627 105108 1639 105111
rect 8938 105108 8944 105120
rect 1627 105080 8944 105108
rect 1627 105077 1639 105080
rect 1581 105071 1639 105077
rect 8938 105068 8944 105080
rect 8996 105068 9002 105120
rect 34146 105068 34152 105120
rect 34204 105108 34210 105120
rect 37277 105111 37335 105117
rect 37277 105108 37289 105111
rect 34204 105080 37289 105108
rect 34204 105068 34210 105080
rect 37277 105077 37289 105080
rect 37323 105077 37335 105111
rect 38010 105108 38016 105120
rect 37971 105080 38016 105108
rect 37277 105071 37335 105077
rect 38010 105068 38016 105080
rect 38068 105068 38074 105120
rect 1104 105018 38824 105040
rect 1104 104966 19606 105018
rect 19658 104966 19670 105018
rect 19722 104966 19734 105018
rect 19786 104966 19798 105018
rect 19850 104966 38824 105018
rect 1104 104944 38824 104966
rect 25958 104904 25964 104916
rect 25919 104876 25964 104904
rect 25958 104864 25964 104876
rect 26016 104864 26022 104916
rect 20438 104796 20444 104848
rect 20496 104836 20502 104848
rect 26050 104836 26056 104848
rect 20496 104808 26056 104836
rect 20496 104796 20502 104808
rect 1854 104768 1860 104780
rect 1815 104740 1860 104768
rect 1854 104728 1860 104740
rect 1912 104728 1918 104780
rect 24854 104768 24860 104780
rect 24815 104740 24860 104768
rect 24854 104728 24860 104740
rect 24912 104728 24918 104780
rect 25700 104777 25728 104808
rect 26050 104796 26056 104808
rect 26108 104796 26114 104848
rect 25317 104771 25375 104777
rect 25317 104737 25329 104771
rect 25363 104737 25375 104771
rect 25317 104731 25375 104737
rect 25685 104771 25743 104777
rect 25685 104737 25697 104771
rect 25731 104737 25743 104771
rect 37182 104768 37188 104780
rect 37143 104740 37188 104768
rect 25685 104731 25743 104737
rect 21266 104660 21272 104712
rect 21324 104700 21330 104712
rect 25332 104700 25360 104731
rect 37182 104728 37188 104740
rect 37240 104728 37246 104780
rect 21324 104672 25360 104700
rect 21324 104660 21330 104672
rect 1949 104567 2007 104573
rect 1949 104533 1961 104567
rect 1995 104564 2007 104567
rect 10318 104564 10324 104576
rect 1995 104536 10324 104564
rect 1995 104533 2007 104536
rect 1949 104527 2007 104533
rect 10318 104524 10324 104536
rect 10376 104524 10382 104576
rect 36998 104524 37004 104576
rect 37056 104564 37062 104576
rect 37277 104567 37335 104573
rect 37277 104564 37289 104567
rect 37056 104536 37289 104564
rect 37056 104524 37062 104536
rect 37277 104533 37289 104536
rect 37323 104533 37335 104567
rect 37277 104527 37335 104533
rect 1104 104474 38824 104496
rect 1104 104422 4246 104474
rect 4298 104422 4310 104474
rect 4362 104422 4374 104474
rect 4426 104422 4438 104474
rect 4490 104422 34966 104474
rect 35018 104422 35030 104474
rect 35082 104422 35094 104474
rect 35146 104422 35158 104474
rect 35210 104422 38824 104474
rect 1104 104400 38824 104422
rect 29549 104363 29607 104369
rect 29549 104329 29561 104363
rect 29595 104360 29607 104363
rect 35342 104360 35348 104372
rect 29595 104332 35348 104360
rect 29595 104329 29607 104332
rect 29549 104323 29607 104329
rect 35342 104320 35348 104332
rect 35400 104320 35406 104372
rect 24946 104184 24952 104236
rect 25004 104224 25010 104236
rect 31386 104224 31392 104236
rect 25004 104196 31392 104224
rect 25004 104184 25010 104196
rect 31386 104184 31392 104196
rect 31444 104184 31450 104236
rect 26878 104116 26884 104168
rect 26936 104156 26942 104168
rect 29365 104159 29423 104165
rect 29365 104156 29377 104159
rect 26936 104128 29377 104156
rect 26936 104116 26942 104128
rect 29365 104125 29377 104128
rect 29411 104125 29423 104159
rect 29365 104119 29423 104125
rect 34238 104116 34244 104168
rect 34296 104156 34302 104168
rect 38010 104156 38016 104168
rect 34296 104128 38016 104156
rect 34296 104116 34302 104128
rect 38010 104116 38016 104128
rect 38068 104116 38074 104168
rect 37182 104088 37188 104100
rect 37143 104060 37188 104088
rect 37182 104048 37188 104060
rect 37240 104048 37246 104100
rect 37366 104088 37372 104100
rect 37327 104060 37372 104088
rect 37366 104048 37372 104060
rect 37424 104048 37430 104100
rect 37918 104088 37924 104100
rect 37879 104060 37924 104088
rect 37918 104048 37924 104060
rect 37976 104048 37982 104100
rect 38010 104020 38016 104032
rect 37971 103992 38016 104020
rect 38010 103980 38016 103992
rect 38068 103980 38074 104032
rect 1104 103930 38824 103952
rect 1104 103878 19606 103930
rect 19658 103878 19670 103930
rect 19722 103878 19734 103930
rect 19786 103878 19798 103930
rect 19850 103878 38824 103930
rect 1104 103856 38824 103878
rect 11054 103776 11060 103828
rect 11112 103816 11118 103828
rect 12529 103819 12587 103825
rect 12529 103816 12541 103819
rect 11112 103788 12541 103816
rect 11112 103776 11118 103788
rect 12529 103785 12541 103788
rect 12575 103785 12587 103819
rect 21266 103816 21272 103828
rect 12529 103779 12587 103785
rect 13096 103788 21272 103816
rect 1854 103748 1860 103760
rect 1815 103720 1860 103748
rect 1854 103708 1860 103720
rect 1912 103708 1918 103760
rect 12526 103680 12532 103692
rect 12487 103652 12532 103680
rect 12526 103640 12532 103652
rect 12584 103640 12590 103692
rect 12618 103640 12624 103692
rect 12676 103680 12682 103692
rect 13096 103689 13124 103788
rect 21266 103776 21272 103788
rect 21324 103776 21330 103828
rect 21634 103816 21640 103828
rect 21595 103788 21640 103816
rect 21634 103776 21640 103788
rect 21692 103776 21698 103828
rect 18322 103748 18328 103760
rect 13280 103720 18328 103748
rect 13280 103689 13308 103720
rect 18322 103708 18328 103720
rect 18380 103748 18386 103760
rect 20438 103748 20444 103760
rect 18380 103720 20444 103748
rect 18380 103708 18386 103720
rect 20438 103708 20444 103720
rect 20496 103708 20502 103760
rect 20530 103708 20536 103760
rect 20588 103748 20594 103760
rect 21478 103751 21536 103757
rect 21478 103748 21490 103751
rect 20588 103720 21490 103748
rect 20588 103708 20594 103720
rect 21478 103717 21490 103720
rect 21524 103748 21536 103751
rect 24854 103748 24860 103760
rect 21524 103720 24860 103748
rect 21524 103717 21536 103720
rect 21478 103711 21536 103717
rect 24854 103708 24860 103720
rect 24912 103708 24918 103760
rect 25133 103751 25191 103757
rect 25133 103717 25145 103751
rect 25179 103748 25191 103751
rect 26786 103748 26792 103760
rect 25179 103720 26792 103748
rect 25179 103717 25191 103720
rect 25133 103711 25191 103717
rect 26786 103708 26792 103720
rect 26844 103708 26850 103760
rect 13081 103683 13139 103689
rect 13081 103680 13093 103683
rect 12676 103652 13093 103680
rect 12676 103640 12682 103652
rect 13081 103649 13093 103652
rect 13127 103649 13139 103683
rect 13081 103643 13139 103649
rect 13265 103683 13323 103689
rect 13265 103649 13277 103683
rect 13311 103649 13323 103683
rect 13265 103643 13323 103649
rect 14458 103640 14464 103692
rect 14516 103680 14522 103692
rect 24949 103683 25007 103689
rect 24949 103680 24961 103683
rect 14516 103652 24961 103680
rect 14516 103640 14522 103652
rect 24949 103649 24961 103652
rect 24995 103649 25007 103683
rect 37182 103680 37188 103692
rect 37143 103652 37188 103680
rect 24949 103643 25007 103649
rect 37182 103640 37188 103652
rect 37240 103640 37246 103692
rect 18046 103572 18052 103624
rect 18104 103612 18110 103624
rect 20993 103615 21051 103621
rect 20993 103612 21005 103615
rect 18104 103584 21005 103612
rect 18104 103572 18110 103584
rect 20993 103581 21005 103584
rect 21039 103581 21051 103615
rect 20993 103575 21051 103581
rect 21361 103615 21419 103621
rect 21361 103581 21373 103615
rect 21407 103581 21419 103615
rect 21361 103575 21419 103581
rect 2041 103547 2099 103553
rect 2041 103513 2053 103547
rect 2087 103544 2099 103547
rect 9030 103544 9036 103556
rect 2087 103516 9036 103544
rect 2087 103513 2099 103516
rect 2041 103507 2099 103513
rect 9030 103504 9036 103516
rect 9088 103504 9094 103556
rect 21376 103544 21404 103575
rect 31202 103572 31208 103624
rect 31260 103612 31266 103624
rect 37369 103615 37427 103621
rect 37369 103612 37381 103615
rect 31260 103584 37381 103612
rect 31260 103572 31266 103584
rect 37369 103581 37381 103584
rect 37415 103581 37427 103615
rect 37369 103575 37427 103581
rect 16592 103516 21404 103544
rect 16592 103488 16620 103516
rect 32306 103504 32312 103556
rect 32364 103544 32370 103556
rect 36906 103544 36912 103556
rect 32364 103516 36912 103544
rect 32364 103504 32370 103516
rect 36906 103504 36912 103516
rect 36964 103504 36970 103556
rect 13538 103436 13544 103488
rect 13596 103476 13602 103488
rect 16574 103476 16580 103488
rect 13596 103448 16580 103476
rect 13596 103436 13602 103448
rect 16574 103436 16580 103448
rect 16632 103436 16638 103488
rect 18322 103436 18328 103488
rect 18380 103476 18386 103488
rect 19334 103476 19340 103488
rect 18380 103448 19340 103476
rect 18380 103436 18386 103448
rect 19334 103436 19340 103448
rect 19392 103436 19398 103488
rect 1104 103386 38824 103408
rect 1104 103334 4246 103386
rect 4298 103334 4310 103386
rect 4362 103334 4374 103386
rect 4426 103334 4438 103386
rect 4490 103334 34966 103386
rect 35018 103334 35030 103386
rect 35082 103334 35094 103386
rect 35146 103334 35158 103386
rect 35210 103334 38824 103386
rect 1104 103312 38824 103334
rect 3510 103232 3516 103284
rect 3568 103272 3574 103284
rect 6365 103275 6423 103281
rect 6365 103272 6377 103275
rect 3568 103244 6377 103272
rect 3568 103232 3574 103244
rect 6365 103241 6377 103244
rect 6411 103241 6423 103275
rect 6365 103235 6423 103241
rect 2038 103164 2044 103216
rect 2096 103204 2102 103216
rect 7009 103207 7067 103213
rect 7009 103204 7021 103207
rect 2096 103176 7021 103204
rect 2096 103164 2102 103176
rect 7009 103173 7021 103176
rect 7055 103173 7067 103207
rect 7009 103167 7067 103173
rect 26605 103207 26663 103213
rect 26605 103173 26617 103207
rect 26651 103204 26663 103207
rect 31294 103204 31300 103216
rect 26651 103176 31300 103204
rect 26651 103173 26663 103176
rect 26605 103167 26663 103173
rect 31294 103164 31300 103176
rect 31352 103164 31358 103216
rect 36078 103096 36084 103148
rect 36136 103136 36142 103148
rect 37553 103139 37611 103145
rect 37553 103136 37565 103139
rect 36136 103108 37565 103136
rect 36136 103096 36142 103108
rect 37553 103105 37565 103108
rect 37599 103105 37611 103139
rect 37553 103099 37611 103105
rect 6178 103068 6184 103080
rect 6139 103040 6184 103068
rect 6178 103028 6184 103040
rect 6236 103028 6242 103080
rect 6822 103068 6828 103080
rect 6783 103040 6828 103068
rect 6822 103028 6828 103040
rect 6880 103028 6886 103080
rect 37274 103068 37280 103080
rect 37235 103040 37280 103068
rect 37274 103028 37280 103040
rect 37332 103028 37338 103080
rect 1854 103000 1860 103012
rect 1815 102972 1860 103000
rect 1854 102960 1860 102972
rect 1912 102960 1918 103012
rect 2041 103003 2099 103009
rect 2041 102969 2053 103003
rect 2087 103000 2099 103003
rect 4798 103000 4804 103012
rect 2087 102972 4804 103000
rect 2087 102969 2099 102972
rect 2041 102963 2099 102969
rect 4798 102960 4804 102972
rect 4856 102960 4862 103012
rect 15194 102960 15200 103012
rect 15252 103000 15258 103012
rect 26421 103003 26479 103009
rect 26421 103000 26433 103003
rect 15252 102972 26433 103000
rect 15252 102960 15258 102972
rect 26421 102969 26433 102972
rect 26467 102969 26479 103003
rect 26421 102963 26479 102969
rect 1104 102842 38824 102864
rect 1104 102790 19606 102842
rect 19658 102790 19670 102842
rect 19722 102790 19734 102842
rect 19786 102790 19798 102842
rect 19850 102790 38824 102842
rect 1104 102768 38824 102790
rect 2682 102688 2688 102740
rect 2740 102728 2746 102740
rect 7837 102731 7895 102737
rect 7837 102728 7849 102731
rect 2740 102700 7849 102728
rect 2740 102688 2746 102700
rect 7837 102697 7849 102700
rect 7883 102697 7895 102731
rect 12434 102728 12440 102740
rect 12347 102700 12440 102728
rect 7837 102691 7895 102697
rect 12434 102688 12440 102700
rect 12492 102728 12498 102740
rect 13538 102728 13544 102740
rect 12492 102700 13544 102728
rect 12492 102688 12498 102700
rect 13538 102688 13544 102700
rect 13596 102688 13602 102740
rect 26786 102728 26792 102740
rect 26747 102700 26792 102728
rect 26786 102688 26792 102700
rect 26844 102688 26850 102740
rect 12618 102620 12624 102672
rect 12676 102620 12682 102672
rect 7653 102595 7711 102601
rect 7653 102592 7665 102595
rect 7484 102564 7665 102592
rect 7484 102388 7512 102564
rect 7653 102561 7665 102564
rect 7699 102561 7711 102595
rect 7653 102555 7711 102561
rect 12345 102595 12403 102601
rect 12345 102561 12357 102595
rect 12391 102592 12403 102595
rect 12636 102592 12664 102620
rect 13170 102592 13176 102604
rect 12391 102564 13176 102592
rect 12391 102561 12403 102564
rect 12345 102555 12403 102561
rect 13170 102552 13176 102564
rect 13228 102552 13234 102604
rect 26694 102592 26700 102604
rect 26655 102564 26700 102592
rect 26694 102552 26700 102564
rect 26752 102552 26758 102604
rect 37182 102592 37188 102604
rect 37143 102564 37188 102592
rect 37182 102552 37188 102564
rect 37240 102552 37246 102604
rect 12066 102524 12072 102536
rect 12027 102496 12072 102524
rect 12066 102484 12072 102496
rect 12124 102484 12130 102536
rect 12526 102484 12532 102536
rect 12584 102533 12590 102536
rect 12584 102527 12612 102533
rect 12600 102493 12612 102527
rect 12584 102487 12612 102493
rect 12584 102484 12590 102487
rect 7558 102416 7564 102468
rect 7616 102456 7622 102468
rect 12713 102459 12771 102465
rect 12713 102456 12725 102459
rect 7616 102428 12725 102456
rect 7616 102416 7622 102428
rect 12713 102425 12725 102428
rect 12759 102425 12771 102459
rect 12713 102419 12771 102425
rect 13354 102388 13360 102400
rect 7484 102360 13360 102388
rect 13354 102348 13360 102360
rect 13412 102348 13418 102400
rect 37274 102388 37280 102400
rect 37235 102360 37280 102388
rect 37274 102348 37280 102360
rect 37332 102348 37338 102400
rect 1104 102298 38824 102320
rect 1104 102246 4246 102298
rect 4298 102246 4310 102298
rect 4362 102246 4374 102298
rect 4426 102246 4438 102298
rect 4490 102246 34966 102298
rect 35018 102246 35030 102298
rect 35082 102246 35094 102298
rect 35146 102246 35158 102298
rect 35210 102246 38824 102298
rect 1104 102224 38824 102246
rect 32490 102144 32496 102196
rect 32548 102184 32554 102196
rect 36538 102184 36544 102196
rect 32548 102156 36544 102184
rect 32548 102144 32554 102156
rect 36538 102144 36544 102156
rect 36596 102144 36602 102196
rect 36906 102144 36912 102196
rect 36964 102184 36970 102196
rect 38010 102184 38016 102196
rect 36964 102156 38016 102184
rect 36964 102144 36970 102156
rect 38010 102144 38016 102156
rect 38068 102144 38074 102196
rect 7742 102076 7748 102128
rect 7800 102116 7806 102128
rect 11885 102119 11943 102125
rect 11885 102116 11897 102119
rect 7800 102088 11897 102116
rect 7800 102076 7806 102088
rect 11885 102085 11897 102088
rect 11931 102085 11943 102119
rect 13446 102116 13452 102128
rect 13407 102088 13452 102116
rect 11885 102079 11943 102085
rect 13446 102076 13452 102088
rect 13504 102076 13510 102128
rect 11517 102051 11575 102057
rect 11517 102017 11529 102051
rect 11563 102048 11575 102051
rect 12618 102048 12624 102060
rect 11563 102020 12624 102048
rect 11563 102017 11575 102020
rect 11517 102011 11575 102017
rect 12618 102008 12624 102020
rect 12676 102008 12682 102060
rect 13173 102051 13231 102057
rect 13173 102017 13185 102051
rect 13219 102048 13231 102051
rect 13538 102048 13544 102060
rect 13219 102020 13544 102048
rect 13219 102017 13231 102020
rect 13173 102011 13231 102017
rect 13538 102008 13544 102020
rect 13596 102008 13602 102060
rect 1854 101980 1860 101992
rect 1815 101952 1860 101980
rect 1854 101940 1860 101952
rect 1912 101940 1918 101992
rect 11241 101983 11299 101989
rect 11241 101949 11253 101983
rect 11287 101980 11299 101983
rect 12066 101980 12072 101992
rect 11287 101952 12072 101980
rect 11287 101949 11299 101952
rect 11241 101943 11299 101949
rect 12066 101940 12072 101952
rect 12124 101980 12130 101992
rect 12805 101983 12863 101989
rect 12805 101980 12817 101983
rect 12124 101952 12817 101980
rect 12124 101940 12130 101952
rect 12805 101949 12817 101952
rect 12851 101980 12863 101983
rect 18046 101980 18052 101992
rect 12851 101952 18052 101980
rect 12851 101949 12863 101952
rect 12805 101943 12863 101949
rect 18046 101940 18052 101952
rect 18104 101940 18110 101992
rect 2038 101912 2044 101924
rect 1999 101884 2044 101912
rect 2038 101872 2044 101884
rect 2096 101872 2102 101924
rect 11726 101915 11784 101921
rect 11726 101881 11738 101915
rect 11772 101912 11784 101915
rect 12250 101912 12256 101924
rect 11772 101884 12256 101912
rect 11772 101881 11784 101884
rect 11726 101875 11784 101881
rect 12250 101872 12256 101884
rect 12308 101872 12314 101924
rect 13290 101915 13348 101921
rect 13290 101881 13302 101915
rect 13336 101912 13348 101915
rect 19426 101912 19432 101924
rect 13336 101884 19432 101912
rect 13336 101881 13348 101884
rect 13290 101875 13348 101881
rect 19426 101872 19432 101884
rect 19484 101872 19490 101924
rect 37918 101912 37924 101924
rect 37879 101884 37924 101912
rect 37918 101872 37924 101884
rect 37976 101872 37982 101924
rect 11609 101847 11667 101853
rect 11609 101813 11621 101847
rect 11655 101844 11667 101847
rect 12434 101844 12440 101856
rect 11655 101816 12440 101844
rect 11655 101813 11667 101816
rect 11609 101807 11667 101813
rect 12434 101804 12440 101816
rect 12492 101804 12498 101856
rect 12618 101804 12624 101856
rect 12676 101844 12682 101856
rect 13081 101847 13139 101853
rect 13081 101844 13093 101847
rect 12676 101816 13093 101844
rect 12676 101804 12682 101816
rect 13081 101813 13093 101816
rect 13127 101844 13139 101847
rect 20622 101844 20628 101856
rect 13127 101816 20628 101844
rect 13127 101813 13139 101816
rect 13081 101807 13139 101813
rect 20622 101804 20628 101816
rect 20680 101804 20686 101856
rect 30466 101804 30472 101856
rect 30524 101844 30530 101856
rect 38013 101847 38071 101853
rect 38013 101844 38025 101847
rect 30524 101816 38025 101844
rect 30524 101804 30530 101816
rect 38013 101813 38025 101816
rect 38059 101813 38071 101847
rect 38013 101807 38071 101813
rect 1104 101754 38824 101776
rect 1104 101702 19606 101754
rect 19658 101702 19670 101754
rect 19722 101702 19734 101754
rect 19786 101702 19798 101754
rect 19850 101702 38824 101754
rect 1104 101680 38824 101702
rect 2130 101600 2136 101652
rect 2188 101640 2194 101652
rect 5905 101643 5963 101649
rect 5905 101640 5917 101643
rect 2188 101612 5917 101640
rect 2188 101600 2194 101612
rect 5905 101609 5917 101612
rect 5951 101609 5963 101643
rect 5905 101603 5963 101609
rect 12434 101600 12440 101652
rect 12492 101640 12498 101652
rect 12710 101640 12716 101652
rect 12492 101612 12537 101640
rect 12671 101612 12716 101640
rect 12492 101600 12498 101612
rect 12710 101600 12716 101612
rect 12768 101600 12774 101652
rect 23290 101640 23296 101652
rect 23251 101612 23296 101640
rect 23290 101600 23296 101612
rect 23348 101600 23354 101652
rect 12345 101575 12403 101581
rect 12345 101541 12357 101575
rect 12391 101572 12403 101575
rect 12618 101572 12624 101584
rect 12391 101544 12624 101572
rect 12391 101541 12403 101544
rect 12345 101535 12403 101541
rect 12618 101532 12624 101544
rect 12676 101532 12682 101584
rect 1854 101504 1860 101516
rect 1815 101476 1860 101504
rect 1854 101464 1860 101476
rect 1912 101464 1918 101516
rect 5718 101504 5724 101516
rect 5679 101476 5724 101504
rect 5718 101464 5724 101476
rect 5776 101464 5782 101516
rect 12069 101507 12127 101513
rect 12069 101473 12081 101507
rect 12115 101504 12127 101507
rect 12894 101504 12900 101516
rect 12115 101476 12900 101504
rect 12115 101473 12127 101476
rect 12069 101467 12127 101473
rect 12894 101464 12900 101476
rect 12952 101464 12958 101516
rect 17218 101464 17224 101516
rect 17276 101504 17282 101516
rect 23201 101507 23259 101513
rect 23201 101504 23213 101507
rect 17276 101476 23213 101504
rect 17276 101464 17282 101476
rect 23201 101473 23213 101476
rect 23247 101473 23259 101507
rect 37182 101504 37188 101516
rect 37143 101476 37188 101504
rect 23201 101467 23259 101473
rect 37182 101464 37188 101476
rect 37240 101464 37246 101516
rect 2406 101396 2412 101448
rect 2464 101436 2470 101448
rect 10870 101436 10876 101448
rect 2464 101408 10876 101436
rect 2464 101396 2470 101408
rect 10870 101396 10876 101408
rect 10928 101396 10934 101448
rect 12526 101396 12532 101448
rect 12584 101445 12590 101448
rect 12584 101439 12612 101445
rect 12600 101405 12612 101439
rect 12584 101399 12612 101405
rect 12584 101396 12590 101399
rect 21450 101396 21456 101448
rect 21508 101436 21514 101448
rect 31110 101436 31116 101448
rect 21508 101408 31116 101436
rect 21508 101396 21514 101408
rect 31110 101396 31116 101408
rect 31168 101396 31174 101448
rect 35342 101396 35348 101448
rect 35400 101436 35406 101448
rect 36630 101436 36636 101448
rect 35400 101408 36636 101436
rect 35400 101396 35406 101408
rect 36630 101396 36636 101408
rect 36688 101396 36694 101448
rect 2041 101371 2099 101377
rect 2041 101337 2053 101371
rect 2087 101368 2099 101371
rect 4062 101368 4068 101380
rect 2087 101340 4068 101368
rect 2087 101337 2099 101340
rect 2041 101331 2099 101337
rect 4062 101328 4068 101340
rect 4120 101328 4126 101380
rect 36538 101260 36544 101312
rect 36596 101300 36602 101312
rect 37277 101303 37335 101309
rect 37277 101300 37289 101303
rect 36596 101272 37289 101300
rect 36596 101260 36602 101272
rect 37277 101269 37289 101272
rect 37323 101269 37335 101303
rect 37277 101263 37335 101269
rect 1104 101210 38824 101232
rect 1104 101158 4246 101210
rect 4298 101158 4310 101210
rect 4362 101158 4374 101210
rect 4426 101158 4438 101210
rect 4490 101158 34966 101210
rect 35018 101158 35030 101210
rect 35082 101158 35094 101210
rect 35146 101158 35158 101210
rect 35210 101158 38824 101210
rect 1104 101136 38824 101158
rect 32122 100920 32128 100972
rect 32180 100960 32186 100972
rect 37366 100960 37372 100972
rect 32180 100932 37372 100960
rect 32180 100920 32186 100932
rect 37366 100920 37372 100932
rect 37424 100920 37430 100972
rect 19426 100852 19432 100904
rect 19484 100892 19490 100904
rect 20530 100892 20536 100904
rect 19484 100864 20536 100892
rect 19484 100852 19490 100864
rect 20530 100852 20536 100864
rect 20588 100852 20594 100904
rect 37918 100892 37924 100904
rect 37879 100864 37924 100892
rect 37918 100852 37924 100864
rect 37976 100852 37982 100904
rect 37182 100824 37188 100836
rect 37143 100796 37188 100824
rect 37182 100784 37188 100796
rect 37240 100784 37246 100836
rect 37369 100827 37427 100833
rect 37369 100793 37381 100827
rect 37415 100824 37427 100827
rect 37642 100824 37648 100836
rect 37415 100796 37648 100824
rect 37415 100793 37427 100796
rect 37369 100787 37427 100793
rect 37642 100784 37648 100796
rect 37700 100784 37706 100836
rect 36722 100716 36728 100768
rect 36780 100756 36786 100768
rect 38013 100759 38071 100765
rect 38013 100756 38025 100759
rect 36780 100728 38025 100756
rect 36780 100716 36786 100728
rect 38013 100725 38025 100728
rect 38059 100725 38071 100759
rect 38013 100719 38071 100725
rect 1104 100666 38824 100688
rect 1104 100614 19606 100666
rect 19658 100614 19670 100666
rect 19722 100614 19734 100666
rect 19786 100614 19798 100666
rect 19850 100614 38824 100666
rect 1104 100592 38824 100614
rect 23106 100552 23112 100564
rect 23067 100524 23112 100552
rect 23106 100512 23112 100524
rect 23164 100512 23170 100564
rect 1854 100484 1860 100496
rect 1815 100456 1860 100484
rect 1854 100444 1860 100456
rect 1912 100444 1918 100496
rect 15930 100376 15936 100428
rect 15988 100416 15994 100428
rect 23017 100419 23075 100425
rect 23017 100416 23029 100419
rect 15988 100388 23029 100416
rect 15988 100376 15994 100388
rect 23017 100385 23029 100388
rect 23063 100385 23075 100419
rect 37182 100416 37188 100428
rect 37143 100388 37188 100416
rect 23017 100379 23075 100385
rect 37182 100376 37188 100388
rect 37240 100376 37246 100428
rect 1949 100215 2007 100221
rect 1949 100181 1961 100215
rect 1995 100212 2007 100215
rect 17310 100212 17316 100224
rect 1995 100184 17316 100212
rect 1995 100181 2007 100184
rect 1949 100175 2007 100181
rect 17310 100172 17316 100184
rect 17368 100172 17374 100224
rect 31110 100172 31116 100224
rect 31168 100212 31174 100224
rect 37277 100215 37335 100221
rect 37277 100212 37289 100215
rect 31168 100184 37289 100212
rect 31168 100172 31174 100184
rect 37277 100181 37289 100184
rect 37323 100181 37335 100215
rect 37277 100175 37335 100181
rect 1104 100122 38824 100144
rect 1104 100070 4246 100122
rect 4298 100070 4310 100122
rect 4362 100070 4374 100122
rect 4426 100070 4438 100122
rect 4490 100070 34966 100122
rect 35018 100070 35030 100122
rect 35082 100070 35094 100122
rect 35146 100070 35158 100122
rect 35210 100070 38824 100122
rect 1104 100048 38824 100070
rect 5718 99968 5724 100020
rect 5776 100008 5782 100020
rect 12066 100008 12072 100020
rect 5776 99980 12072 100008
rect 5776 99968 5782 99980
rect 12066 99968 12072 99980
rect 12124 99968 12130 100020
rect 32214 99968 32220 100020
rect 32272 100008 32278 100020
rect 34701 100011 34759 100017
rect 34701 100008 34713 100011
rect 32272 99980 34713 100008
rect 32272 99968 32278 99980
rect 34701 99977 34713 99980
rect 34747 99977 34759 100011
rect 34701 99971 34759 99977
rect 33965 99943 34023 99949
rect 33965 99909 33977 99943
rect 34011 99940 34023 99943
rect 35618 99940 35624 99952
rect 34011 99912 35624 99940
rect 34011 99909 34023 99912
rect 33965 99903 34023 99909
rect 35618 99900 35624 99912
rect 35676 99900 35682 99952
rect 29638 99764 29644 99816
rect 29696 99804 29702 99816
rect 33781 99807 33839 99813
rect 33781 99804 33793 99807
rect 29696 99776 33793 99804
rect 29696 99764 29702 99776
rect 33781 99773 33793 99776
rect 33827 99804 33839 99807
rect 34609 99807 34667 99813
rect 34609 99804 34621 99807
rect 33827 99776 34621 99804
rect 33827 99773 33839 99776
rect 33781 99767 33839 99773
rect 34609 99773 34621 99776
rect 34655 99773 34667 99807
rect 34609 99767 34667 99773
rect 1854 99736 1860 99748
rect 1815 99708 1860 99736
rect 1854 99696 1860 99708
rect 1912 99696 1918 99748
rect 2041 99739 2099 99745
rect 2041 99705 2053 99739
rect 2087 99736 2099 99739
rect 6270 99736 6276 99748
rect 2087 99708 6276 99736
rect 2087 99705 2099 99708
rect 2041 99699 2099 99705
rect 6270 99696 6276 99708
rect 6328 99696 6334 99748
rect 18598 99696 18604 99748
rect 18656 99736 18662 99748
rect 21913 99739 21971 99745
rect 21913 99736 21925 99739
rect 18656 99708 21925 99736
rect 18656 99696 18662 99708
rect 21913 99705 21925 99708
rect 21959 99705 21971 99739
rect 21913 99699 21971 99705
rect 22097 99739 22155 99745
rect 22097 99705 22109 99739
rect 22143 99736 22155 99739
rect 31018 99736 31024 99748
rect 22143 99708 31024 99736
rect 22143 99705 22155 99708
rect 22097 99699 22155 99705
rect 31018 99696 31024 99708
rect 31076 99696 31082 99748
rect 33594 99736 33600 99748
rect 33555 99708 33600 99736
rect 33594 99696 33600 99708
rect 33652 99696 33658 99748
rect 34422 99736 34428 99748
rect 34383 99708 34428 99736
rect 34422 99696 34428 99708
rect 34480 99696 34486 99748
rect 37918 99736 37924 99748
rect 37879 99708 37924 99736
rect 37918 99696 37924 99708
rect 37976 99696 37982 99748
rect 37826 99628 37832 99680
rect 37884 99668 37890 99680
rect 38013 99671 38071 99677
rect 38013 99668 38025 99671
rect 37884 99640 38025 99668
rect 37884 99628 37890 99640
rect 38013 99637 38025 99640
rect 38059 99637 38071 99671
rect 38013 99631 38071 99637
rect 1104 99578 38824 99600
rect 1104 99526 19606 99578
rect 19658 99526 19670 99578
rect 19722 99526 19734 99578
rect 19786 99526 19798 99578
rect 19850 99526 38824 99578
rect 1104 99504 38824 99526
rect 13722 99356 13728 99408
rect 13780 99396 13786 99408
rect 15194 99396 15200 99408
rect 13780 99368 15200 99396
rect 13780 99356 13786 99368
rect 15194 99356 15200 99368
rect 15252 99356 15258 99408
rect 29638 99356 29644 99408
rect 29696 99396 29702 99408
rect 29914 99396 29920 99408
rect 29696 99368 29920 99396
rect 29696 99356 29702 99368
rect 29914 99356 29920 99368
rect 29972 99356 29978 99408
rect 13265 99331 13323 99337
rect 13265 99297 13277 99331
rect 13311 99328 13323 99331
rect 16390 99328 16396 99340
rect 13311 99300 16396 99328
rect 13311 99297 13323 99300
rect 13265 99291 13323 99297
rect 16390 99288 16396 99300
rect 16448 99288 16454 99340
rect 37182 99328 37188 99340
rect 37143 99300 37188 99328
rect 37182 99288 37188 99300
rect 37240 99288 37246 99340
rect 12894 99260 12900 99272
rect 12807 99232 12900 99260
rect 12894 99220 12900 99232
rect 12952 99220 12958 99272
rect 13170 99260 13176 99272
rect 13131 99232 13176 99260
rect 13170 99220 13176 99232
rect 13228 99220 13234 99272
rect 13357 99263 13415 99269
rect 13357 99229 13369 99263
rect 13403 99260 13415 99263
rect 15194 99260 15200 99272
rect 13403 99232 15200 99260
rect 13403 99229 13415 99232
rect 13357 99223 13415 99229
rect 15194 99220 15200 99232
rect 15252 99220 15258 99272
rect 12912 99192 12940 99220
rect 20070 99192 20076 99204
rect 12912 99164 20076 99192
rect 20070 99152 20076 99164
rect 20128 99152 20134 99204
rect 3418 99084 3424 99136
rect 3476 99124 3482 99136
rect 13541 99127 13599 99133
rect 13541 99124 13553 99127
rect 3476 99096 13553 99124
rect 3476 99084 3482 99096
rect 13541 99093 13553 99096
rect 13587 99093 13599 99127
rect 13541 99087 13599 99093
rect 31570 99084 31576 99136
rect 31628 99124 31634 99136
rect 37277 99127 37335 99133
rect 37277 99124 37289 99127
rect 31628 99096 37289 99124
rect 31628 99084 31634 99096
rect 37277 99093 37289 99096
rect 37323 99093 37335 99127
rect 37277 99087 37335 99093
rect 1104 99034 38824 99056
rect 1104 98982 4246 99034
rect 4298 98982 4310 99034
rect 4362 98982 4374 99034
rect 4426 98982 4438 99034
rect 4490 98982 34966 99034
rect 35018 98982 35030 99034
rect 35082 98982 35094 99034
rect 35146 98982 35158 99034
rect 35210 98982 38824 99034
rect 1104 98960 38824 98982
rect 21450 98852 21456 98864
rect 21411 98824 21456 98852
rect 21450 98812 21456 98824
rect 21508 98812 21514 98864
rect 22189 98855 22247 98861
rect 22189 98821 22201 98855
rect 22235 98852 22247 98855
rect 28258 98852 28264 98864
rect 22235 98824 28264 98852
rect 22235 98821 22247 98824
rect 22189 98815 22247 98821
rect 28258 98812 28264 98824
rect 28316 98812 28322 98864
rect 1854 98716 1860 98728
rect 1815 98688 1860 98716
rect 1854 98676 1860 98688
rect 1912 98676 1918 98728
rect 13814 98676 13820 98728
rect 13872 98716 13878 98728
rect 26694 98716 26700 98728
rect 13872 98688 26700 98716
rect 13872 98676 13878 98688
rect 26694 98676 26700 98688
rect 26752 98676 26758 98728
rect 37182 98716 37188 98728
rect 37143 98688 37188 98716
rect 37182 98676 37188 98688
rect 37240 98676 37246 98728
rect 2041 98651 2099 98657
rect 2041 98617 2053 98651
rect 2087 98648 2099 98651
rect 3510 98648 3516 98660
rect 2087 98620 3516 98648
rect 2087 98617 2099 98620
rect 2041 98611 2099 98617
rect 3510 98608 3516 98620
rect 3568 98608 3574 98660
rect 21266 98648 21272 98660
rect 21227 98620 21272 98648
rect 21266 98608 21272 98620
rect 21324 98608 21330 98660
rect 22002 98648 22008 98660
rect 21963 98620 22008 98648
rect 22002 98608 22008 98620
rect 22060 98608 22066 98660
rect 23658 98608 23664 98660
rect 23716 98648 23722 98660
rect 31478 98648 31484 98660
rect 23716 98620 31484 98648
rect 23716 98608 23722 98620
rect 31478 98608 31484 98620
rect 31536 98608 31542 98660
rect 37369 98651 37427 98657
rect 37369 98617 37381 98651
rect 37415 98648 37427 98651
rect 37734 98648 37740 98660
rect 37415 98620 37740 98648
rect 37415 98617 37427 98620
rect 37369 98611 37427 98617
rect 37734 98608 37740 98620
rect 37792 98608 37798 98660
rect 37918 98648 37924 98660
rect 37879 98620 37924 98648
rect 37918 98608 37924 98620
rect 37976 98608 37982 98660
rect 36630 98540 36636 98592
rect 36688 98580 36694 98592
rect 38013 98583 38071 98589
rect 38013 98580 38025 98583
rect 36688 98552 38025 98580
rect 36688 98540 36694 98552
rect 38013 98549 38025 98552
rect 38059 98549 38071 98583
rect 38013 98543 38071 98549
rect 1104 98490 38824 98512
rect 1104 98438 19606 98490
rect 19658 98438 19670 98490
rect 19722 98438 19734 98490
rect 19786 98438 19798 98490
rect 19850 98438 38824 98490
rect 1104 98416 38824 98438
rect 2222 98336 2228 98388
rect 2280 98376 2286 98388
rect 5169 98379 5227 98385
rect 5169 98376 5181 98379
rect 2280 98348 5181 98376
rect 2280 98336 2286 98348
rect 5169 98345 5181 98348
rect 5215 98345 5227 98379
rect 5169 98339 5227 98345
rect 1854 98240 1860 98252
rect 1815 98212 1860 98240
rect 1854 98200 1860 98212
rect 1912 98200 1918 98252
rect 4982 98240 4988 98252
rect 4943 98212 4988 98240
rect 4982 98200 4988 98212
rect 5040 98200 5046 98252
rect 37182 98240 37188 98252
rect 37143 98212 37188 98240
rect 37182 98200 37188 98212
rect 37240 98200 37246 98252
rect 2041 98107 2099 98113
rect 2041 98073 2053 98107
rect 2087 98104 2099 98107
rect 9122 98104 9128 98116
rect 2087 98076 9128 98104
rect 2087 98073 2099 98076
rect 2041 98067 2099 98073
rect 9122 98064 9128 98076
rect 9180 98064 9186 98116
rect 32398 98064 32404 98116
rect 32456 98104 32462 98116
rect 33318 98104 33324 98116
rect 32456 98076 33324 98104
rect 32456 98064 32462 98076
rect 33318 98064 33324 98076
rect 33376 98064 33382 98116
rect 35618 98064 35624 98116
rect 35676 98104 35682 98116
rect 36814 98104 36820 98116
rect 35676 98076 36820 98104
rect 35676 98064 35682 98076
rect 36814 98064 36820 98076
rect 36872 98064 36878 98116
rect 29454 97996 29460 98048
rect 29512 98036 29518 98048
rect 37277 98039 37335 98045
rect 37277 98036 37289 98039
rect 29512 98008 37289 98036
rect 29512 97996 29518 98008
rect 37277 98005 37289 98008
rect 37323 98005 37335 98039
rect 37277 97999 37335 98005
rect 1104 97946 38824 97968
rect 1104 97894 4246 97946
rect 4298 97894 4310 97946
rect 4362 97894 4374 97946
rect 4426 97894 4438 97946
rect 4490 97894 34966 97946
rect 35018 97894 35030 97946
rect 35082 97894 35094 97946
rect 35146 97894 35158 97946
rect 35210 97894 38824 97946
rect 1104 97872 38824 97894
rect 16574 97724 16580 97776
rect 16632 97764 16638 97776
rect 16632 97736 16677 97764
rect 16632 97724 16638 97736
rect 16390 97628 16396 97640
rect 16351 97600 16396 97628
rect 16390 97588 16396 97600
rect 16448 97628 16454 97640
rect 18230 97628 18236 97640
rect 16448 97600 18236 97628
rect 16448 97588 16454 97600
rect 18230 97588 18236 97600
rect 18288 97588 18294 97640
rect 37918 97628 37924 97640
rect 37879 97600 37924 97628
rect 37918 97588 37924 97600
rect 37976 97588 37982 97640
rect 14829 97563 14887 97569
rect 14829 97529 14841 97563
rect 14875 97560 14887 97563
rect 15194 97560 15200 97572
rect 14875 97532 15200 97560
rect 14875 97529 14887 97532
rect 14829 97523 14887 97529
rect 15194 97520 15200 97532
rect 15252 97560 15258 97572
rect 15838 97560 15844 97572
rect 15252 97532 15844 97560
rect 15252 97520 15258 97532
rect 15838 97520 15844 97532
rect 15896 97520 15902 97572
rect 12526 97452 12532 97504
rect 12584 97492 12590 97504
rect 15102 97492 15108 97504
rect 12584 97464 15108 97492
rect 12584 97452 12590 97464
rect 15102 97452 15108 97464
rect 15160 97452 15166 97504
rect 33502 97452 33508 97504
rect 33560 97492 33566 97504
rect 38013 97495 38071 97501
rect 38013 97492 38025 97495
rect 33560 97464 38025 97492
rect 33560 97452 33566 97464
rect 38013 97461 38025 97464
rect 38059 97461 38071 97495
rect 38013 97455 38071 97461
rect 1104 97402 38824 97424
rect 1104 97350 19606 97402
rect 19658 97350 19670 97402
rect 19722 97350 19734 97402
rect 19786 97350 19798 97402
rect 19850 97350 38824 97402
rect 1104 97328 38824 97350
rect 6822 97248 6828 97300
rect 6880 97288 6886 97300
rect 13998 97288 14004 97300
rect 6880 97260 14004 97288
rect 6880 97248 6886 97260
rect 13998 97248 14004 97260
rect 14056 97248 14062 97300
rect 1854 97152 1860 97164
rect 1815 97124 1860 97152
rect 1854 97112 1860 97124
rect 1912 97112 1918 97164
rect 37182 97152 37188 97164
rect 37143 97124 37188 97152
rect 37182 97112 37188 97124
rect 37240 97112 37246 97164
rect 1949 96951 2007 96957
rect 1949 96917 1961 96951
rect 1995 96948 2007 96951
rect 11698 96948 11704 96960
rect 1995 96920 11704 96948
rect 1995 96917 2007 96920
rect 1949 96911 2007 96917
rect 11698 96908 11704 96920
rect 11756 96908 11762 96960
rect 31294 96908 31300 96960
rect 31352 96948 31358 96960
rect 37277 96951 37335 96957
rect 37277 96948 37289 96951
rect 31352 96920 37289 96948
rect 31352 96908 31358 96920
rect 37277 96917 37289 96920
rect 37323 96917 37335 96951
rect 37277 96911 37335 96917
rect 1104 96858 38824 96880
rect 1104 96806 4246 96858
rect 4298 96806 4310 96858
rect 4362 96806 4374 96858
rect 4426 96806 4438 96858
rect 4490 96806 34966 96858
rect 35018 96806 35030 96858
rect 35082 96806 35094 96858
rect 35146 96806 35158 96858
rect 35210 96806 38824 96858
rect 1104 96784 38824 96806
rect 18325 96747 18383 96753
rect 18325 96713 18337 96747
rect 18371 96744 18383 96747
rect 19334 96744 19340 96756
rect 18371 96716 19340 96744
rect 18371 96713 18383 96716
rect 18325 96707 18383 96713
rect 19334 96704 19340 96716
rect 19392 96704 19398 96756
rect 18230 96540 18236 96552
rect 18191 96512 18236 96540
rect 18230 96500 18236 96512
rect 18288 96500 18294 96552
rect 37182 96540 37188 96552
rect 37143 96512 37188 96540
rect 37182 96500 37188 96512
rect 37240 96500 37246 96552
rect 37918 96540 37924 96552
rect 37879 96512 37924 96540
rect 37918 96500 37924 96512
rect 37976 96500 37982 96552
rect 1854 96472 1860 96484
rect 1815 96444 1860 96472
rect 1854 96432 1860 96444
rect 1912 96432 1918 96484
rect 18046 96472 18052 96484
rect 18007 96444 18052 96472
rect 18046 96432 18052 96444
rect 18104 96432 18110 96484
rect 36814 96432 36820 96484
rect 36872 96472 36878 96484
rect 38105 96475 38163 96481
rect 38105 96472 38117 96475
rect 36872 96444 38117 96472
rect 36872 96432 36878 96444
rect 38105 96441 38117 96444
rect 38151 96441 38163 96475
rect 38105 96435 38163 96441
rect 1949 96407 2007 96413
rect 1949 96373 1961 96407
rect 1995 96404 2007 96407
rect 16574 96404 16580 96416
rect 1995 96376 16580 96404
rect 1995 96373 2007 96376
rect 1949 96367 2007 96373
rect 16574 96364 16580 96376
rect 16632 96364 16638 96416
rect 28902 96364 28908 96416
rect 28960 96404 28966 96416
rect 37369 96407 37427 96413
rect 37369 96404 37381 96407
rect 28960 96376 37381 96404
rect 28960 96364 28966 96376
rect 37369 96373 37381 96376
rect 37415 96373 37427 96407
rect 37369 96367 37427 96373
rect 1104 96314 38824 96336
rect 1104 96262 19606 96314
rect 19658 96262 19670 96314
rect 19722 96262 19734 96314
rect 19786 96262 19798 96314
rect 19850 96262 38824 96314
rect 1104 96240 38824 96262
rect 37182 96064 37188 96076
rect 37143 96036 37188 96064
rect 37182 96024 37188 96036
rect 37240 96024 37246 96076
rect 4062 95888 4068 95940
rect 4120 95928 4126 95940
rect 28442 95928 28448 95940
rect 4120 95900 28448 95928
rect 4120 95888 4126 95900
rect 28442 95888 28448 95900
rect 28500 95888 28506 95940
rect 1946 95820 1952 95872
rect 2004 95860 2010 95872
rect 27062 95860 27068 95872
rect 2004 95832 27068 95860
rect 2004 95820 2010 95832
rect 27062 95820 27068 95832
rect 27120 95820 27126 95872
rect 36170 95820 36176 95872
rect 36228 95860 36234 95872
rect 37369 95863 37427 95869
rect 37369 95860 37381 95863
rect 36228 95832 37381 95860
rect 36228 95820 36234 95832
rect 37369 95829 37381 95832
rect 37415 95829 37427 95863
rect 37369 95823 37427 95829
rect 1104 95770 38824 95792
rect 1104 95718 4246 95770
rect 4298 95718 4310 95770
rect 4362 95718 4374 95770
rect 4426 95718 4438 95770
rect 4490 95718 34966 95770
rect 35018 95718 35030 95770
rect 35082 95718 35094 95770
rect 35146 95718 35158 95770
rect 35210 95718 38824 95770
rect 1104 95696 38824 95718
rect 1946 95656 1952 95668
rect 1907 95628 1952 95656
rect 1946 95616 1952 95628
rect 2004 95616 2010 95668
rect 35986 95548 35992 95600
rect 36044 95588 36050 95600
rect 38105 95591 38163 95597
rect 38105 95588 38117 95591
rect 36044 95560 38117 95588
rect 36044 95548 36050 95560
rect 38105 95557 38117 95560
rect 38151 95557 38163 95591
rect 38105 95551 38163 95557
rect 19334 95480 19340 95532
rect 19392 95520 19398 95532
rect 19392 95492 23704 95520
rect 19392 95480 19398 95492
rect 1854 95452 1860 95464
rect 1815 95424 1860 95452
rect 1854 95412 1860 95424
rect 1912 95412 1918 95464
rect 15102 95412 15108 95464
rect 15160 95452 15166 95464
rect 23676 95461 23704 95492
rect 22833 95455 22891 95461
rect 22833 95452 22845 95455
rect 15160 95424 22845 95452
rect 15160 95412 15166 95424
rect 22833 95421 22845 95424
rect 22879 95421 22891 95455
rect 22833 95415 22891 95421
rect 23293 95455 23351 95461
rect 23293 95421 23305 95455
rect 23339 95421 23351 95455
rect 23293 95415 23351 95421
rect 23661 95455 23719 95461
rect 23661 95421 23673 95455
rect 23707 95421 23719 95455
rect 37274 95452 37280 95464
rect 37235 95424 37280 95452
rect 23661 95415 23719 95421
rect 19978 95344 19984 95396
rect 20036 95384 20042 95396
rect 20622 95384 20628 95396
rect 20036 95356 20628 95384
rect 20036 95344 20042 95356
rect 20622 95344 20628 95356
rect 20680 95384 20686 95396
rect 23308 95384 23336 95415
rect 37274 95412 37280 95424
rect 37332 95412 37338 95464
rect 37918 95452 37924 95464
rect 37879 95424 37924 95452
rect 37918 95412 37924 95424
rect 37976 95412 37982 95464
rect 20680 95356 23336 95384
rect 20680 95344 20686 95356
rect 23934 95316 23940 95328
rect 23895 95288 23940 95316
rect 23934 95276 23940 95288
rect 23992 95276 23998 95328
rect 30926 95276 30932 95328
rect 30984 95316 30990 95328
rect 37461 95319 37519 95325
rect 37461 95316 37473 95319
rect 30984 95288 37473 95316
rect 30984 95276 30990 95288
rect 37461 95285 37473 95288
rect 37507 95285 37519 95319
rect 37461 95279 37519 95285
rect 1104 95226 38824 95248
rect 1104 95174 19606 95226
rect 19658 95174 19670 95226
rect 19722 95174 19734 95226
rect 19786 95174 19798 95226
rect 19850 95174 38824 95226
rect 1104 95152 38824 95174
rect 1854 94976 1860 94988
rect 1815 94948 1860 94976
rect 1854 94936 1860 94948
rect 1912 94936 1918 94988
rect 37182 94976 37188 94988
rect 37143 94948 37188 94976
rect 37182 94936 37188 94948
rect 37240 94936 37246 94988
rect 1949 94775 2007 94781
rect 1949 94741 1961 94775
rect 1995 94772 2007 94775
rect 25498 94772 25504 94784
rect 1995 94744 25504 94772
rect 1995 94741 2007 94744
rect 1949 94735 2007 94741
rect 25498 94732 25504 94744
rect 25556 94732 25562 94784
rect 28258 94732 28264 94784
rect 28316 94772 28322 94784
rect 37369 94775 37427 94781
rect 37369 94772 37381 94775
rect 28316 94744 37381 94772
rect 28316 94732 28322 94744
rect 37369 94741 37381 94744
rect 37415 94741 37427 94775
rect 37369 94735 37427 94741
rect 37642 94732 37648 94784
rect 37700 94772 37706 94784
rect 38654 94772 38660 94784
rect 37700 94744 38660 94772
rect 37700 94732 37706 94744
rect 38654 94732 38660 94744
rect 38712 94732 38718 94784
rect 1104 94682 38824 94704
rect 1104 94630 4246 94682
rect 4298 94630 4310 94682
rect 4362 94630 4374 94682
rect 4426 94630 4438 94682
rect 4490 94630 34966 94682
rect 35018 94630 35030 94682
rect 35082 94630 35094 94682
rect 35146 94630 35158 94682
rect 35210 94630 38824 94682
rect 1104 94608 38824 94630
rect 32766 94528 32772 94580
rect 32824 94568 32830 94580
rect 33042 94568 33048 94580
rect 32824 94540 33048 94568
rect 32824 94528 32830 94540
rect 33042 94528 33048 94540
rect 33100 94528 33106 94580
rect 38378 94528 38384 94580
rect 38436 94568 38442 94580
rect 38838 94568 38844 94580
rect 38436 94540 38844 94568
rect 38436 94528 38442 94540
rect 38838 94528 38844 94540
rect 38896 94528 38902 94580
rect 35894 94460 35900 94512
rect 35952 94500 35958 94512
rect 38105 94503 38163 94509
rect 38105 94500 38117 94503
rect 35952 94472 38117 94500
rect 35952 94460 35958 94472
rect 38105 94469 38117 94472
rect 38151 94469 38163 94503
rect 38105 94463 38163 94469
rect 37550 94392 37556 94444
rect 37608 94432 37614 94444
rect 38562 94432 38568 94444
rect 37608 94404 38568 94432
rect 37608 94392 37614 94404
rect 38562 94392 38568 94404
rect 38620 94392 38626 94444
rect 37274 94364 37280 94376
rect 37235 94336 37280 94364
rect 37274 94324 37280 94336
rect 37332 94324 37338 94376
rect 37918 94364 37924 94376
rect 37879 94336 37924 94364
rect 37918 94324 37924 94336
rect 37976 94324 37982 94376
rect 37458 94228 37464 94240
rect 37419 94200 37464 94228
rect 37458 94188 37464 94200
rect 37516 94188 37522 94240
rect 1104 94138 38824 94160
rect 1104 94086 19606 94138
rect 19658 94086 19670 94138
rect 19722 94086 19734 94138
rect 19786 94086 19798 94138
rect 19850 94086 38824 94138
rect 1104 94064 38824 94086
rect 1854 93888 1860 93900
rect 1815 93860 1860 93888
rect 1854 93848 1860 93860
rect 1912 93848 1918 93900
rect 2041 93891 2099 93897
rect 2041 93857 2053 93891
rect 2087 93888 2099 93891
rect 26970 93888 26976 93900
rect 2087 93860 26976 93888
rect 2087 93857 2099 93860
rect 2041 93851 2099 93857
rect 26970 93848 26976 93860
rect 27028 93848 27034 93900
rect 1104 93594 38824 93616
rect 1104 93542 4246 93594
rect 4298 93542 4310 93594
rect 4362 93542 4374 93594
rect 4426 93542 4438 93594
rect 4490 93542 34966 93594
rect 35018 93542 35030 93594
rect 35082 93542 35094 93594
rect 35146 93542 35158 93594
rect 35210 93542 38824 93594
rect 1104 93520 38824 93542
rect 2038 93236 2044 93288
rect 2096 93276 2102 93288
rect 27338 93276 27344 93288
rect 2096 93248 27344 93276
rect 2096 93236 2102 93248
rect 27338 93236 27344 93248
rect 27396 93236 27402 93288
rect 37274 93276 37280 93288
rect 37235 93248 37280 93276
rect 37274 93236 37280 93248
rect 37332 93236 37338 93288
rect 37921 93279 37979 93285
rect 37921 93245 37933 93279
rect 37967 93276 37979 93279
rect 38933 93279 38991 93285
rect 38933 93276 38945 93279
rect 37967 93248 38945 93276
rect 37967 93245 37979 93248
rect 37921 93239 37979 93245
rect 38933 93245 38945 93248
rect 38979 93245 38991 93279
rect 38933 93239 38991 93245
rect 1854 93208 1860 93220
rect 1815 93180 1860 93208
rect 1854 93168 1860 93180
rect 1912 93168 1918 93220
rect 1949 93143 2007 93149
rect 1949 93109 1961 93143
rect 1995 93140 2007 93143
rect 24854 93140 24860 93152
rect 1995 93112 24860 93140
rect 1995 93109 2007 93112
rect 1949 93103 2007 93109
rect 24854 93100 24860 93112
rect 24912 93100 24918 93152
rect 37461 93143 37519 93149
rect 37461 93109 37473 93143
rect 37507 93140 37519 93143
rect 37642 93140 37648 93152
rect 37507 93112 37648 93140
rect 37507 93109 37519 93112
rect 37461 93103 37519 93109
rect 37642 93100 37648 93112
rect 37700 93100 37706 93152
rect 38105 93143 38163 93149
rect 38105 93109 38117 93143
rect 38151 93140 38163 93143
rect 38378 93140 38384 93152
rect 38151 93112 38384 93140
rect 38151 93109 38163 93112
rect 38105 93103 38163 93109
rect 38378 93100 38384 93112
rect 38436 93100 38442 93152
rect 1104 93050 38824 93072
rect 1104 92998 19606 93050
rect 19658 92998 19670 93050
rect 19722 92998 19734 93050
rect 19786 92998 19798 93050
rect 19850 92998 38824 93050
rect 1104 92976 38824 92998
rect 37182 92800 37188 92812
rect 37143 92772 37188 92800
rect 37182 92760 37188 92772
rect 37240 92760 37246 92812
rect 37366 92596 37372 92608
rect 37327 92568 37372 92596
rect 37366 92556 37372 92568
rect 37424 92556 37430 92608
rect 38930 92528 38936 92540
rect 1104 92506 38824 92528
rect 1104 92454 4246 92506
rect 4298 92454 4310 92506
rect 4362 92454 4374 92506
rect 4426 92454 4438 92506
rect 4490 92454 34966 92506
rect 35018 92454 35030 92506
rect 35082 92454 35094 92506
rect 35146 92454 35158 92506
rect 35210 92454 38824 92506
rect 38891 92500 38936 92528
rect 38930 92488 38936 92500
rect 38988 92488 38994 92540
rect 1104 92432 38824 92454
rect 19978 92352 19984 92404
rect 20036 92392 20042 92404
rect 20165 92395 20223 92401
rect 20165 92392 20177 92395
rect 20036 92364 20177 92392
rect 20036 92352 20042 92364
rect 20165 92361 20177 92364
rect 20211 92361 20223 92395
rect 20165 92355 20223 92361
rect 35802 92284 35808 92336
rect 35860 92324 35866 92336
rect 38105 92327 38163 92333
rect 38105 92324 38117 92327
rect 35860 92296 38117 92324
rect 35860 92284 35866 92296
rect 38105 92293 38117 92296
rect 38151 92293 38163 92327
rect 38105 92287 38163 92293
rect 1854 92188 1860 92200
rect 1815 92160 1860 92188
rect 1854 92148 1860 92160
rect 1912 92148 1918 92200
rect 29178 92188 29184 92200
rect 6886 92160 29184 92188
rect 1949 92055 2007 92061
rect 1949 92021 1961 92055
rect 1995 92052 2007 92055
rect 6886 92052 6914 92160
rect 29178 92148 29184 92160
rect 29236 92148 29242 92200
rect 37274 92188 37280 92200
rect 37235 92160 37280 92188
rect 37274 92148 37280 92160
rect 37332 92148 37338 92200
rect 37918 92188 37924 92200
rect 37879 92160 37924 92188
rect 37918 92148 37924 92160
rect 37976 92148 37982 92200
rect 20070 92120 20076 92132
rect 20031 92092 20076 92120
rect 20070 92080 20076 92092
rect 20128 92080 20134 92132
rect 1995 92024 6914 92052
rect 1995 92021 2007 92024
rect 1949 92015 2007 92021
rect 30282 92012 30288 92064
rect 30340 92052 30346 92064
rect 37461 92055 37519 92061
rect 37461 92052 37473 92055
rect 30340 92024 37473 92052
rect 30340 92012 30346 92024
rect 37461 92021 37473 92024
rect 37507 92021 37519 92055
rect 37461 92015 37519 92021
rect 1104 91962 38824 91984
rect 1104 91910 19606 91962
rect 19658 91910 19670 91962
rect 19722 91910 19734 91962
rect 19786 91910 19798 91962
rect 19850 91910 38824 91962
rect 1104 91888 38824 91910
rect 10870 91848 10876 91860
rect 10831 91820 10876 91848
rect 10870 91808 10876 91820
rect 10928 91808 10934 91860
rect 15838 91848 15844 91860
rect 15799 91820 15844 91848
rect 15838 91808 15844 91820
rect 15896 91808 15902 91860
rect 16022 91808 16028 91860
rect 16080 91848 16086 91860
rect 23382 91848 23388 91860
rect 16080 91820 23388 91848
rect 16080 91808 16086 91820
rect 23382 91808 23388 91820
rect 23440 91808 23446 91860
rect 19058 91740 19064 91792
rect 19116 91780 19122 91792
rect 26878 91780 26884 91792
rect 19116 91752 26884 91780
rect 19116 91740 19122 91752
rect 26878 91740 26884 91752
rect 26936 91740 26942 91792
rect 1854 91712 1860 91724
rect 1815 91684 1860 91712
rect 1854 91672 1860 91684
rect 1912 91672 1918 91724
rect 10778 91712 10784 91724
rect 10739 91684 10784 91712
rect 10778 91672 10784 91684
rect 10836 91672 10842 91724
rect 15749 91715 15807 91721
rect 15749 91681 15761 91715
rect 15795 91712 15807 91715
rect 16482 91712 16488 91724
rect 15795 91684 16488 91712
rect 15795 91681 15807 91684
rect 15749 91675 15807 91681
rect 16482 91672 16488 91684
rect 16540 91672 16546 91724
rect 1946 91508 1952 91520
rect 1907 91480 1952 91508
rect 1946 91468 1952 91480
rect 2004 91468 2010 91520
rect 1104 91418 38824 91440
rect 1104 91366 4246 91418
rect 4298 91366 4310 91418
rect 4362 91366 4374 91418
rect 4426 91366 4438 91418
rect 4490 91366 34966 91418
rect 35018 91366 35030 91418
rect 35082 91366 35094 91418
rect 35146 91366 35158 91418
rect 35210 91366 38824 91418
rect 1104 91344 38824 91366
rect 1946 91264 1952 91316
rect 2004 91304 2010 91316
rect 25038 91304 25044 91316
rect 2004 91276 25044 91304
rect 2004 91264 2010 91276
rect 25038 91264 25044 91276
rect 25096 91264 25102 91316
rect 29638 91264 29644 91316
rect 29696 91304 29702 91316
rect 38105 91307 38163 91313
rect 38105 91304 38117 91307
rect 29696 91276 38117 91304
rect 29696 91264 29702 91276
rect 38105 91273 38117 91276
rect 38151 91273 38163 91307
rect 38105 91267 38163 91273
rect 37461 91239 37519 91245
rect 31726 91208 33180 91236
rect 28350 91100 28356 91112
rect 28311 91072 28356 91100
rect 28350 91060 28356 91072
rect 28408 91060 28414 91112
rect 28442 91060 28448 91112
rect 28500 91100 28506 91112
rect 28626 91100 28632 91112
rect 28500 91072 28545 91100
rect 28587 91072 28632 91100
rect 28500 91060 28506 91072
rect 28626 91060 28632 91072
rect 28684 91060 28690 91112
rect 28859 91103 28917 91109
rect 28859 91069 28871 91103
rect 28905 91100 28917 91103
rect 31726 91100 31754 91208
rect 32858 91128 32864 91180
rect 32916 91168 32922 91180
rect 33045 91171 33103 91177
rect 33045 91168 33057 91171
rect 32916 91140 33057 91168
rect 32916 91128 32922 91140
rect 33045 91137 33057 91140
rect 33091 91137 33103 91171
rect 33152 91168 33180 91208
rect 37461 91205 37473 91239
rect 37507 91236 37519 91239
rect 37550 91236 37556 91248
rect 37507 91208 37556 91236
rect 37507 91205 37519 91208
rect 37461 91199 37519 91205
rect 37550 91196 37556 91208
rect 37608 91196 37614 91248
rect 33152 91140 37504 91168
rect 33045 91131 33103 91137
rect 37476 91112 37504 91140
rect 28905 91072 31754 91100
rect 32585 91103 32643 91109
rect 28905 91069 28917 91072
rect 28859 91063 28917 91069
rect 32585 91069 32597 91103
rect 32631 91069 32643 91103
rect 32585 91063 32643 91069
rect 32677 91103 32735 91109
rect 32677 91069 32689 91103
rect 32723 91100 32735 91103
rect 32766 91100 32772 91112
rect 32723 91072 32772 91100
rect 32723 91069 32735 91072
rect 32677 91063 32735 91069
rect 28718 91032 28724 91044
rect 28679 91004 28724 91032
rect 28718 90992 28724 91004
rect 28776 90992 28782 91044
rect 31938 91032 31944 91044
rect 31899 91004 31944 91032
rect 31938 90992 31944 91004
rect 31996 90992 32002 91044
rect 28997 90967 29055 90973
rect 28997 90933 29009 90967
rect 29043 90964 29055 90967
rect 32600 90964 32628 91063
rect 32766 91060 32772 91072
rect 32824 91060 32830 91112
rect 32953 91103 33011 91109
rect 32953 91069 32965 91103
rect 32999 91069 33011 91103
rect 37274 91100 37280 91112
rect 37235 91072 37280 91100
rect 32953 91063 33011 91069
rect 32968 90976 32996 91063
rect 37274 91060 37280 91072
rect 37332 91060 37338 91112
rect 37458 91060 37464 91112
rect 37516 91060 37522 91112
rect 37918 91100 37924 91112
rect 37879 91072 37924 91100
rect 37918 91060 37924 91072
rect 37976 91060 37982 91112
rect 29043 90936 32628 90964
rect 29043 90933 29055 90936
rect 28997 90927 29055 90933
rect 32950 90924 32956 90976
rect 33008 90924 33014 90976
rect 1104 90874 38824 90896
rect 1104 90822 19606 90874
rect 19658 90822 19670 90874
rect 19722 90822 19734 90874
rect 19786 90822 19798 90874
rect 19850 90822 38824 90874
rect 1104 90800 38824 90822
rect 13170 90720 13176 90772
rect 13228 90760 13234 90772
rect 18233 90763 18291 90769
rect 18233 90760 18245 90763
rect 13228 90732 18245 90760
rect 13228 90720 13234 90732
rect 18233 90729 18245 90732
rect 18279 90729 18291 90763
rect 18233 90723 18291 90729
rect 27338 90652 27344 90704
rect 27396 90692 27402 90704
rect 28626 90692 28632 90704
rect 27396 90664 28488 90692
rect 28587 90664 28632 90692
rect 27396 90652 27402 90664
rect 1854 90624 1860 90636
rect 1815 90596 1860 90624
rect 1854 90584 1860 90596
rect 1912 90584 1918 90636
rect 18141 90627 18199 90633
rect 18141 90593 18153 90627
rect 18187 90624 18199 90627
rect 19886 90624 19892 90636
rect 18187 90596 19892 90624
rect 18187 90593 18199 90596
rect 18141 90587 18199 90593
rect 19886 90584 19892 90596
rect 19944 90584 19950 90636
rect 26786 90584 26792 90636
rect 26844 90624 26850 90636
rect 28460 90633 28488 90664
rect 28626 90652 28632 90664
rect 28684 90652 28690 90704
rect 35986 90692 35992 90704
rect 31496 90664 35992 90692
rect 28353 90627 28411 90633
rect 28353 90624 28365 90627
rect 26844 90596 28365 90624
rect 26844 90584 26850 90596
rect 28353 90593 28365 90596
rect 28399 90593 28411 90627
rect 28353 90587 28411 90593
rect 28446 90627 28504 90633
rect 28446 90593 28458 90627
rect 28492 90593 28504 90627
rect 28718 90624 28724 90636
rect 28679 90596 28724 90624
rect 28446 90587 28504 90593
rect 28718 90584 28724 90596
rect 28776 90584 28782 90636
rect 28859 90627 28917 90633
rect 28859 90593 28871 90627
rect 28905 90624 28917 90627
rect 31496 90624 31524 90664
rect 35986 90652 35992 90664
rect 36044 90652 36050 90704
rect 28905 90596 31524 90624
rect 31573 90627 31631 90633
rect 28905 90593 28917 90596
rect 28859 90587 28917 90593
rect 31573 90593 31585 90627
rect 31619 90593 31631 90627
rect 31573 90587 31631 90593
rect 29086 90516 29092 90568
rect 29144 90556 29150 90568
rect 31588 90556 31616 90587
rect 31846 90584 31852 90636
rect 31904 90624 31910 90636
rect 31941 90627 31999 90633
rect 31941 90624 31953 90627
rect 31904 90596 31953 90624
rect 31904 90584 31910 90596
rect 31941 90593 31953 90596
rect 31987 90593 31999 90627
rect 31941 90587 31999 90593
rect 32125 90627 32183 90633
rect 32125 90593 32137 90627
rect 32171 90624 32183 90627
rect 32306 90624 32312 90636
rect 32171 90596 32312 90624
rect 32171 90593 32183 90596
rect 32125 90587 32183 90593
rect 32306 90584 32312 90596
rect 32364 90584 32370 90636
rect 32858 90584 32864 90636
rect 32916 90624 32922 90636
rect 33045 90627 33103 90633
rect 33045 90624 33057 90627
rect 32916 90596 33057 90624
rect 32916 90584 32922 90596
rect 33045 90593 33057 90596
rect 33091 90624 33103 90627
rect 33226 90624 33232 90636
rect 33091 90596 33232 90624
rect 33091 90593 33103 90596
rect 33045 90587 33103 90593
rect 33226 90584 33232 90596
rect 33284 90584 33290 90636
rect 37182 90624 37188 90636
rect 37143 90596 37188 90624
rect 37182 90584 37188 90596
rect 37240 90584 37246 90636
rect 29144 90528 31616 90556
rect 31665 90559 31723 90565
rect 29144 90516 29150 90528
rect 31665 90525 31677 90559
rect 31711 90525 31723 90559
rect 31665 90519 31723 90525
rect 31386 90448 31392 90500
rect 31444 90488 31450 90500
rect 31680 90488 31708 90519
rect 31444 90460 31708 90488
rect 31444 90448 31450 90460
rect 1946 90420 1952 90432
rect 1907 90392 1952 90420
rect 1946 90380 1952 90392
rect 2004 90380 2010 90432
rect 28994 90420 29000 90432
rect 28955 90392 29000 90420
rect 28994 90380 29000 90392
rect 29052 90380 29058 90432
rect 30558 90380 30564 90432
rect 30616 90420 30622 90432
rect 31021 90423 31079 90429
rect 31021 90420 31033 90423
rect 30616 90392 31033 90420
rect 30616 90380 30622 90392
rect 31021 90389 31033 90392
rect 31067 90389 31079 90423
rect 31021 90383 31079 90389
rect 32858 90380 32864 90432
rect 32916 90420 32922 90432
rect 33229 90423 33287 90429
rect 33229 90420 33241 90423
rect 32916 90392 33241 90420
rect 32916 90380 32922 90392
rect 33229 90389 33241 90392
rect 33275 90389 33287 90423
rect 33229 90383 33287 90389
rect 37369 90423 37427 90429
rect 37369 90389 37381 90423
rect 37415 90420 37427 90423
rect 38010 90420 38016 90432
rect 37415 90392 38016 90420
rect 37415 90389 37427 90392
rect 37369 90383 37427 90389
rect 38010 90380 38016 90392
rect 38068 90380 38074 90432
rect 1104 90330 38824 90352
rect 1104 90278 4246 90330
rect 4298 90278 4310 90330
rect 4362 90278 4374 90330
rect 4426 90278 4438 90330
rect 4490 90278 34966 90330
rect 35018 90278 35030 90330
rect 35082 90278 35094 90330
rect 35146 90278 35158 90330
rect 35210 90278 38824 90330
rect 1104 90256 38824 90278
rect 1946 90176 1952 90228
rect 2004 90216 2010 90228
rect 24118 90216 24124 90228
rect 2004 90188 24124 90216
rect 2004 90176 2010 90188
rect 24118 90176 24124 90188
rect 24176 90176 24182 90228
rect 35894 90216 35900 90228
rect 28828 90188 35900 90216
rect 17310 90040 17316 90092
rect 17368 90080 17374 90092
rect 17368 90052 28488 90080
rect 17368 90040 17374 90052
rect 16482 89972 16488 90024
rect 16540 90012 16546 90024
rect 18693 90015 18751 90021
rect 18693 90012 18705 90015
rect 16540 89984 18705 90012
rect 16540 89972 16546 89984
rect 18693 89981 18705 89984
rect 18739 89981 18751 90015
rect 18693 89975 18751 89981
rect 27798 89972 27804 90024
rect 27856 90012 27862 90024
rect 28460 90021 28488 90052
rect 28353 90015 28411 90021
rect 28353 90012 28365 90015
rect 27856 89984 28365 90012
rect 27856 89972 27862 89984
rect 28353 89981 28365 89984
rect 28399 89981 28411 90015
rect 28353 89975 28411 89981
rect 28446 90015 28504 90021
rect 28446 89981 28458 90015
rect 28492 89981 28504 90015
rect 28626 90012 28632 90024
rect 28539 89984 28632 90012
rect 28446 89975 28504 89981
rect 19061 89947 19119 89953
rect 19061 89913 19073 89947
rect 19107 89944 19119 89947
rect 19334 89944 19340 89956
rect 19107 89916 19340 89944
rect 19107 89913 19119 89916
rect 19061 89907 19119 89913
rect 19334 89904 19340 89916
rect 19392 89904 19398 89956
rect 28552 89944 28580 89984
rect 28626 89972 28632 89984
rect 28684 89972 28690 90024
rect 28828 90021 28856 90188
rect 35894 90176 35900 90188
rect 35952 90176 35958 90228
rect 33042 90108 33048 90160
rect 33100 90108 33106 90160
rect 33318 90108 33324 90160
rect 33376 90148 33382 90160
rect 38105 90151 38163 90157
rect 38105 90148 38117 90151
rect 33376 90120 38117 90148
rect 33376 90108 33382 90120
rect 38105 90117 38117 90120
rect 38151 90117 38163 90151
rect 38105 90111 38163 90117
rect 32766 90080 32772 90092
rect 32727 90052 32772 90080
rect 32766 90040 32772 90052
rect 32824 90040 32830 90092
rect 33060 90080 33088 90108
rect 33137 90083 33195 90089
rect 33137 90080 33149 90083
rect 33060 90052 33149 90080
rect 33137 90049 33149 90052
rect 33183 90049 33195 90083
rect 33137 90043 33195 90049
rect 28818 90015 28876 90021
rect 28818 89981 28830 90015
rect 28864 89981 28876 90015
rect 28818 89975 28876 89981
rect 28994 89972 29000 90024
rect 29052 90012 29058 90024
rect 32677 90015 32735 90021
rect 32677 90012 32689 90015
rect 29052 89984 32689 90012
rect 29052 89972 29058 89984
rect 32677 89981 32689 89984
rect 32723 89981 32735 90015
rect 32677 89975 32735 89981
rect 32950 89972 32956 90024
rect 33008 90012 33014 90024
rect 33045 90015 33103 90021
rect 33045 90012 33057 90015
rect 33008 89984 33057 90012
rect 33008 89972 33014 89984
rect 33045 89981 33057 89984
rect 33091 89981 33103 90015
rect 37274 90012 37280 90024
rect 37235 89984 37280 90012
rect 33045 89975 33103 89981
rect 37274 89972 37280 89984
rect 37332 89972 37338 90024
rect 37918 90012 37924 90024
rect 37879 89984 37924 90012
rect 37918 89972 37924 89984
rect 37976 89972 37982 90024
rect 28718 89944 28724 89956
rect 28460 89916 28580 89944
rect 28679 89916 28724 89944
rect 28460 89888 28488 89916
rect 28718 89904 28724 89916
rect 28776 89904 28782 89956
rect 32033 89947 32091 89953
rect 32033 89913 32045 89947
rect 32079 89944 32091 89947
rect 32214 89944 32220 89956
rect 32079 89916 32220 89944
rect 32079 89913 32091 89916
rect 32033 89907 32091 89913
rect 32214 89904 32220 89916
rect 32272 89904 32278 89956
rect 28442 89836 28448 89888
rect 28500 89836 28506 89888
rect 28997 89879 29055 89885
rect 28997 89845 29009 89879
rect 29043 89876 29055 89879
rect 32582 89876 32588 89888
rect 29043 89848 32588 89876
rect 29043 89845 29055 89848
rect 28997 89839 29055 89845
rect 32582 89836 32588 89848
rect 32640 89836 32646 89888
rect 37458 89876 37464 89888
rect 37419 89848 37464 89876
rect 37458 89836 37464 89848
rect 37516 89836 37522 89888
rect 1104 89786 38824 89808
rect 1104 89734 19606 89786
rect 19658 89734 19670 89786
rect 19722 89734 19734 89786
rect 19786 89734 19798 89786
rect 19850 89734 38824 89786
rect 1104 89712 38824 89734
rect 28905 89675 28963 89681
rect 28905 89641 28917 89675
rect 28951 89672 28963 89675
rect 29086 89672 29092 89684
rect 28951 89644 29092 89672
rect 28951 89641 28963 89644
rect 28905 89635 28963 89641
rect 29086 89632 29092 89644
rect 29144 89632 29150 89684
rect 32306 89632 32312 89684
rect 32364 89672 32370 89684
rect 32766 89672 32772 89684
rect 32364 89644 32772 89672
rect 32364 89632 32370 89644
rect 32766 89632 32772 89644
rect 32824 89632 32830 89684
rect 33318 89632 33324 89684
rect 33376 89672 33382 89684
rect 33686 89672 33692 89684
rect 33376 89644 33692 89672
rect 33376 89632 33382 89644
rect 33686 89632 33692 89644
rect 33744 89632 33750 89684
rect 1854 89604 1860 89616
rect 1815 89576 1860 89604
rect 1854 89564 1860 89576
rect 1912 89564 1918 89616
rect 38470 89604 38476 89616
rect 6886 89576 28396 89604
rect 6270 89496 6276 89548
rect 6328 89536 6334 89548
rect 6886 89536 6914 89576
rect 6328 89508 6914 89536
rect 6328 89496 6334 89508
rect 27706 89496 27712 89548
rect 27764 89536 27770 89548
rect 28368 89545 28396 89576
rect 32140 89576 38476 89604
rect 28261 89539 28319 89545
rect 28261 89536 28273 89539
rect 27764 89508 28273 89536
rect 27764 89496 27770 89508
rect 28261 89505 28273 89508
rect 28307 89505 28319 89539
rect 28261 89499 28319 89505
rect 28354 89539 28412 89545
rect 28354 89505 28366 89539
rect 28400 89505 28412 89539
rect 28354 89499 28412 89505
rect 28442 89496 28448 89548
rect 28500 89536 28506 89548
rect 28537 89539 28595 89545
rect 28537 89536 28549 89539
rect 28500 89508 28549 89536
rect 28500 89496 28506 89508
rect 28537 89505 28549 89508
rect 28583 89505 28595 89539
rect 28537 89499 28595 89505
rect 28626 89496 28632 89548
rect 28684 89536 28690 89548
rect 28810 89545 28816 89548
rect 28767 89539 28816 89545
rect 28684 89508 28729 89536
rect 28684 89496 28690 89508
rect 28767 89505 28779 89539
rect 28813 89505 28816 89539
rect 28767 89499 28816 89505
rect 28810 89496 28816 89499
rect 28868 89496 28874 89548
rect 28902 89496 28908 89548
rect 28960 89536 28966 89548
rect 31573 89539 31631 89545
rect 31573 89536 31585 89539
rect 28960 89508 31585 89536
rect 28960 89496 28966 89508
rect 31573 89505 31585 89508
rect 31619 89505 31631 89539
rect 31573 89499 31631 89505
rect 31846 89496 31852 89548
rect 31904 89536 31910 89548
rect 32140 89545 32168 89576
rect 38470 89564 38476 89576
rect 38528 89564 38534 89616
rect 31941 89539 31999 89545
rect 31941 89536 31953 89539
rect 31904 89508 31953 89536
rect 31904 89496 31910 89508
rect 31941 89505 31953 89508
rect 31987 89505 31999 89539
rect 31941 89499 31999 89505
rect 32125 89539 32183 89545
rect 32125 89505 32137 89539
rect 32171 89505 32183 89539
rect 32125 89499 32183 89505
rect 33689 89539 33747 89545
rect 33689 89505 33701 89539
rect 33735 89505 33747 89539
rect 33689 89499 33747 89505
rect 31478 89468 31484 89480
rect 31439 89440 31484 89468
rect 31478 89428 31484 89440
rect 31536 89428 31542 89480
rect 32766 89428 32772 89480
rect 32824 89468 32830 89480
rect 33597 89471 33655 89477
rect 33597 89468 33609 89471
rect 32824 89440 33609 89468
rect 32824 89428 32830 89440
rect 33597 89437 33609 89440
rect 33643 89437 33655 89471
rect 33597 89431 33655 89437
rect 2041 89403 2099 89409
rect 2041 89369 2053 89403
rect 2087 89400 2099 89403
rect 3418 89400 3424 89412
rect 2087 89372 3424 89400
rect 2087 89369 2099 89372
rect 2041 89363 2099 89369
rect 3418 89360 3424 89372
rect 3476 89360 3482 89412
rect 29822 89360 29828 89412
rect 29880 89400 29886 89412
rect 33704 89400 33732 89499
rect 33962 89496 33968 89548
rect 34020 89536 34026 89548
rect 34057 89539 34115 89545
rect 34057 89536 34069 89539
rect 34020 89508 34069 89536
rect 34020 89496 34026 89508
rect 34057 89505 34069 89508
rect 34103 89505 34115 89539
rect 34057 89499 34115 89505
rect 34146 89496 34152 89548
rect 34204 89536 34210 89548
rect 34204 89508 34249 89536
rect 34204 89496 34210 89508
rect 36354 89428 36360 89480
rect 36412 89468 36418 89480
rect 36630 89468 36636 89480
rect 36412 89440 36636 89468
rect 36412 89428 36418 89440
rect 36630 89428 36636 89440
rect 36688 89428 36694 89480
rect 29880 89372 33732 89400
rect 29880 89360 29886 89372
rect 30374 89292 30380 89344
rect 30432 89332 30438 89344
rect 31021 89335 31079 89341
rect 31021 89332 31033 89335
rect 30432 89304 31033 89332
rect 30432 89292 30438 89304
rect 31021 89301 31033 89304
rect 31067 89301 31079 89335
rect 31021 89295 31079 89301
rect 31846 89292 31852 89344
rect 31904 89332 31910 89344
rect 32950 89332 32956 89344
rect 31904 89304 32956 89332
rect 31904 89292 31910 89304
rect 32950 89292 32956 89304
rect 33008 89292 33014 89344
rect 33137 89335 33195 89341
rect 33137 89301 33149 89335
rect 33183 89332 33195 89335
rect 33318 89332 33324 89344
rect 33183 89304 33324 89332
rect 33183 89301 33195 89304
rect 33137 89295 33195 89301
rect 33318 89292 33324 89304
rect 33376 89292 33382 89344
rect 36630 89292 36636 89344
rect 36688 89332 36694 89344
rect 37182 89332 37188 89344
rect 36688 89304 37188 89332
rect 36688 89292 36694 89304
rect 37182 89292 37188 89304
rect 37240 89292 37246 89344
rect 1104 89242 38824 89264
rect 1104 89190 4246 89242
rect 4298 89190 4310 89242
rect 4362 89190 4374 89242
rect 4426 89190 4438 89242
rect 4490 89190 34966 89242
rect 35018 89190 35030 89242
rect 35082 89190 35094 89242
rect 35146 89190 35158 89242
rect 35210 89190 38824 89242
rect 1104 89168 38824 89190
rect 28902 89128 28908 89140
rect 28863 89100 28908 89128
rect 28902 89088 28908 89100
rect 28960 89088 28966 89140
rect 28994 89088 29000 89140
rect 29052 89128 29058 89140
rect 38378 89128 38384 89140
rect 29052 89100 38384 89128
rect 29052 89088 29058 89100
rect 38378 89088 38384 89100
rect 38436 89088 38442 89140
rect 28810 89020 28816 89072
rect 28868 89020 28874 89072
rect 31478 89020 31484 89072
rect 31536 89060 31542 89072
rect 32766 89060 32772 89072
rect 31536 89032 32772 89060
rect 31536 89020 31542 89032
rect 32766 89020 32772 89032
rect 32824 89020 32830 89072
rect 37642 89060 37648 89072
rect 32968 89032 37648 89060
rect 28828 88992 28856 89020
rect 32968 88992 32996 89032
rect 37642 89020 37648 89032
rect 37700 89020 37706 89072
rect 6886 88964 28396 88992
rect 28828 88964 32996 88992
rect 33045 88995 33103 89001
rect 3510 88884 3516 88936
rect 3568 88924 3574 88936
rect 6886 88924 6914 88964
rect 3568 88896 6914 88924
rect 3568 88884 3574 88896
rect 23382 88884 23388 88936
rect 23440 88924 23446 88936
rect 23569 88927 23627 88933
rect 23569 88924 23581 88927
rect 23440 88896 23581 88924
rect 23440 88884 23446 88896
rect 23569 88893 23581 88896
rect 23615 88893 23627 88927
rect 23569 88887 23627 88893
rect 27890 88884 27896 88936
rect 27948 88924 27954 88936
rect 28368 88933 28396 88964
rect 33045 88961 33057 88995
rect 33091 88992 33103 88995
rect 38562 88992 38568 89004
rect 33091 88964 38568 88992
rect 33091 88961 33103 88964
rect 33045 88955 33103 88961
rect 38562 88952 38568 88964
rect 38620 88952 38626 89004
rect 28261 88927 28319 88933
rect 28261 88924 28273 88927
rect 27948 88896 28273 88924
rect 27948 88884 27954 88896
rect 28261 88893 28273 88896
rect 28307 88893 28319 88927
rect 28261 88887 28319 88893
rect 28354 88927 28412 88933
rect 28354 88893 28366 88927
rect 28400 88893 28412 88927
rect 28354 88887 28412 88893
rect 28767 88927 28825 88933
rect 28767 88893 28779 88927
rect 28813 88924 28825 88927
rect 32582 88924 32588 88936
rect 28813 88896 32444 88924
rect 32543 88896 32588 88924
rect 28813 88893 28825 88896
rect 28767 88887 28825 88893
rect 1854 88856 1860 88868
rect 1815 88828 1860 88856
rect 1854 88816 1860 88828
rect 1912 88816 1918 88868
rect 2041 88859 2099 88865
rect 2041 88825 2053 88859
rect 2087 88856 2099 88859
rect 9214 88856 9220 88868
rect 2087 88828 9220 88856
rect 2087 88825 2099 88828
rect 2041 88819 2099 88825
rect 9214 88816 9220 88828
rect 9272 88816 9278 88868
rect 23753 88859 23811 88865
rect 23753 88825 23765 88859
rect 23799 88856 23811 88859
rect 27154 88856 27160 88868
rect 23799 88828 27160 88856
rect 23799 88825 23811 88828
rect 23753 88819 23811 88825
rect 27154 88816 27160 88828
rect 27212 88816 27218 88868
rect 27798 88816 27804 88868
rect 27856 88856 27862 88868
rect 28442 88856 28448 88868
rect 27856 88828 28448 88856
rect 27856 88816 27862 88828
rect 28442 88816 28448 88828
rect 28500 88856 28506 88868
rect 28537 88859 28595 88865
rect 28537 88856 28549 88859
rect 28500 88828 28549 88856
rect 28500 88816 28506 88828
rect 28537 88825 28549 88828
rect 28583 88825 28595 88859
rect 28537 88819 28595 88825
rect 28626 88816 28632 88868
rect 28684 88856 28690 88868
rect 28684 88828 28729 88856
rect 28684 88816 28690 88828
rect 29362 88816 29368 88868
rect 29420 88856 29426 88868
rect 31294 88856 31300 88868
rect 29420 88828 31300 88856
rect 29420 88816 29426 88828
rect 31294 88816 31300 88828
rect 31352 88816 31358 88868
rect 31846 88816 31852 88868
rect 31904 88856 31910 88868
rect 31941 88859 31999 88865
rect 31941 88856 31953 88859
rect 31904 88828 31953 88856
rect 31904 88816 31910 88828
rect 31941 88825 31953 88828
rect 31987 88825 31999 88859
rect 32416 88856 32444 88896
rect 32582 88884 32588 88896
rect 32640 88884 32646 88936
rect 32677 88927 32735 88933
rect 32677 88893 32689 88927
rect 32723 88924 32735 88927
rect 32766 88924 32772 88936
rect 32723 88896 32772 88924
rect 32723 88893 32735 88896
rect 32677 88887 32735 88893
rect 32766 88884 32772 88896
rect 32824 88884 32830 88936
rect 32950 88924 32956 88936
rect 32911 88896 32956 88924
rect 32950 88884 32956 88896
rect 33008 88884 33014 88936
rect 37274 88924 37280 88936
rect 37235 88896 37280 88924
rect 37274 88884 37280 88896
rect 37332 88884 37338 88936
rect 37918 88924 37924 88936
rect 37879 88896 37924 88924
rect 37918 88884 37924 88896
rect 37976 88884 37982 88936
rect 38102 88884 38108 88936
rect 38160 88924 38166 88936
rect 38378 88924 38384 88936
rect 38160 88896 38384 88924
rect 38160 88884 38166 88896
rect 38378 88884 38384 88896
rect 38436 88884 38442 88936
rect 37366 88856 37372 88868
rect 32416 88828 37372 88856
rect 31941 88819 31999 88825
rect 37366 88816 37372 88828
rect 37424 88816 37430 88868
rect 30742 88748 30748 88800
rect 30800 88788 30806 88800
rect 35802 88788 35808 88800
rect 30800 88760 35808 88788
rect 30800 88748 30806 88760
rect 35802 88748 35808 88760
rect 35860 88748 35866 88800
rect 36078 88748 36084 88800
rect 36136 88788 36142 88800
rect 37461 88791 37519 88797
rect 37461 88788 37473 88791
rect 36136 88760 37473 88788
rect 36136 88748 36142 88760
rect 37461 88757 37473 88760
rect 37507 88757 37519 88791
rect 38102 88788 38108 88800
rect 38063 88760 38108 88788
rect 37461 88751 37519 88757
rect 38102 88748 38108 88760
rect 38160 88748 38166 88800
rect 1104 88698 38824 88720
rect 1104 88646 19606 88698
rect 19658 88646 19670 88698
rect 19722 88646 19734 88698
rect 19786 88646 19798 88698
rect 19850 88646 38824 88698
rect 1104 88624 38824 88646
rect 9122 88544 9128 88596
rect 9180 88584 9186 88596
rect 28166 88584 28172 88596
rect 9180 88556 28172 88584
rect 9180 88544 9186 88556
rect 28166 88544 28172 88556
rect 28224 88544 28230 88596
rect 28721 88587 28779 88593
rect 28721 88553 28733 88587
rect 28767 88584 28779 88587
rect 31662 88584 31668 88596
rect 28767 88556 31668 88584
rect 28767 88553 28779 88556
rect 28721 88547 28779 88553
rect 31662 88544 31668 88556
rect 31720 88544 31726 88596
rect 32306 88544 32312 88596
rect 32364 88584 32370 88596
rect 32766 88584 32772 88596
rect 32364 88556 32772 88584
rect 32364 88544 32370 88556
rect 32766 88544 32772 88556
rect 32824 88544 32830 88596
rect 33042 88544 33048 88596
rect 33100 88584 33106 88596
rect 37369 88587 37427 88593
rect 37369 88584 37381 88587
rect 33100 88556 37381 88584
rect 33100 88544 33106 88556
rect 37369 88553 37381 88556
rect 37415 88553 37427 88587
rect 37369 88547 37427 88553
rect 16574 88476 16580 88528
rect 16632 88516 16638 88528
rect 28810 88516 28816 88528
rect 16632 88488 28816 88516
rect 16632 88476 16638 88488
rect 28810 88476 28816 88488
rect 28868 88476 28874 88528
rect 28994 88476 29000 88528
rect 29052 88516 29058 88528
rect 29052 88488 31616 88516
rect 29052 88476 29058 88488
rect 27430 88408 27436 88460
rect 27488 88448 27494 88460
rect 28077 88451 28135 88457
rect 28077 88448 28089 88451
rect 27488 88420 28089 88448
rect 27488 88408 27494 88420
rect 28077 88417 28089 88420
rect 28123 88417 28135 88451
rect 28077 88411 28135 88417
rect 28166 88408 28172 88460
rect 28224 88448 28230 88460
rect 28353 88451 28411 88457
rect 28224 88420 28269 88448
rect 28224 88408 28230 88420
rect 28353 88417 28365 88451
rect 28399 88417 28411 88451
rect 28353 88411 28411 88417
rect 27246 88272 27252 88324
rect 27304 88312 27310 88324
rect 28368 88312 28396 88411
rect 28442 88408 28448 88460
rect 28500 88448 28506 88460
rect 28583 88451 28641 88457
rect 28500 88420 28545 88448
rect 28500 88408 28506 88420
rect 28583 88417 28595 88451
rect 28629 88448 28641 88451
rect 28902 88448 28908 88460
rect 28629 88420 28908 88448
rect 28629 88417 28641 88420
rect 28583 88411 28641 88417
rect 28902 88408 28908 88420
rect 28960 88408 28966 88460
rect 29086 88408 29092 88460
rect 29144 88448 29150 88460
rect 29181 88451 29239 88457
rect 29181 88448 29193 88451
rect 29144 88420 29193 88448
rect 29144 88408 29150 88420
rect 29181 88417 29193 88420
rect 29227 88417 29239 88451
rect 29181 88411 29239 88417
rect 29274 88451 29332 88457
rect 29274 88417 29286 88451
rect 29320 88417 29332 88451
rect 29457 88451 29515 88457
rect 29457 88448 29469 88451
rect 29274 88411 29332 88417
rect 29380 88420 29469 88448
rect 28810 88340 28816 88392
rect 28868 88380 28874 88392
rect 29288 88380 29316 88411
rect 28868 88352 29316 88380
rect 28868 88340 28874 88352
rect 29380 88312 29408 88420
rect 29457 88417 29469 88420
rect 29503 88417 29515 88451
rect 29457 88411 29515 88417
rect 29549 88451 29607 88457
rect 29549 88417 29561 88451
rect 29595 88417 29607 88451
rect 29549 88411 29607 88417
rect 29687 88451 29745 88457
rect 29687 88417 29699 88451
rect 29733 88448 29745 88451
rect 30742 88448 30748 88460
rect 29733 88420 30748 88448
rect 29733 88417 29745 88420
rect 29687 88411 29745 88417
rect 29564 88380 29592 88411
rect 30742 88408 30748 88420
rect 30800 88408 30806 88460
rect 30929 88451 30987 88457
rect 30929 88417 30941 88451
rect 30975 88448 30987 88451
rect 31386 88448 31392 88460
rect 30975 88420 31392 88448
rect 30975 88417 30987 88420
rect 30929 88411 30987 88417
rect 31386 88408 31392 88420
rect 31444 88408 31450 88460
rect 31588 88457 31616 88488
rect 31680 88488 33824 88516
rect 31573 88451 31631 88457
rect 31573 88417 31585 88451
rect 31619 88417 31631 88451
rect 31573 88411 31631 88417
rect 27304 88284 29408 88312
rect 29472 88352 29592 88380
rect 27304 88272 27310 88284
rect 27614 88204 27620 88256
rect 27672 88244 27678 88256
rect 28442 88244 28448 88256
rect 27672 88216 28448 88244
rect 27672 88204 27678 88216
rect 28442 88204 28448 88216
rect 28500 88244 28506 88256
rect 29472 88244 29500 88352
rect 29822 88340 29828 88392
rect 29880 88340 29886 88392
rect 30834 88340 30840 88392
rect 30892 88380 30898 88392
rect 31202 88380 31208 88392
rect 30892 88352 31208 88380
rect 30892 88340 30898 88352
rect 31202 88340 31208 88352
rect 31260 88340 31266 88392
rect 31478 88380 31484 88392
rect 31439 88352 31484 88380
rect 31478 88340 31484 88352
rect 31536 88340 31542 88392
rect 31680 88380 31708 88488
rect 31941 88451 31999 88457
rect 31941 88417 31953 88451
rect 31987 88417 31999 88451
rect 31941 88411 31999 88417
rect 32125 88451 32183 88457
rect 32125 88417 32137 88451
rect 32171 88448 32183 88451
rect 32398 88448 32404 88460
rect 32171 88420 32404 88448
rect 32171 88417 32183 88420
rect 32125 88411 32183 88417
rect 31588 88352 31708 88380
rect 31956 88380 31984 88411
rect 32398 88408 32404 88420
rect 32456 88408 32462 88460
rect 32582 88408 32588 88460
rect 32640 88448 32646 88460
rect 33226 88448 33232 88460
rect 32640 88420 33232 88448
rect 32640 88408 32646 88420
rect 33226 88408 33232 88420
rect 33284 88408 33290 88460
rect 33796 88457 33824 88488
rect 35802 88476 35808 88528
rect 35860 88516 35866 88528
rect 38102 88516 38108 88528
rect 35860 88488 38108 88516
rect 35860 88476 35866 88488
rect 38102 88476 38108 88488
rect 38160 88476 38166 88528
rect 33689 88451 33747 88457
rect 33689 88417 33701 88451
rect 33735 88417 33747 88451
rect 33689 88411 33747 88417
rect 33781 88451 33839 88457
rect 33781 88417 33793 88451
rect 33827 88417 33839 88451
rect 33781 88411 33839 88417
rect 32306 88380 32312 88392
rect 31956 88352 32312 88380
rect 29840 88253 29868 88340
rect 31018 88272 31024 88324
rect 31076 88312 31082 88324
rect 31588 88312 31616 88352
rect 32306 88340 32312 88352
rect 32364 88340 32370 88392
rect 31076 88284 31616 88312
rect 31076 88272 31082 88284
rect 32398 88272 32404 88324
rect 32456 88312 32462 88324
rect 33704 88312 33732 88411
rect 33962 88408 33968 88460
rect 34020 88448 34026 88460
rect 34057 88451 34115 88457
rect 34057 88448 34069 88451
rect 34020 88420 34069 88448
rect 34020 88408 34026 88420
rect 34057 88417 34069 88420
rect 34103 88417 34115 88451
rect 34238 88448 34244 88460
rect 34199 88420 34244 88448
rect 34057 88411 34115 88417
rect 34238 88408 34244 88420
rect 34296 88408 34302 88460
rect 37182 88448 37188 88460
rect 37143 88420 37188 88448
rect 37182 88408 37188 88420
rect 37240 88408 37246 88460
rect 32456 88284 33732 88312
rect 32456 88272 32462 88284
rect 28500 88216 29500 88244
rect 29825 88247 29883 88253
rect 28500 88204 28506 88216
rect 29825 88213 29837 88247
rect 29871 88213 29883 88247
rect 29825 88207 29883 88213
rect 33137 88247 33195 88253
rect 33137 88213 33149 88247
rect 33183 88244 33195 88247
rect 33226 88244 33232 88256
rect 33183 88216 33232 88244
rect 33183 88213 33195 88216
rect 33137 88207 33195 88213
rect 33226 88204 33232 88216
rect 33284 88204 33290 88256
rect 1104 88154 38824 88176
rect 1104 88102 4246 88154
rect 4298 88102 4310 88154
rect 4362 88102 4374 88154
rect 4426 88102 4438 88154
rect 4490 88102 34966 88154
rect 35018 88102 35030 88154
rect 35082 88102 35094 88154
rect 35146 88102 35158 88154
rect 35210 88102 38824 88154
rect 1104 88080 38824 88102
rect 24118 88000 24124 88052
rect 24176 88040 24182 88052
rect 28721 88043 28779 88049
rect 24176 88012 28396 88040
rect 24176 88000 24182 88012
rect 27617 87975 27675 87981
rect 27617 87941 27629 87975
rect 27663 87972 27675 87975
rect 28166 87972 28172 87984
rect 27663 87944 28172 87972
rect 27663 87941 27675 87944
rect 27617 87935 27675 87941
rect 28166 87932 28172 87944
rect 28224 87932 28230 87984
rect 11698 87864 11704 87916
rect 11756 87904 11762 87916
rect 28368 87904 28396 88012
rect 28721 88009 28733 88043
rect 28767 88040 28779 88043
rect 28994 88040 29000 88052
rect 28767 88012 29000 88040
rect 28767 88009 28779 88012
rect 28721 88003 28779 88009
rect 28994 88000 29000 88012
rect 29052 88000 29058 88052
rect 28810 87932 28816 87984
rect 28868 87972 28874 87984
rect 28868 87944 30604 87972
rect 28868 87932 28874 87944
rect 28994 87904 29000 87916
rect 11756 87876 28212 87904
rect 28368 87876 29000 87904
rect 11756 87864 11762 87876
rect 1854 87836 1860 87848
rect 1815 87808 1860 87836
rect 1854 87796 1860 87808
rect 1912 87796 1918 87848
rect 26234 87796 26240 87848
rect 26292 87836 26298 87848
rect 26973 87839 27031 87845
rect 26973 87836 26985 87839
rect 26292 87808 26985 87836
rect 26292 87796 26298 87808
rect 26973 87805 26985 87808
rect 27019 87805 27031 87839
rect 26973 87799 27031 87805
rect 27062 87796 27068 87848
rect 27120 87836 27126 87848
rect 27522 87845 27528 87848
rect 27479 87839 27528 87845
rect 27120 87808 27165 87836
rect 27120 87796 27126 87808
rect 27479 87805 27491 87839
rect 27525 87805 27528 87839
rect 27479 87799 27528 87805
rect 27522 87796 27528 87799
rect 27580 87796 27586 87848
rect 28074 87836 28080 87848
rect 28035 87808 28080 87836
rect 28074 87796 28080 87808
rect 28132 87796 28138 87848
rect 28184 87845 28212 87876
rect 28994 87864 29000 87876
rect 29052 87864 29058 87916
rect 30576 87904 30604 87944
rect 30650 87932 30656 87984
rect 30708 87972 30714 87984
rect 30929 87975 30987 87981
rect 30929 87972 30941 87975
rect 30708 87944 30941 87972
rect 30708 87932 30714 87944
rect 30929 87941 30941 87944
rect 30975 87941 30987 87975
rect 32398 87972 32404 87984
rect 30929 87935 30987 87941
rect 31036 87944 32404 87972
rect 31036 87904 31064 87944
rect 32398 87932 32404 87944
rect 32456 87932 32462 87984
rect 32490 87932 32496 87984
rect 32548 87932 32554 87984
rect 36170 87932 36176 87984
rect 36228 87972 36234 87984
rect 38105 87975 38163 87981
rect 38105 87972 38117 87975
rect 36228 87944 38117 87972
rect 36228 87932 36234 87944
rect 38105 87941 38117 87944
rect 38151 87941 38163 87975
rect 38105 87935 38163 87941
rect 30576 87876 31064 87904
rect 31478 87864 31484 87916
rect 31536 87904 31542 87916
rect 32033 87907 32091 87913
rect 32033 87904 32045 87907
rect 31536 87876 32045 87904
rect 31536 87864 31542 87876
rect 32033 87873 32045 87876
rect 32079 87873 32091 87907
rect 32508 87904 32536 87932
rect 32585 87907 32643 87913
rect 32585 87904 32597 87907
rect 32508 87876 32597 87904
rect 32033 87867 32091 87873
rect 32585 87873 32597 87876
rect 32631 87873 32643 87907
rect 32585 87867 32643 87873
rect 28170 87839 28228 87845
rect 28170 87805 28182 87839
rect 28216 87805 28228 87839
rect 28170 87799 28228 87805
rect 28583 87839 28641 87845
rect 28583 87805 28595 87839
rect 28629 87836 28641 87839
rect 30282 87836 30288 87848
rect 28629 87808 30288 87836
rect 28629 87805 28641 87808
rect 28583 87799 28641 87805
rect 30282 87796 30288 87808
rect 30340 87796 30346 87848
rect 30745 87839 30803 87845
rect 30745 87805 30757 87839
rect 30791 87836 30803 87839
rect 30791 87808 31616 87836
rect 30791 87805 30803 87808
rect 30745 87799 30803 87805
rect 2041 87771 2099 87777
rect 2041 87737 2053 87771
rect 2087 87768 2099 87771
rect 3510 87768 3516 87780
rect 2087 87740 3516 87768
rect 2087 87737 2099 87740
rect 2041 87731 2099 87737
rect 3510 87728 3516 87740
rect 3568 87728 3574 87780
rect 27246 87768 27252 87780
rect 27207 87740 27252 87768
rect 27246 87728 27252 87740
rect 27304 87728 27310 87780
rect 27341 87771 27399 87777
rect 27341 87737 27353 87771
rect 27387 87768 27399 87771
rect 27614 87768 27620 87780
rect 27387 87740 27620 87768
rect 27387 87737 27399 87740
rect 27341 87731 27399 87737
rect 27614 87728 27620 87740
rect 27672 87728 27678 87780
rect 28353 87771 28411 87777
rect 28353 87768 28365 87771
rect 27724 87740 28365 87768
rect 27264 87700 27292 87728
rect 27724 87700 27752 87740
rect 28353 87737 28365 87740
rect 28399 87737 28411 87771
rect 28353 87731 28411 87737
rect 28442 87728 28448 87780
rect 28500 87768 28506 87780
rect 28810 87768 28816 87780
rect 28500 87740 28816 87768
rect 28500 87728 28506 87740
rect 28810 87728 28816 87740
rect 28868 87728 28874 87780
rect 31294 87728 31300 87780
rect 31352 87768 31358 87780
rect 31481 87771 31539 87777
rect 31481 87768 31493 87771
rect 31352 87740 31493 87768
rect 31352 87728 31358 87740
rect 31481 87737 31493 87740
rect 31527 87737 31539 87771
rect 31588 87768 31616 87808
rect 31662 87796 31668 87848
rect 31720 87836 31726 87848
rect 32125 87839 32183 87845
rect 32125 87836 32137 87839
rect 31720 87808 32137 87836
rect 31720 87796 31726 87808
rect 32125 87805 32137 87808
rect 32171 87805 32183 87839
rect 32125 87799 32183 87805
rect 32306 87796 32312 87848
rect 32364 87836 32370 87848
rect 32493 87839 32551 87845
rect 32493 87836 32505 87839
rect 32364 87808 32505 87836
rect 32364 87796 32370 87808
rect 32493 87805 32505 87808
rect 32539 87836 32551 87839
rect 33962 87836 33968 87848
rect 32539 87808 33968 87836
rect 32539 87805 32551 87808
rect 32493 87799 32551 87805
rect 33962 87796 33968 87808
rect 34020 87796 34026 87848
rect 34146 87796 34152 87848
rect 34204 87836 34210 87848
rect 35894 87836 35900 87848
rect 34204 87808 35900 87836
rect 34204 87796 34210 87808
rect 35894 87796 35900 87808
rect 35952 87796 35958 87848
rect 37274 87836 37280 87848
rect 37235 87808 37280 87836
rect 37274 87796 37280 87808
rect 37332 87796 37338 87848
rect 37918 87836 37924 87848
rect 37879 87808 37924 87836
rect 37918 87796 37924 87808
rect 37976 87796 37982 87848
rect 32582 87768 32588 87780
rect 31588 87740 32588 87768
rect 31481 87731 31539 87737
rect 32582 87728 32588 87740
rect 32640 87768 32646 87780
rect 33229 87771 33287 87777
rect 33229 87768 33241 87771
rect 32640 87740 33241 87768
rect 32640 87728 32646 87740
rect 33229 87737 33241 87740
rect 33275 87737 33287 87771
rect 33229 87731 33287 87737
rect 27264 87672 27752 87700
rect 28166 87660 28172 87712
rect 28224 87700 28230 87712
rect 32398 87700 32404 87712
rect 28224 87672 32404 87700
rect 28224 87660 28230 87672
rect 32398 87660 32404 87672
rect 32456 87660 32462 87712
rect 32490 87660 32496 87712
rect 32548 87700 32554 87712
rect 33321 87703 33379 87709
rect 33321 87700 33333 87703
rect 32548 87672 33333 87700
rect 32548 87660 32554 87672
rect 33321 87669 33333 87672
rect 33367 87669 33379 87703
rect 33321 87663 33379 87669
rect 35894 87660 35900 87712
rect 35952 87700 35958 87712
rect 37461 87703 37519 87709
rect 37461 87700 37473 87703
rect 35952 87672 37473 87700
rect 35952 87660 35958 87672
rect 37461 87669 37473 87672
rect 37507 87669 37519 87703
rect 37461 87663 37519 87669
rect 1104 87610 38824 87632
rect 1104 87558 19606 87610
rect 19658 87558 19670 87610
rect 19722 87558 19734 87610
rect 19786 87558 19798 87610
rect 19850 87558 38824 87610
rect 1104 87536 38824 87558
rect 26142 87456 26148 87508
rect 26200 87496 26206 87508
rect 28629 87499 28687 87505
rect 26200 87468 28488 87496
rect 26200 87456 26206 87468
rect 9030 87388 9036 87440
rect 9088 87428 9094 87440
rect 9088 87400 28120 87428
rect 9088 87388 9094 87400
rect 1854 87360 1860 87372
rect 1815 87332 1860 87360
rect 1854 87320 1860 87332
rect 1912 87320 1918 87372
rect 23382 87360 23388 87372
rect 23343 87332 23388 87360
rect 23382 87320 23388 87332
rect 23440 87320 23446 87372
rect 27338 87320 27344 87372
rect 27396 87360 27402 87372
rect 28092 87369 28120 87400
rect 28166 87388 28172 87440
rect 28224 87428 28230 87440
rect 28353 87431 28411 87437
rect 28353 87428 28365 87431
rect 28224 87400 28365 87428
rect 28224 87388 28230 87400
rect 28353 87397 28365 87400
rect 28399 87397 28411 87431
rect 28460 87428 28488 87468
rect 28629 87465 28641 87499
rect 28675 87496 28687 87499
rect 31202 87496 31208 87508
rect 28675 87468 31208 87496
rect 28675 87465 28687 87468
rect 28629 87459 28687 87465
rect 31202 87456 31208 87468
rect 31260 87456 31266 87508
rect 32950 87456 32956 87508
rect 33008 87496 33014 87508
rect 33229 87499 33287 87505
rect 33229 87496 33241 87499
rect 33008 87468 33241 87496
rect 33008 87456 33014 87468
rect 33229 87465 33241 87468
rect 33275 87465 33287 87499
rect 33229 87459 33287 87465
rect 33962 87456 33968 87508
rect 34020 87496 34026 87508
rect 36998 87496 37004 87508
rect 34020 87468 37004 87496
rect 34020 87456 34026 87468
rect 36998 87456 37004 87468
rect 37056 87456 37062 87508
rect 29273 87431 29331 87437
rect 29273 87428 29285 87431
rect 28460 87400 29285 87428
rect 28353 87391 28411 87397
rect 29273 87397 29285 87400
rect 29319 87397 29331 87431
rect 30926 87428 30932 87440
rect 29273 87391 29331 87397
rect 29472 87400 30932 87428
rect 27985 87363 28043 87369
rect 27985 87360 27997 87363
rect 27396 87332 27997 87360
rect 27396 87320 27402 87332
rect 27985 87329 27997 87332
rect 28031 87329 28043 87363
rect 27985 87323 28043 87329
rect 28078 87363 28136 87369
rect 28078 87329 28090 87363
rect 28124 87329 28136 87363
rect 28078 87323 28136 87329
rect 28261 87363 28319 87369
rect 28261 87329 28273 87363
rect 28307 87329 28319 87363
rect 28261 87323 28319 87329
rect 28491 87363 28549 87369
rect 28491 87329 28503 87363
rect 28537 87360 28549 87363
rect 29472 87360 29500 87400
rect 30926 87388 30932 87400
rect 30984 87388 30990 87440
rect 32398 87388 32404 87440
rect 32456 87428 32462 87440
rect 37550 87428 37556 87440
rect 32456 87400 37556 87428
rect 32456 87388 32462 87400
rect 37550 87388 37556 87400
rect 37608 87388 37614 87440
rect 28537 87332 29500 87360
rect 28537 87329 28549 87332
rect 28491 87323 28549 87329
rect 28276 87292 28304 87323
rect 29546 87320 29552 87372
rect 29604 87360 29610 87372
rect 29917 87363 29975 87369
rect 29917 87360 29929 87363
rect 29604 87332 29929 87360
rect 29604 87320 29610 87332
rect 29917 87329 29929 87332
rect 29963 87329 29975 87363
rect 29917 87323 29975 87329
rect 30285 87363 30343 87369
rect 30285 87329 30297 87363
rect 30331 87329 30343 87363
rect 30285 87323 30343 87329
rect 30469 87363 30527 87369
rect 30469 87329 30481 87363
rect 30515 87360 30527 87363
rect 30834 87360 30840 87372
rect 30515 87332 30840 87360
rect 30515 87329 30527 87332
rect 30469 87323 30527 87329
rect 28902 87292 28908 87304
rect 28276 87264 28908 87292
rect 28902 87252 28908 87264
rect 28960 87252 28966 87304
rect 30009 87295 30067 87301
rect 30009 87261 30021 87295
rect 30055 87292 30067 87295
rect 30098 87292 30104 87304
rect 30055 87264 30104 87292
rect 30055 87261 30067 87264
rect 30009 87255 30067 87261
rect 30098 87252 30104 87264
rect 30156 87252 30162 87304
rect 30300 87292 30328 87323
rect 30834 87320 30840 87332
rect 30892 87320 30898 87372
rect 31573 87363 31631 87369
rect 31573 87360 31585 87363
rect 30944 87332 31585 87360
rect 30300 87264 30512 87292
rect 23569 87227 23627 87233
rect 23569 87193 23581 87227
rect 23615 87224 23627 87227
rect 28718 87224 28724 87236
rect 23615 87196 28724 87224
rect 23615 87193 23627 87196
rect 23569 87187 23627 87193
rect 28718 87184 28724 87196
rect 28776 87184 28782 87236
rect 30484 87224 30512 87264
rect 30742 87252 30748 87304
rect 30800 87292 30806 87304
rect 30944 87292 30972 87332
rect 31573 87329 31585 87332
rect 31619 87329 31631 87363
rect 31573 87323 31631 87329
rect 31941 87363 31999 87369
rect 31941 87329 31953 87363
rect 31987 87360 31999 87363
rect 32306 87360 32312 87372
rect 31987 87332 32312 87360
rect 31987 87329 31999 87332
rect 31941 87323 31999 87329
rect 32306 87320 32312 87332
rect 32364 87320 32370 87372
rect 32490 87320 32496 87372
rect 32548 87360 32554 87372
rect 32950 87360 32956 87372
rect 32548 87332 32956 87360
rect 32548 87320 32554 87332
rect 32950 87320 32956 87332
rect 33008 87360 33014 87372
rect 33045 87363 33103 87369
rect 33045 87360 33057 87363
rect 33008 87332 33057 87360
rect 33008 87320 33014 87332
rect 33045 87329 33057 87332
rect 33091 87329 33103 87363
rect 33045 87323 33103 87329
rect 34606 87320 34612 87372
rect 34664 87320 34670 87372
rect 35250 87320 35256 87372
rect 35308 87360 35314 87372
rect 35434 87360 35440 87372
rect 35308 87332 35440 87360
rect 35308 87320 35314 87332
rect 35434 87320 35440 87332
rect 35492 87320 35498 87372
rect 30800 87264 30972 87292
rect 30800 87252 30806 87264
rect 31018 87252 31024 87304
rect 31076 87292 31082 87304
rect 31481 87295 31539 87301
rect 31481 87292 31493 87295
rect 31076 87264 31493 87292
rect 31076 87252 31082 87264
rect 31481 87261 31493 87264
rect 31527 87261 31539 87295
rect 31481 87255 31539 87261
rect 32033 87295 32091 87301
rect 32033 87261 32045 87295
rect 32079 87292 32091 87295
rect 33962 87292 33968 87304
rect 32079 87264 33968 87292
rect 32079 87261 32091 87264
rect 32033 87255 32091 87261
rect 33962 87252 33968 87264
rect 34020 87252 34026 87304
rect 34624 87236 34652 87320
rect 30484 87196 31156 87224
rect 1946 87156 1952 87168
rect 1907 87128 1952 87156
rect 1946 87116 1952 87128
rect 2004 87116 2010 87168
rect 28258 87116 28264 87168
rect 28316 87156 28322 87168
rect 28534 87156 28540 87168
rect 28316 87128 28540 87156
rect 28316 87116 28322 87128
rect 28534 87116 28540 87128
rect 28592 87116 28598 87168
rect 29270 87116 29276 87168
rect 29328 87156 29334 87168
rect 30742 87156 30748 87168
rect 29328 87128 30748 87156
rect 29328 87116 29334 87128
rect 30742 87116 30748 87128
rect 30800 87116 30806 87168
rect 30834 87116 30840 87168
rect 30892 87156 30898 87168
rect 31021 87159 31079 87165
rect 31021 87156 31033 87159
rect 30892 87128 31033 87156
rect 30892 87116 30898 87128
rect 31021 87125 31033 87128
rect 31067 87125 31079 87159
rect 31128 87156 31156 87196
rect 34606 87184 34612 87236
rect 34664 87184 34670 87236
rect 35158 87184 35164 87236
rect 35216 87224 35222 87236
rect 35216 87196 35296 87224
rect 35216 87184 35222 87196
rect 35268 87168 35296 87196
rect 32398 87156 32404 87168
rect 31128 87128 32404 87156
rect 31021 87119 31079 87125
rect 32398 87116 32404 87128
rect 32456 87156 32462 87168
rect 32858 87156 32864 87168
rect 32456 87128 32864 87156
rect 32456 87116 32462 87128
rect 32858 87116 32864 87128
rect 32916 87116 32922 87168
rect 35250 87116 35256 87168
rect 35308 87116 35314 87168
rect 1104 87066 38824 87088
rect 1104 87014 4246 87066
rect 4298 87014 4310 87066
rect 4362 87014 4374 87066
rect 4426 87014 4438 87066
rect 4490 87014 34966 87066
rect 35018 87014 35030 87066
rect 35082 87014 35094 87066
rect 35146 87014 35158 87066
rect 35210 87014 38824 87066
rect 1104 86992 38824 87014
rect 4798 86912 4804 86964
rect 4856 86952 4862 86964
rect 26789 86955 26847 86961
rect 26789 86952 26801 86955
rect 4856 86924 26801 86952
rect 4856 86912 4862 86924
rect 26789 86921 26801 86924
rect 26835 86921 26847 86955
rect 26789 86915 26847 86921
rect 27525 86955 27583 86961
rect 27525 86921 27537 86955
rect 27571 86952 27583 86955
rect 27614 86952 27620 86964
rect 27571 86924 27620 86952
rect 27571 86921 27583 86924
rect 27525 86915 27583 86921
rect 27614 86912 27620 86924
rect 27672 86912 27678 86964
rect 32490 86952 32496 86964
rect 27816 86924 32496 86952
rect 20070 86776 20076 86828
rect 20128 86816 20134 86828
rect 20128 86788 23244 86816
rect 20128 86776 20134 86788
rect 19334 86708 19340 86760
rect 19392 86748 19398 86760
rect 23216 86757 23244 86788
rect 24854 86776 24860 86828
rect 24912 86816 24918 86828
rect 27522 86816 27528 86828
rect 24912 86788 27016 86816
rect 24912 86776 24918 86788
rect 23017 86751 23075 86757
rect 23017 86748 23029 86751
rect 19392 86720 23029 86748
rect 19392 86708 19398 86720
rect 23017 86717 23029 86720
rect 23063 86717 23075 86751
rect 23017 86711 23075 86717
rect 23201 86751 23259 86757
rect 23201 86717 23213 86751
rect 23247 86717 23259 86751
rect 23201 86711 23259 86717
rect 23382 86708 23388 86760
rect 23440 86748 23446 86760
rect 23937 86751 23995 86757
rect 23937 86748 23949 86751
rect 23440 86720 23949 86748
rect 23440 86708 23446 86720
rect 23937 86717 23949 86720
rect 23983 86717 23995 86751
rect 23937 86711 23995 86717
rect 26602 86708 26608 86760
rect 26660 86748 26666 86760
rect 26988 86757 27016 86788
rect 27264 86788 27528 86816
rect 26881 86751 26939 86757
rect 26881 86748 26893 86751
rect 26660 86720 26893 86748
rect 26660 86708 26666 86720
rect 26881 86717 26893 86720
rect 26927 86717 26939 86751
rect 26881 86711 26939 86717
rect 26974 86751 27032 86757
rect 26974 86717 26986 86751
rect 27020 86717 27032 86751
rect 27154 86748 27160 86760
rect 27115 86720 27160 86748
rect 26974 86711 27032 86717
rect 27154 86708 27160 86720
rect 27212 86708 27218 86760
rect 27264 86757 27292 86788
rect 27522 86776 27528 86788
rect 27580 86776 27586 86828
rect 27249 86751 27307 86757
rect 27249 86717 27261 86751
rect 27295 86717 27307 86751
rect 27249 86711 27307 86717
rect 27387 86751 27445 86757
rect 27387 86717 27399 86751
rect 27433 86748 27445 86751
rect 27816 86748 27844 86924
rect 32490 86912 32496 86924
rect 32548 86912 32554 86964
rect 32582 86912 32588 86964
rect 32640 86952 32646 86964
rect 32640 86924 33824 86952
rect 32640 86912 32646 86924
rect 28166 86844 28172 86896
rect 28224 86884 28230 86896
rect 28224 86856 28396 86884
rect 28224 86844 28230 86856
rect 28258 86816 28264 86828
rect 28000 86788 28264 86816
rect 28000 86757 28028 86788
rect 28258 86776 28264 86788
rect 28316 86776 28322 86828
rect 28368 86757 28396 86856
rect 30098 86844 30104 86896
rect 30156 86884 30162 86896
rect 31018 86884 31024 86896
rect 30156 86856 31024 86884
rect 30156 86844 30162 86856
rect 31018 86844 31024 86856
rect 31076 86884 31082 86896
rect 31662 86884 31668 86896
rect 31076 86856 31668 86884
rect 31076 86844 31082 86856
rect 28902 86816 28908 86828
rect 28828 86788 28908 86816
rect 28534 86757 28540 86760
rect 27433 86720 27844 86748
rect 27985 86751 28043 86757
rect 27433 86717 27445 86720
rect 27387 86711 27445 86717
rect 27985 86717 27997 86751
rect 28031 86717 28043 86751
rect 27985 86711 28043 86717
rect 28078 86751 28136 86757
rect 28078 86717 28090 86751
rect 28124 86717 28136 86751
rect 28078 86711 28136 86717
rect 28353 86751 28411 86757
rect 28353 86717 28365 86751
rect 28399 86717 28411 86751
rect 28353 86711 28411 86717
rect 28491 86751 28540 86757
rect 28491 86717 28503 86751
rect 28537 86717 28540 86751
rect 28491 86711 28540 86717
rect 19426 86640 19432 86692
rect 19484 86680 19490 86692
rect 20162 86680 20168 86692
rect 19484 86652 20168 86680
rect 19484 86640 19490 86652
rect 20162 86640 20168 86652
rect 20220 86680 20226 86692
rect 22557 86683 22615 86689
rect 22557 86680 22569 86683
rect 20220 86652 22569 86680
rect 20220 86640 20226 86652
rect 22557 86649 22569 86652
rect 22603 86649 22615 86683
rect 22557 86643 22615 86649
rect 22649 86683 22707 86689
rect 22649 86649 22661 86683
rect 22695 86680 22707 86683
rect 22738 86680 22744 86692
rect 22695 86652 22744 86680
rect 22695 86649 22707 86652
rect 22649 86643 22707 86649
rect 22738 86640 22744 86652
rect 22796 86640 22802 86692
rect 23109 86683 23167 86689
rect 23109 86649 23121 86683
rect 23155 86649 23167 86683
rect 23109 86643 23167 86649
rect 24121 86683 24179 86689
rect 24121 86649 24133 86683
rect 24167 86680 24179 86683
rect 26694 86680 26700 86692
rect 24167 86652 26700 86680
rect 24167 86649 24179 86652
rect 24121 86643 24179 86649
rect 18230 86572 18236 86624
rect 18288 86612 18294 86624
rect 19334 86612 19340 86624
rect 18288 86584 19340 86612
rect 18288 86572 18294 86584
rect 19334 86572 19340 86584
rect 19392 86612 19398 86624
rect 23124 86612 23152 86643
rect 26694 86640 26700 86652
rect 26752 86640 26758 86692
rect 26789 86683 26847 86689
rect 26789 86649 26801 86683
rect 26835 86680 26847 86683
rect 28093 86680 28121 86711
rect 28534 86708 28540 86711
rect 28592 86708 28598 86760
rect 26835 86652 28121 86680
rect 28261 86683 28319 86689
rect 26835 86649 26847 86652
rect 26789 86643 26847 86649
rect 28261 86649 28273 86683
rect 28307 86680 28319 86683
rect 28828 86680 28856 86788
rect 28902 86776 28908 86788
rect 28960 86776 28966 86828
rect 31588 86825 31616 86856
rect 31662 86844 31668 86856
rect 31720 86844 31726 86896
rect 32766 86844 32772 86896
rect 32824 86884 32830 86896
rect 32950 86884 32956 86896
rect 32824 86856 32956 86884
rect 32824 86844 32830 86856
rect 32950 86844 32956 86856
rect 33008 86884 33014 86896
rect 33008 86856 33272 86884
rect 33008 86844 33014 86856
rect 31573 86819 31631 86825
rect 31573 86785 31585 86819
rect 31619 86785 31631 86819
rect 32122 86816 32128 86828
rect 32083 86788 32128 86816
rect 31573 86779 31631 86785
rect 32122 86776 32128 86788
rect 32180 86776 32186 86828
rect 32508 86788 33180 86816
rect 28966 86720 29096 86748
rect 28966 86692 28994 86720
rect 28307 86652 28856 86680
rect 28307 86649 28319 86652
rect 28261 86643 28319 86649
rect 28552 86624 28580 86652
rect 28902 86640 28908 86692
rect 28960 86652 28994 86692
rect 29068 86680 29096 86720
rect 29822 86708 29828 86760
rect 29880 86748 29886 86760
rect 31665 86751 31723 86757
rect 31665 86748 31677 86751
rect 29880 86720 31677 86748
rect 29880 86708 29886 86720
rect 31665 86717 31677 86720
rect 31711 86717 31723 86751
rect 31665 86711 31723 86717
rect 32033 86751 32091 86757
rect 32033 86717 32045 86751
rect 32079 86748 32091 86751
rect 32398 86748 32404 86760
rect 32079 86720 32404 86748
rect 32079 86717 32091 86720
rect 32033 86711 32091 86717
rect 32398 86708 32404 86720
rect 32456 86708 32462 86760
rect 30282 86680 30288 86692
rect 29068 86652 30288 86680
rect 28960 86640 28966 86652
rect 30282 86640 30288 86652
rect 30340 86640 30346 86692
rect 30926 86640 30932 86692
rect 30984 86680 30990 86692
rect 31021 86683 31079 86689
rect 31021 86680 31033 86683
rect 30984 86652 31033 86680
rect 30984 86640 30990 86652
rect 31021 86649 31033 86652
rect 31067 86649 31079 86683
rect 31021 86643 31079 86649
rect 31202 86640 31208 86692
rect 31260 86680 31266 86692
rect 32508 86680 32536 86788
rect 32766 86708 32772 86760
rect 32824 86748 32830 86760
rect 32953 86751 33011 86757
rect 32953 86748 32965 86751
rect 32824 86720 32965 86748
rect 32824 86708 32830 86720
rect 32953 86717 32965 86720
rect 32999 86717 33011 86751
rect 32953 86711 33011 86717
rect 33045 86751 33103 86757
rect 33045 86717 33057 86751
rect 33091 86717 33103 86751
rect 33045 86711 33103 86717
rect 31260 86652 32536 86680
rect 31260 86640 31266 86652
rect 32582 86640 32588 86692
rect 32640 86680 32646 86692
rect 33060 86680 33088 86711
rect 32640 86652 33088 86680
rect 33152 86680 33180 86788
rect 33244 86757 33272 86856
rect 33796 86757 33824 86924
rect 33962 86912 33968 86964
rect 34020 86952 34026 86964
rect 37458 86952 37464 86964
rect 34020 86924 37464 86952
rect 34020 86912 34026 86924
rect 37458 86912 37464 86924
rect 37516 86912 37522 86964
rect 33229 86751 33287 86757
rect 33229 86717 33241 86751
rect 33275 86717 33287 86751
rect 33229 86711 33287 86717
rect 33321 86751 33379 86757
rect 33321 86717 33333 86751
rect 33367 86717 33379 86751
rect 33321 86711 33379 86717
rect 33781 86751 33839 86757
rect 33781 86717 33793 86751
rect 33827 86748 33839 86751
rect 33962 86748 33968 86760
rect 33827 86720 33968 86748
rect 33827 86717 33839 86720
rect 33781 86711 33839 86717
rect 33336 86680 33364 86711
rect 33962 86708 33968 86720
rect 34020 86708 34026 86760
rect 37274 86748 37280 86760
rect 37235 86720 37280 86748
rect 37274 86708 37280 86720
rect 37332 86708 37338 86760
rect 37918 86748 37924 86760
rect 37879 86720 37924 86748
rect 37918 86708 37924 86720
rect 37976 86708 37982 86760
rect 33152 86652 33364 86680
rect 32640 86640 32646 86652
rect 19392 86584 23152 86612
rect 19392 86572 19398 86584
rect 28534 86572 28540 86624
rect 28592 86572 28598 86624
rect 28629 86615 28687 86621
rect 28629 86581 28641 86615
rect 28675 86612 28687 86615
rect 32398 86612 32404 86624
rect 28675 86584 32404 86612
rect 28675 86581 28687 86584
rect 28629 86575 28687 86581
rect 32398 86572 32404 86584
rect 32456 86572 32462 86624
rect 32766 86612 32772 86624
rect 32727 86584 32772 86612
rect 32766 86572 32772 86584
rect 32824 86572 32830 86624
rect 33965 86615 34023 86621
rect 33965 86581 33977 86615
rect 34011 86612 34023 86615
rect 34238 86612 34244 86624
rect 34011 86584 34244 86612
rect 34011 86581 34023 86584
rect 33965 86575 34023 86581
rect 34238 86572 34244 86584
rect 34296 86572 34302 86624
rect 37461 86615 37519 86621
rect 37461 86581 37473 86615
rect 37507 86612 37519 86615
rect 37550 86612 37556 86624
rect 37507 86584 37556 86612
rect 37507 86581 37519 86584
rect 37461 86575 37519 86581
rect 37550 86572 37556 86584
rect 37608 86572 37614 86624
rect 37642 86572 37648 86624
rect 37700 86612 37706 86624
rect 38105 86615 38163 86621
rect 38105 86612 38117 86615
rect 37700 86584 38117 86612
rect 37700 86572 37706 86584
rect 38105 86581 38117 86584
rect 38151 86581 38163 86615
rect 38105 86575 38163 86581
rect 1104 86522 38824 86544
rect 1104 86470 19606 86522
rect 19658 86470 19670 86522
rect 19722 86470 19734 86522
rect 19786 86470 19798 86522
rect 19850 86470 38824 86522
rect 1104 86448 38824 86470
rect 19981 86411 20039 86417
rect 19981 86377 19993 86411
rect 20027 86408 20039 86411
rect 20070 86408 20076 86420
rect 20027 86380 20076 86408
rect 20027 86377 20039 86380
rect 19981 86371 20039 86377
rect 20070 86368 20076 86380
rect 20128 86368 20134 86420
rect 26789 86411 26847 86417
rect 26789 86377 26801 86411
rect 26835 86408 26847 86411
rect 27798 86408 27804 86420
rect 26835 86380 27804 86408
rect 26835 86377 26847 86380
rect 26789 86371 26847 86377
rect 27798 86368 27804 86380
rect 27856 86368 27862 86420
rect 28629 86411 28687 86417
rect 28629 86377 28641 86411
rect 28675 86408 28687 86411
rect 29270 86408 29276 86420
rect 28675 86380 29276 86408
rect 28675 86377 28687 86380
rect 28629 86371 28687 86377
rect 29270 86368 29276 86380
rect 29328 86368 29334 86420
rect 29733 86411 29791 86417
rect 29733 86377 29745 86411
rect 29779 86408 29791 86411
rect 29822 86408 29828 86420
rect 29779 86380 29828 86408
rect 29779 86377 29791 86380
rect 29733 86371 29791 86377
rect 29822 86368 29828 86380
rect 29880 86368 29886 86420
rect 32306 86368 32312 86420
rect 32364 86408 32370 86420
rect 33229 86411 33287 86417
rect 33229 86408 33241 86411
rect 32364 86380 33241 86408
rect 32364 86368 32370 86380
rect 33229 86377 33241 86380
rect 33275 86377 33287 86411
rect 33229 86371 33287 86377
rect 1854 86340 1860 86352
rect 1815 86312 1860 86340
rect 1854 86300 1860 86312
rect 1912 86300 1918 86352
rect 25498 86300 25504 86352
rect 25556 86340 25562 86352
rect 28810 86340 28816 86352
rect 25556 86312 28120 86340
rect 25556 86300 25562 86312
rect 19886 86272 19892 86284
rect 19847 86244 19892 86272
rect 19886 86232 19892 86244
rect 19944 86232 19950 86284
rect 23382 86272 23388 86284
rect 23343 86244 23388 86272
rect 23382 86232 23388 86244
rect 23440 86232 23446 86284
rect 26694 86272 26700 86284
rect 26655 86244 26700 86272
rect 26694 86232 26700 86244
rect 26752 86232 26758 86284
rect 28092 86281 28120 86312
rect 28368 86312 28816 86340
rect 28368 86281 28396 86312
rect 28810 86300 28816 86312
rect 28868 86300 28874 86352
rect 29457 86343 29515 86349
rect 28920 86312 29317 86340
rect 27985 86275 28043 86281
rect 27985 86272 27997 86275
rect 26804 86244 27997 86272
rect 26326 86164 26332 86216
rect 26384 86204 26390 86216
rect 26804 86204 26832 86244
rect 27985 86241 27997 86244
rect 28031 86241 28043 86275
rect 27985 86235 28043 86241
rect 28078 86275 28136 86281
rect 28078 86241 28090 86275
rect 28124 86241 28136 86275
rect 28078 86235 28136 86241
rect 28261 86275 28319 86281
rect 28261 86241 28273 86275
rect 28307 86241 28319 86275
rect 28261 86235 28319 86241
rect 28353 86275 28411 86281
rect 28353 86241 28365 86275
rect 28399 86241 28411 86275
rect 28353 86235 28411 86241
rect 28491 86275 28549 86281
rect 28491 86241 28503 86275
rect 28537 86272 28549 86275
rect 28920 86272 28948 86312
rect 29289 86284 29317 86312
rect 29457 86309 29469 86343
rect 29503 86340 29515 86343
rect 29503 86312 29868 86340
rect 29503 86309 29515 86312
rect 29457 86303 29515 86309
rect 29089 86275 29147 86281
rect 29089 86272 29101 86275
rect 28537 86244 28948 86272
rect 29013 86244 29101 86272
rect 28537 86241 28549 86244
rect 28491 86235 28549 86241
rect 26384 86176 26832 86204
rect 26384 86164 26390 86176
rect 27246 86164 27252 86216
rect 27304 86204 27310 86216
rect 28276 86204 28304 86235
rect 27304 86176 28304 86204
rect 27304 86164 27310 86176
rect 2038 86136 2044 86148
rect 1999 86108 2044 86136
rect 2038 86096 2044 86108
rect 2096 86096 2102 86148
rect 28258 86096 28264 86148
rect 28316 86136 28322 86148
rect 28368 86136 28396 86235
rect 28810 86164 28816 86216
rect 28868 86204 28874 86216
rect 29013 86204 29041 86244
rect 29089 86241 29101 86244
rect 29135 86241 29147 86275
rect 29089 86235 29147 86241
rect 29182 86275 29240 86281
rect 29182 86241 29194 86275
rect 29228 86241 29240 86275
rect 29182 86235 29240 86241
rect 28868 86176 29041 86204
rect 28868 86164 28874 86176
rect 28316 86108 28396 86136
rect 28316 86096 28322 86108
rect 23290 86028 23296 86080
rect 23348 86068 23354 86080
rect 23569 86071 23627 86077
rect 23569 86068 23581 86071
rect 23348 86040 23581 86068
rect 23348 86028 23354 86040
rect 23569 86037 23581 86040
rect 23615 86037 23627 86071
rect 23569 86031 23627 86037
rect 26970 86028 26976 86080
rect 27028 86068 27034 86080
rect 29196 86068 29224 86235
rect 29271 86232 29277 86284
rect 29329 86232 29335 86284
rect 29638 86281 29644 86284
rect 29365 86275 29423 86281
rect 29365 86241 29377 86275
rect 29411 86241 29423 86275
rect 29365 86235 29423 86241
rect 29593 86275 29644 86281
rect 29593 86241 29605 86275
rect 29639 86241 29644 86275
rect 29593 86235 29644 86241
rect 29380 86204 29408 86235
rect 29638 86232 29644 86235
rect 29696 86232 29702 86284
rect 29840 86216 29868 86312
rect 30742 86300 30748 86352
rect 30800 86340 30806 86352
rect 35986 86340 35992 86352
rect 30800 86312 35992 86340
rect 30800 86300 30806 86312
rect 35986 86300 35992 86312
rect 36044 86300 36050 86352
rect 30193 86275 30251 86281
rect 30193 86241 30205 86275
rect 30239 86241 30251 86275
rect 30193 86235 30251 86241
rect 29288 86176 29408 86204
rect 29288 86148 29316 86176
rect 29822 86164 29828 86216
rect 29880 86164 29886 86216
rect 30006 86164 30012 86216
rect 30064 86204 30070 86216
rect 30208 86204 30236 86235
rect 30282 86232 30288 86284
rect 30340 86272 30346 86284
rect 31495 86275 31553 86281
rect 31495 86272 31507 86275
rect 30340 86244 31507 86272
rect 30340 86232 30346 86244
rect 31495 86241 31507 86244
rect 31541 86241 31553 86275
rect 31495 86235 31553 86241
rect 31941 86275 31999 86281
rect 31941 86241 31953 86275
rect 31987 86272 31999 86275
rect 32122 86272 32128 86284
rect 31987 86244 32128 86272
rect 31987 86241 31999 86244
rect 31941 86235 31999 86241
rect 32122 86232 32128 86244
rect 32180 86272 32186 86284
rect 32490 86272 32496 86284
rect 32180 86244 32496 86272
rect 32180 86232 32186 86244
rect 32490 86232 32496 86244
rect 32548 86232 32554 86284
rect 32858 86232 32864 86284
rect 32916 86272 32922 86284
rect 33045 86275 33103 86281
rect 33045 86272 33057 86275
rect 32916 86244 33057 86272
rect 32916 86232 32922 86244
rect 33045 86241 33057 86244
rect 33091 86241 33103 86275
rect 37182 86272 37188 86284
rect 37143 86244 37188 86272
rect 33045 86235 33103 86241
rect 37182 86232 37188 86244
rect 37240 86232 37246 86284
rect 30064 86176 30236 86204
rect 31573 86207 31631 86213
rect 30064 86164 30070 86176
rect 31573 86173 31585 86207
rect 31619 86204 31631 86207
rect 32033 86207 32091 86213
rect 31619 86176 31708 86204
rect 31619 86173 31631 86176
rect 31573 86167 31631 86173
rect 31680 86148 31708 86176
rect 32033 86173 32045 86207
rect 32079 86204 32091 86207
rect 37090 86204 37096 86216
rect 32079 86176 37096 86204
rect 32079 86173 32091 86176
rect 32033 86167 32091 86173
rect 37090 86164 37096 86176
rect 37148 86164 37154 86216
rect 29270 86096 29276 86148
rect 29328 86096 29334 86148
rect 30377 86139 30435 86145
rect 30377 86105 30389 86139
rect 30423 86136 30435 86139
rect 31478 86136 31484 86148
rect 30423 86108 31484 86136
rect 30423 86105 30435 86108
rect 30377 86099 30435 86105
rect 31478 86096 31484 86108
rect 31536 86096 31542 86148
rect 31662 86096 31668 86148
rect 31720 86096 31726 86148
rect 31018 86068 31024 86080
rect 27028 86040 29224 86068
rect 30979 86040 31024 86068
rect 27028 86028 27034 86040
rect 31018 86028 31024 86040
rect 31076 86028 31082 86080
rect 31202 86028 31208 86080
rect 31260 86068 31266 86080
rect 33686 86068 33692 86080
rect 31260 86040 33692 86068
rect 31260 86028 31266 86040
rect 33686 86028 33692 86040
rect 33744 86028 33750 86080
rect 37366 86068 37372 86080
rect 37327 86040 37372 86068
rect 37366 86028 37372 86040
rect 37424 86028 37430 86080
rect 1104 85978 38824 86000
rect 1104 85926 4246 85978
rect 4298 85926 4310 85978
rect 4362 85926 4374 85978
rect 4426 85926 4438 85978
rect 4490 85926 34966 85978
rect 35018 85926 35030 85978
rect 35082 85926 35094 85978
rect 35146 85926 35158 85978
rect 35210 85926 38824 85978
rect 1104 85904 38824 85926
rect 28534 85864 28540 85876
rect 28092 85836 28540 85864
rect 1854 85660 1860 85672
rect 1815 85632 1860 85660
rect 1854 85620 1860 85632
rect 1912 85620 1918 85672
rect 21818 85620 21824 85672
rect 21876 85660 21882 85672
rect 28092 85669 28120 85836
rect 28534 85824 28540 85836
rect 28592 85824 28598 85876
rect 28810 85824 28816 85876
rect 28868 85864 28874 85876
rect 29638 85864 29644 85876
rect 28868 85836 29644 85864
rect 28868 85824 28874 85836
rect 29638 85824 29644 85836
rect 29696 85824 29702 85876
rect 30742 85796 30748 85808
rect 28322 85768 30748 85796
rect 28322 85669 28350 85768
rect 30742 85756 30748 85768
rect 30800 85756 30806 85808
rect 34146 85796 34152 85808
rect 32324 85768 34152 85796
rect 29178 85688 29184 85740
rect 29236 85688 29242 85740
rect 29822 85728 29828 85740
rect 29288 85700 29828 85728
rect 27801 85663 27859 85669
rect 27801 85660 27813 85663
rect 21876 85632 27813 85660
rect 21876 85620 21882 85632
rect 27801 85629 27813 85632
rect 27847 85629 27859 85663
rect 27801 85623 27859 85629
rect 27894 85663 27952 85669
rect 27894 85629 27906 85663
rect 27940 85629 27952 85663
rect 28077 85663 28135 85669
rect 28077 85660 28089 85663
rect 27894 85623 27952 85629
rect 28000 85632 28089 85660
rect 2041 85595 2099 85601
rect 2041 85561 2053 85595
rect 2087 85592 2099 85595
rect 2682 85592 2688 85604
rect 2087 85564 2688 85592
rect 2087 85561 2099 85564
rect 2041 85555 2099 85561
rect 2682 85552 2688 85564
rect 2740 85552 2746 85604
rect 10318 85552 10324 85604
rect 10376 85592 10382 85604
rect 27909 85592 27937 85623
rect 10376 85564 27937 85592
rect 10376 85552 10382 85564
rect 27798 85484 27804 85536
rect 27856 85524 27862 85536
rect 28000 85524 28028 85632
rect 28077 85629 28089 85632
rect 28123 85629 28135 85663
rect 28077 85623 28135 85629
rect 28307 85663 28365 85669
rect 28307 85629 28319 85663
rect 28353 85629 28365 85663
rect 28307 85623 28365 85629
rect 28534 85620 28540 85672
rect 28592 85660 28598 85672
rect 28905 85663 28963 85669
rect 28905 85660 28917 85663
rect 28592 85632 28917 85660
rect 28592 85620 28598 85632
rect 28905 85629 28917 85632
rect 28951 85629 28963 85663
rect 28905 85623 28963 85629
rect 29053 85663 29111 85669
rect 29053 85629 29065 85663
rect 29099 85660 29111 85663
rect 29196 85660 29224 85688
rect 29288 85669 29316 85700
rect 29822 85688 29828 85700
rect 29880 85688 29886 85740
rect 32122 85728 32128 85740
rect 31772 85700 32128 85728
rect 29099 85632 29224 85660
rect 29273 85663 29331 85669
rect 29099 85629 29111 85632
rect 29053 85623 29111 85629
rect 29273 85629 29285 85663
rect 29319 85629 29331 85663
rect 29273 85623 29331 85629
rect 29411 85663 29469 85669
rect 29411 85629 29423 85663
rect 29457 85660 29469 85663
rect 31202 85660 31208 85672
rect 29457 85632 31208 85660
rect 29457 85629 29469 85632
rect 29411 85623 29469 85629
rect 28166 85592 28172 85604
rect 28127 85564 28172 85592
rect 28166 85552 28172 85564
rect 28224 85552 28230 85604
rect 28810 85552 28816 85604
rect 28868 85592 28874 85604
rect 29181 85595 29239 85601
rect 29181 85592 29193 85595
rect 28868 85564 29193 85592
rect 28868 85552 28874 85564
rect 29181 85561 29193 85564
rect 29227 85561 29239 85595
rect 29181 85555 29239 85561
rect 27856 85496 28028 85524
rect 28445 85527 28503 85533
rect 27856 85484 27862 85496
rect 28445 85493 28457 85527
rect 28491 85524 28503 85527
rect 28902 85524 28908 85536
rect 28491 85496 28908 85524
rect 28491 85493 28503 85496
rect 28445 85487 28503 85493
rect 28902 85484 28908 85496
rect 28960 85484 28966 85536
rect 29288 85524 29316 85623
rect 31202 85620 31208 85632
rect 31260 85620 31266 85672
rect 31389 85663 31447 85669
rect 31389 85629 31401 85663
rect 31435 85629 31447 85663
rect 31389 85623 31447 85629
rect 30742 85592 30748 85604
rect 30703 85564 30748 85592
rect 30742 85552 30748 85564
rect 30800 85552 30806 85604
rect 29362 85524 29368 85536
rect 29288 85496 29368 85524
rect 29362 85484 29368 85496
rect 29420 85484 29426 85536
rect 29546 85524 29552 85536
rect 29507 85496 29552 85524
rect 29546 85484 29552 85496
rect 29604 85484 29610 85536
rect 30374 85484 30380 85536
rect 30432 85524 30438 85536
rect 31404 85524 31432 85623
rect 31478 85620 31484 85672
rect 31536 85660 31542 85672
rect 31772 85669 31800 85700
rect 32122 85688 32128 85700
rect 32180 85688 32186 85740
rect 31757 85663 31815 85669
rect 31536 85632 31581 85660
rect 31536 85620 31542 85632
rect 31757 85629 31769 85663
rect 31803 85629 31815 85663
rect 31757 85623 31815 85629
rect 31941 85663 31999 85669
rect 31941 85629 31953 85663
rect 31987 85660 31999 85663
rect 32324 85660 32352 85768
rect 34146 85756 34152 85768
rect 34204 85756 34210 85808
rect 36906 85756 36912 85808
rect 36964 85796 36970 85808
rect 37461 85799 37519 85805
rect 37461 85796 37473 85799
rect 36964 85768 37473 85796
rect 36964 85756 36970 85768
rect 37461 85765 37473 85768
rect 37507 85765 37519 85799
rect 37461 85759 37519 85765
rect 32398 85688 32404 85740
rect 32456 85728 32462 85740
rect 32456 85700 33088 85728
rect 32456 85688 32462 85700
rect 32674 85660 32680 85672
rect 31987 85632 32352 85660
rect 32635 85632 32680 85660
rect 31987 85629 31999 85632
rect 31941 85623 31999 85629
rect 32674 85620 32680 85632
rect 32732 85620 32738 85672
rect 32769 85663 32827 85669
rect 32769 85629 32781 85663
rect 32815 85629 32827 85663
rect 32950 85660 32956 85672
rect 32911 85632 32956 85660
rect 32769 85623 32827 85629
rect 32582 85552 32588 85604
rect 32640 85592 32646 85604
rect 32784 85592 32812 85623
rect 32950 85620 32956 85632
rect 33008 85620 33014 85672
rect 33060 85669 33088 85700
rect 33045 85663 33103 85669
rect 33045 85629 33057 85663
rect 33091 85629 33103 85663
rect 33045 85623 33103 85629
rect 33505 85663 33563 85669
rect 33505 85629 33517 85663
rect 33551 85660 33563 85663
rect 33962 85660 33968 85672
rect 33551 85632 33968 85660
rect 33551 85629 33563 85632
rect 33505 85623 33563 85629
rect 33962 85620 33968 85632
rect 34020 85620 34026 85672
rect 37274 85660 37280 85672
rect 37235 85632 37280 85660
rect 37274 85620 37280 85632
rect 37332 85620 37338 85672
rect 37918 85660 37924 85672
rect 37879 85632 37924 85660
rect 37918 85620 37924 85632
rect 37976 85620 37982 85672
rect 32640 85564 33732 85592
rect 32640 85552 32646 85564
rect 32490 85524 32496 85536
rect 30432 85496 31432 85524
rect 32451 85496 32496 85524
rect 30432 85484 30438 85496
rect 32490 85484 32496 85496
rect 32548 85484 32554 85536
rect 33704 85533 33732 85564
rect 33689 85527 33747 85533
rect 33689 85493 33701 85527
rect 33735 85493 33747 85527
rect 33689 85487 33747 85493
rect 33870 85484 33876 85536
rect 33928 85524 33934 85536
rect 38105 85527 38163 85533
rect 38105 85524 38117 85527
rect 33928 85496 38117 85524
rect 33928 85484 33934 85496
rect 38105 85493 38117 85496
rect 38151 85493 38163 85527
rect 38105 85487 38163 85493
rect 1104 85434 38824 85456
rect 1104 85382 19606 85434
rect 19658 85382 19670 85434
rect 19722 85382 19734 85434
rect 19786 85382 19798 85434
rect 19850 85382 38824 85434
rect 1104 85360 38824 85382
rect 26789 85323 26847 85329
rect 26789 85289 26801 85323
rect 26835 85320 26847 85323
rect 27246 85320 27252 85332
rect 26835 85292 27252 85320
rect 26835 85289 26847 85292
rect 26789 85283 26847 85289
rect 27246 85280 27252 85292
rect 27304 85280 27310 85332
rect 27798 85280 27804 85332
rect 27856 85320 27862 85332
rect 27856 85292 28028 85320
rect 27856 85280 27862 85292
rect 8938 85212 8944 85264
rect 8996 85252 9002 85264
rect 28000 85252 28028 85292
rect 28350 85280 28356 85332
rect 28408 85320 28414 85332
rect 28810 85320 28816 85332
rect 28408 85292 28816 85320
rect 28408 85280 28414 85292
rect 28810 85280 28816 85292
rect 28868 85280 28874 85332
rect 28902 85280 28908 85332
rect 28960 85280 28966 85332
rect 29270 85320 29276 85332
rect 29196 85292 29276 85320
rect 28077 85255 28135 85261
rect 28077 85252 28089 85255
rect 8996 85224 27937 85252
rect 8996 85212 9002 85224
rect 23201 85187 23259 85193
rect 23201 85153 23213 85187
rect 23247 85184 23259 85187
rect 23382 85184 23388 85196
rect 23247 85156 23388 85184
rect 23247 85153 23259 85156
rect 23201 85147 23259 85153
rect 23382 85144 23388 85156
rect 23440 85144 23446 85196
rect 26418 85144 26424 85196
rect 26476 85184 26482 85196
rect 26694 85184 26700 85196
rect 26476 85156 26700 85184
rect 26476 85144 26482 85156
rect 26694 85144 26700 85156
rect 26752 85144 26758 85196
rect 27154 85144 27160 85196
rect 27212 85184 27218 85196
rect 27909 85193 27937 85224
rect 28000 85224 28089 85252
rect 27801 85187 27859 85193
rect 27801 85184 27813 85187
rect 27212 85156 27813 85184
rect 27212 85144 27218 85156
rect 27801 85153 27813 85156
rect 27847 85153 27859 85187
rect 27801 85147 27859 85153
rect 27894 85187 27952 85193
rect 27894 85153 27906 85187
rect 27940 85153 27952 85187
rect 27894 85147 27952 85153
rect 23290 85076 23296 85128
rect 23348 85116 23354 85128
rect 28000 85116 28028 85224
rect 28077 85221 28089 85224
rect 28123 85221 28135 85255
rect 28920 85252 28948 85280
rect 29196 85261 29224 85292
rect 29270 85280 29276 85292
rect 29328 85280 29334 85332
rect 30193 85323 30251 85329
rect 30193 85289 30205 85323
rect 30239 85320 30251 85323
rect 32950 85320 32956 85332
rect 30239 85292 32956 85320
rect 30239 85289 30251 85292
rect 30193 85283 30251 85289
rect 32950 85280 32956 85292
rect 33008 85280 33014 85332
rect 33410 85280 33416 85332
rect 33468 85320 33474 85332
rect 33505 85323 33563 85329
rect 33505 85320 33517 85323
rect 33468 85292 33517 85320
rect 33468 85280 33474 85292
rect 33505 85289 33517 85292
rect 33551 85289 33563 85323
rect 33505 85283 33563 85289
rect 28077 85215 28135 85221
rect 28736 85224 28948 85252
rect 29181 85255 29239 85261
rect 28166 85184 28172 85196
rect 28079 85156 28172 85184
rect 28166 85144 28172 85156
rect 28224 85144 28230 85196
rect 28307 85187 28365 85193
rect 28307 85153 28319 85187
rect 28353 85184 28365 85187
rect 28442 85184 28448 85196
rect 28353 85156 28448 85184
rect 28353 85153 28365 85156
rect 28307 85147 28365 85153
rect 28442 85144 28448 85156
rect 28500 85144 28506 85196
rect 23348 85088 28028 85116
rect 28184 85116 28212 85144
rect 28184 85088 28396 85116
rect 23348 85076 23354 85088
rect 28368 85060 28396 85088
rect 23385 85051 23443 85057
rect 23385 85017 23397 85051
rect 23431 85048 23443 85051
rect 25866 85048 25872 85060
rect 23431 85020 25872 85048
rect 23431 85017 23443 85020
rect 23385 85011 23443 85017
rect 25866 85008 25872 85020
rect 25924 85008 25930 85060
rect 28350 85008 28356 85060
rect 28408 85008 28414 85060
rect 28166 84940 28172 84992
rect 28224 84980 28230 84992
rect 28445 84983 28503 84989
rect 28445 84980 28457 84983
rect 28224 84952 28457 84980
rect 28224 84940 28230 84952
rect 28445 84949 28457 84952
rect 28491 84949 28503 84983
rect 28736 84980 28764 85224
rect 29181 85221 29193 85255
rect 29227 85221 29239 85255
rect 33042 85252 33048 85264
rect 29181 85215 29239 85221
rect 29426 85224 33048 85252
rect 28902 85184 28908 85196
rect 28863 85156 28908 85184
rect 28902 85144 28908 85156
rect 28960 85144 28966 85196
rect 28994 85144 29000 85196
rect 29052 85184 29058 85196
rect 29426 85193 29454 85224
rect 33042 85212 33048 85224
rect 33100 85212 33106 85264
rect 29273 85187 29331 85193
rect 29052 85156 29097 85184
rect 29052 85144 29058 85156
rect 29273 85153 29285 85187
rect 29319 85153 29331 85187
rect 29273 85147 29331 85153
rect 29411 85187 29469 85193
rect 29411 85153 29423 85187
rect 29457 85153 29469 85187
rect 29411 85147 29469 85153
rect 30009 85187 30067 85193
rect 30009 85153 30021 85187
rect 30055 85184 30067 85187
rect 30098 85184 30104 85196
rect 30055 85156 30104 85184
rect 30055 85153 30067 85156
rect 30009 85147 30067 85153
rect 29288 85116 29316 85147
rect 30098 85144 30104 85156
rect 30156 85144 30162 85196
rect 31389 85187 31447 85193
rect 31389 85153 31401 85187
rect 31435 85153 31447 85187
rect 31389 85147 31447 85153
rect 31757 85187 31815 85193
rect 31757 85153 31769 85187
rect 31803 85184 31815 85187
rect 32122 85184 32128 85196
rect 31803 85156 32128 85184
rect 31803 85153 31815 85156
rect 31757 85147 31815 85153
rect 31404 85116 31432 85147
rect 32122 85144 32128 85156
rect 32180 85144 32186 85196
rect 33410 85184 33416 85196
rect 33371 85156 33416 85184
rect 33410 85144 33416 85156
rect 33468 85144 33474 85196
rect 29288 85088 29408 85116
rect 29380 85060 29408 85088
rect 29564 85088 31432 85116
rect 29362 85008 29368 85060
rect 29420 85008 29426 85060
rect 29564 85057 29592 85088
rect 31478 85076 31484 85128
rect 31536 85116 31542 85128
rect 31849 85119 31907 85125
rect 31536 85088 31629 85116
rect 31536 85076 31542 85088
rect 31849 85085 31861 85119
rect 31895 85116 31907 85119
rect 36630 85116 36636 85128
rect 31895 85088 36636 85116
rect 31895 85085 31907 85088
rect 31849 85079 31907 85085
rect 36630 85076 36636 85088
rect 36688 85076 36694 85128
rect 29549 85051 29607 85057
rect 29549 85017 29561 85051
rect 29595 85017 29607 85051
rect 29549 85011 29607 85017
rect 29822 85008 29828 85060
rect 29880 85048 29886 85060
rect 30837 85051 30895 85057
rect 30837 85048 30849 85051
rect 29880 85020 30849 85048
rect 29880 85008 29886 85020
rect 30837 85017 30849 85020
rect 30883 85017 30895 85051
rect 30837 85011 30895 85017
rect 31202 85008 31208 85060
rect 31260 85048 31266 85060
rect 31496 85048 31524 85076
rect 31260 85020 31524 85048
rect 31260 85008 31266 85020
rect 32950 84980 32956 84992
rect 28736 84952 32956 84980
rect 28445 84943 28503 84949
rect 32950 84940 32956 84952
rect 33008 84940 33014 84992
rect 1104 84890 38824 84912
rect 1104 84838 4246 84890
rect 4298 84838 4310 84890
rect 4362 84838 4374 84890
rect 4426 84838 4438 84890
rect 4490 84838 34966 84890
rect 35018 84838 35030 84890
rect 35082 84838 35094 84890
rect 35146 84838 35158 84890
rect 35210 84838 38824 84890
rect 1104 84816 38824 84838
rect 36078 84776 36084 84788
rect 28322 84748 36084 84776
rect 27522 84668 27528 84720
rect 27580 84708 27586 84720
rect 27580 84680 28212 84708
rect 27580 84668 27586 84680
rect 25038 84600 25044 84652
rect 25096 84640 25102 84652
rect 25096 84612 27937 84640
rect 25096 84600 25102 84612
rect 1854 84572 1860 84584
rect 1815 84544 1860 84572
rect 1854 84532 1860 84544
rect 1912 84532 1918 84584
rect 27062 84532 27068 84584
rect 27120 84572 27126 84584
rect 27909 84581 27937 84612
rect 28184 84581 28212 84680
rect 28322 84581 28350 84748
rect 36078 84736 36084 84748
rect 36136 84736 36142 84788
rect 37734 84736 37740 84788
rect 37792 84776 37798 84788
rect 38194 84776 38200 84788
rect 37792 84748 38200 84776
rect 37792 84736 37798 84748
rect 38194 84736 38200 84748
rect 38252 84736 38258 84788
rect 28626 84668 28632 84720
rect 28684 84708 28690 84720
rect 29181 84711 29239 84717
rect 29181 84708 29193 84711
rect 28684 84680 29193 84708
rect 28684 84668 28690 84680
rect 29181 84677 29193 84680
rect 29227 84677 29239 84711
rect 29181 84671 29239 84677
rect 30650 84668 30656 84720
rect 30708 84708 30714 84720
rect 31478 84708 31484 84720
rect 30708 84680 31484 84708
rect 30708 84668 30714 84680
rect 31478 84668 31484 84680
rect 31536 84708 31542 84720
rect 31536 84680 33180 84708
rect 31536 84668 31542 84680
rect 28442 84600 28448 84652
rect 28500 84640 28506 84652
rect 29822 84640 29828 84652
rect 28500 84612 29828 84640
rect 28500 84600 28506 84612
rect 29822 84600 29828 84612
rect 29880 84600 29886 84652
rect 30466 84600 30472 84652
rect 30524 84640 30530 84652
rect 31573 84643 31631 84649
rect 31573 84640 31585 84643
rect 30524 84612 31585 84640
rect 30524 84600 30530 84612
rect 31573 84609 31585 84612
rect 31619 84609 31631 84643
rect 32677 84643 32735 84649
rect 32677 84640 32689 84643
rect 31573 84603 31631 84609
rect 31726 84612 32689 84640
rect 27801 84575 27859 84581
rect 27801 84572 27813 84575
rect 27120 84544 27813 84572
rect 27120 84532 27126 84544
rect 27801 84541 27813 84544
rect 27847 84541 27859 84575
rect 27801 84535 27859 84541
rect 27894 84575 27952 84581
rect 27894 84541 27906 84575
rect 27940 84541 27952 84575
rect 27894 84535 27952 84541
rect 28169 84575 28227 84581
rect 28169 84541 28181 84575
rect 28215 84541 28227 84575
rect 28169 84535 28227 84541
rect 28307 84575 28365 84581
rect 28307 84541 28319 84575
rect 28353 84541 28365 84575
rect 28307 84535 28365 84541
rect 28626 84532 28632 84584
rect 28684 84572 28690 84584
rect 28997 84575 29055 84581
rect 28997 84572 29009 84575
rect 28684 84544 29009 84572
rect 28684 84532 28690 84544
rect 28997 84541 29009 84544
rect 29043 84541 29055 84575
rect 28997 84535 29055 84541
rect 29638 84532 29644 84584
rect 29696 84572 29702 84584
rect 31113 84575 31171 84581
rect 31113 84572 31125 84575
rect 29696 84544 31125 84572
rect 29696 84532 29702 84544
rect 31113 84541 31125 84544
rect 31159 84541 31171 84575
rect 31113 84535 31171 84541
rect 31202 84532 31208 84584
rect 31260 84572 31266 84584
rect 31478 84572 31484 84584
rect 31260 84544 31305 84572
rect 31439 84544 31484 84572
rect 31260 84532 31266 84544
rect 31478 84532 31484 84544
rect 31536 84532 31542 84584
rect 2041 84507 2099 84513
rect 2041 84473 2053 84507
rect 2087 84504 2099 84507
rect 2590 84504 2596 84516
rect 2087 84476 2596 84504
rect 2087 84473 2099 84476
rect 2041 84467 2099 84473
rect 2590 84464 2596 84476
rect 2648 84464 2654 84516
rect 28077 84507 28135 84513
rect 28077 84473 28089 84507
rect 28123 84504 28135 84507
rect 29270 84504 29276 84516
rect 28123 84476 29276 84504
rect 28123 84473 28135 84476
rect 28077 84467 28135 84473
rect 29270 84464 29276 84476
rect 29328 84464 29334 84516
rect 29822 84464 29828 84516
rect 29880 84504 29886 84516
rect 29880 84476 30420 84504
rect 29880 84464 29886 84476
rect 28445 84439 28503 84445
rect 28445 84405 28457 84439
rect 28491 84436 28503 84439
rect 28994 84436 29000 84448
rect 28491 84408 29000 84436
rect 28491 84405 28503 84408
rect 28445 84399 28503 84405
rect 28994 84396 29000 84408
rect 29052 84396 29058 84448
rect 30392 84436 30420 84476
rect 30466 84464 30472 84516
rect 30524 84504 30530 84516
rect 31220 84504 31248 84532
rect 31726 84504 31754 84612
rect 32677 84609 32689 84612
rect 32723 84609 32735 84643
rect 32677 84603 32735 84609
rect 33152 84581 33180 84680
rect 33962 84668 33968 84720
rect 34020 84708 34026 84720
rect 38105 84711 38163 84717
rect 38105 84708 38117 84711
rect 34020 84680 38117 84708
rect 34020 84668 34026 84680
rect 38105 84677 38117 84680
rect 38151 84677 38163 84711
rect 38105 84671 38163 84677
rect 32769 84575 32827 84581
rect 32769 84541 32781 84575
rect 32815 84541 32827 84575
rect 32769 84535 32827 84541
rect 33137 84575 33195 84581
rect 33137 84541 33149 84575
rect 33183 84541 33195 84575
rect 33137 84535 33195 84541
rect 33321 84575 33379 84581
rect 33321 84541 33333 84575
rect 33367 84572 33379 84575
rect 36722 84572 36728 84584
rect 33367 84544 36728 84572
rect 33367 84541 33379 84544
rect 33321 84535 33379 84541
rect 30524 84476 30569 84504
rect 31220 84476 31754 84504
rect 32125 84507 32183 84513
rect 30524 84464 30530 84476
rect 32125 84473 32137 84507
rect 32171 84504 32183 84507
rect 32306 84504 32312 84516
rect 32171 84476 32312 84504
rect 32171 84473 32183 84476
rect 32125 84467 32183 84473
rect 32306 84464 32312 84476
rect 32364 84464 32370 84516
rect 32784 84436 32812 84535
rect 36722 84532 36728 84544
rect 36780 84532 36786 84584
rect 37274 84572 37280 84584
rect 37235 84544 37280 84572
rect 37274 84532 37280 84544
rect 37332 84532 37338 84584
rect 37918 84572 37924 84584
rect 37879 84544 37924 84572
rect 37918 84532 37924 84544
rect 37976 84532 37982 84584
rect 34238 84464 34244 84516
rect 34296 84504 34302 84516
rect 38654 84504 38660 84516
rect 34296 84476 38660 84504
rect 34296 84464 34302 84476
rect 38654 84464 38660 84476
rect 38712 84464 38718 84516
rect 30392 84408 32812 84436
rect 37461 84439 37519 84445
rect 37461 84405 37473 84439
rect 37507 84436 37519 84439
rect 37734 84436 37740 84448
rect 37507 84408 37740 84436
rect 37507 84405 37519 84408
rect 37461 84399 37519 84405
rect 37734 84396 37740 84408
rect 37792 84396 37798 84448
rect 1104 84346 38824 84368
rect 1104 84294 19606 84346
rect 19658 84294 19670 84346
rect 19722 84294 19734 84346
rect 19786 84294 19798 84346
rect 19850 84294 38824 84346
rect 1104 84272 38824 84294
rect 28445 84235 28503 84241
rect 28445 84201 28457 84235
rect 28491 84232 28503 84235
rect 28491 84204 30328 84232
rect 28491 84201 28503 84204
rect 28445 84195 28503 84201
rect 9214 84124 9220 84176
rect 9272 84164 9278 84176
rect 28077 84167 28135 84173
rect 9272 84136 27937 84164
rect 9272 84124 9278 84136
rect 1854 84096 1860 84108
rect 1815 84068 1860 84096
rect 1854 84056 1860 84068
rect 1912 84056 1918 84108
rect 27798 84096 27804 84108
rect 27759 84068 27804 84096
rect 27798 84056 27804 84068
rect 27856 84056 27862 84108
rect 27909 84105 27937 84136
rect 28077 84133 28089 84167
rect 28123 84164 28135 84167
rect 28718 84164 28724 84176
rect 28123 84136 28724 84164
rect 28123 84133 28135 84136
rect 28077 84127 28135 84133
rect 28718 84124 28724 84136
rect 28776 84124 28782 84176
rect 29086 84124 29092 84176
rect 29144 84164 29150 84176
rect 29362 84164 29368 84176
rect 29144 84136 29368 84164
rect 29144 84124 29150 84136
rect 29362 84124 29368 84136
rect 29420 84124 29426 84176
rect 27894 84099 27952 84105
rect 27894 84065 27906 84099
rect 27940 84065 27952 84099
rect 27894 84059 27952 84065
rect 28169 84099 28227 84105
rect 28169 84065 28181 84099
rect 28215 84065 28227 84099
rect 28169 84059 28227 84065
rect 28266 84099 28324 84105
rect 28266 84065 28278 84099
rect 28312 84065 28324 84099
rect 28266 84059 28324 84065
rect 2041 83963 2099 83969
rect 2041 83929 2053 83963
rect 2087 83960 2099 83963
rect 4062 83960 4068 83972
rect 2087 83932 4068 83960
rect 2087 83929 2099 83932
rect 2041 83923 2099 83929
rect 4062 83920 4068 83932
rect 4120 83920 4126 83972
rect 28184 83892 28212 84059
rect 28283 83960 28311 84059
rect 28442 84056 28448 84108
rect 28500 84096 28506 84108
rect 28626 84096 28632 84108
rect 28500 84068 28632 84096
rect 28500 84056 28506 84068
rect 28626 84056 28632 84068
rect 28684 84096 28690 84108
rect 28905 84099 28963 84105
rect 28905 84096 28917 84099
rect 28684 84068 28917 84096
rect 28684 84056 28690 84068
rect 28905 84065 28917 84068
rect 28951 84065 28963 84099
rect 28905 84059 28963 84065
rect 29013 84068 29224 84096
rect 29013 83960 29041 84068
rect 29086 83988 29092 84040
rect 29144 83988 29150 84040
rect 28283 83932 29041 83960
rect 28994 83892 29000 83904
rect 28184 83864 29000 83892
rect 28994 83852 29000 83864
rect 29052 83852 29058 83904
rect 29104 83901 29132 83988
rect 29196 83960 29224 84068
rect 29270 84056 29276 84108
rect 29328 84096 29334 84108
rect 29641 84099 29699 84105
rect 29641 84096 29653 84099
rect 29328 84068 29653 84096
rect 29328 84056 29334 84068
rect 29641 84065 29653 84068
rect 29687 84096 29699 84099
rect 30006 84096 30012 84108
rect 29687 84068 30012 84096
rect 29687 84065 29699 84068
rect 29641 84059 29699 84065
rect 30006 84056 30012 84068
rect 30064 84056 30070 84108
rect 30300 84096 30328 84204
rect 30374 84192 30380 84244
rect 30432 84232 30438 84244
rect 31662 84232 31668 84244
rect 30432 84204 31668 84232
rect 30432 84192 30438 84204
rect 31662 84192 31668 84204
rect 31720 84192 31726 84244
rect 31021 84099 31079 84105
rect 31021 84096 31033 84099
rect 30300 84068 31033 84096
rect 31021 84065 31033 84068
rect 31067 84065 31079 84099
rect 31021 84059 31079 84065
rect 31389 84099 31447 84105
rect 31389 84065 31401 84099
rect 31435 84096 31447 84099
rect 31478 84096 31484 84108
rect 31435 84068 31484 84096
rect 31435 84065 31447 84068
rect 31389 84059 31447 84065
rect 31478 84056 31484 84068
rect 31536 84056 31542 84108
rect 31573 84099 31631 84105
rect 31573 84065 31585 84099
rect 31619 84096 31631 84099
rect 36538 84096 36544 84108
rect 31619 84068 36544 84096
rect 31619 84065 31631 84068
rect 31573 84059 31631 84065
rect 36538 84056 36544 84068
rect 36596 84056 36602 84108
rect 37182 84096 37188 84108
rect 37143 84068 37188 84096
rect 37182 84056 37188 84068
rect 37240 84056 37246 84108
rect 30650 83988 30656 84040
rect 30708 84028 30714 84040
rect 30929 84031 30987 84037
rect 30929 84028 30941 84031
rect 30708 84000 30941 84028
rect 30708 83988 30714 84000
rect 30929 83997 30941 84000
rect 30975 84028 30987 84031
rect 31202 84028 31208 84040
rect 30975 84000 31208 84028
rect 30975 83997 30987 84000
rect 30929 83991 30987 83997
rect 31202 83988 31208 84000
rect 31260 83988 31266 84040
rect 33686 83988 33692 84040
rect 33744 84028 33750 84040
rect 36354 84028 36360 84040
rect 33744 84000 36360 84028
rect 33744 83988 33750 84000
rect 36354 83988 36360 84000
rect 36412 83988 36418 84040
rect 35894 83960 35900 83972
rect 29196 83932 35900 83960
rect 35894 83920 35900 83932
rect 35952 83920 35958 83972
rect 29089 83895 29147 83901
rect 29089 83861 29101 83895
rect 29135 83861 29147 83895
rect 29089 83855 29147 83861
rect 29825 83895 29883 83901
rect 29825 83861 29837 83895
rect 29871 83892 29883 83895
rect 30374 83892 30380 83904
rect 29871 83864 30380 83892
rect 29871 83861 29883 83864
rect 29825 83855 29883 83861
rect 30374 83852 30380 83864
rect 30432 83852 30438 83904
rect 30469 83895 30527 83901
rect 30469 83861 30481 83895
rect 30515 83892 30527 83895
rect 31478 83892 31484 83904
rect 30515 83864 31484 83892
rect 30515 83861 30527 83864
rect 30469 83855 30527 83861
rect 31478 83852 31484 83864
rect 31536 83852 31542 83904
rect 36354 83852 36360 83904
rect 36412 83892 36418 83904
rect 37369 83895 37427 83901
rect 37369 83892 37381 83895
rect 36412 83864 37381 83892
rect 36412 83852 36418 83864
rect 37369 83861 37381 83864
rect 37415 83861 37427 83895
rect 37369 83855 37427 83861
rect 1104 83802 38824 83824
rect 1104 83750 4246 83802
rect 4298 83750 4310 83802
rect 4362 83750 4374 83802
rect 4426 83750 4438 83802
rect 4490 83750 34966 83802
rect 35018 83750 35030 83802
rect 35082 83750 35094 83802
rect 35146 83750 35158 83802
rect 35210 83750 38824 83802
rect 1104 83728 38824 83750
rect 25130 83648 25136 83700
rect 25188 83688 25194 83700
rect 30466 83688 30472 83700
rect 25188 83660 27752 83688
rect 25188 83648 25194 83660
rect 3418 83580 3424 83632
rect 3476 83620 3482 83632
rect 27724 83620 27752 83660
rect 29380 83660 30472 83688
rect 29380 83620 29408 83660
rect 30466 83648 30472 83660
rect 30524 83648 30530 83700
rect 30561 83691 30619 83697
rect 30561 83657 30573 83691
rect 30607 83688 30619 83691
rect 31662 83688 31668 83700
rect 30607 83660 31668 83688
rect 30607 83657 30619 83660
rect 30561 83651 30619 83657
rect 31662 83648 31668 83660
rect 31720 83648 31726 83700
rect 3476 83592 27660 83620
rect 27724 83592 29408 83620
rect 29457 83623 29515 83629
rect 3476 83580 3482 83592
rect 26878 83444 26884 83496
rect 26936 83484 26942 83496
rect 27632 83493 27660 83592
rect 29457 83589 29469 83623
rect 29503 83620 29515 83623
rect 30650 83620 30656 83632
rect 29503 83592 30656 83620
rect 29503 83589 29515 83592
rect 29457 83583 29515 83589
rect 30650 83580 30656 83592
rect 30708 83580 30714 83632
rect 31202 83580 31208 83632
rect 31260 83580 31266 83632
rect 28166 83552 28172 83564
rect 27816 83524 28172 83552
rect 27816 83493 27844 83524
rect 28166 83512 28172 83524
rect 28224 83552 28230 83564
rect 28718 83552 28724 83564
rect 28224 83524 28724 83552
rect 28224 83512 28230 83524
rect 28718 83512 28724 83524
rect 28776 83512 28782 83564
rect 28994 83512 29000 83564
rect 29052 83552 29058 83564
rect 31220 83552 31248 83580
rect 29052 83524 31156 83552
rect 31220 83524 31524 83552
rect 29052 83512 29058 83524
rect 27525 83487 27583 83493
rect 27525 83484 27537 83487
rect 26936 83456 27537 83484
rect 26936 83444 26942 83456
rect 27525 83453 27537 83456
rect 27571 83453 27583 83487
rect 27525 83447 27583 83453
rect 27618 83487 27676 83493
rect 27618 83453 27630 83487
rect 27664 83453 27676 83487
rect 27618 83447 27676 83453
rect 27801 83487 27859 83493
rect 27801 83453 27813 83487
rect 27847 83453 27859 83487
rect 27801 83447 27859 83453
rect 28031 83487 28089 83493
rect 28031 83453 28043 83487
rect 28077 83484 28089 83487
rect 28077 83456 29224 83484
rect 28077 83453 28089 83456
rect 28031 83447 28089 83453
rect 27893 83419 27951 83425
rect 27893 83385 27905 83419
rect 27939 83416 27951 83419
rect 29086 83416 29092 83428
rect 27939 83388 29092 83416
rect 27939 83385 27951 83388
rect 27893 83379 27951 83385
rect 29086 83376 29092 83388
rect 29144 83376 29150 83428
rect 28169 83351 28227 83357
rect 28169 83317 28181 83351
rect 28215 83348 28227 83351
rect 28626 83348 28632 83360
rect 28215 83320 28632 83348
rect 28215 83317 28227 83320
rect 28169 83311 28227 83317
rect 28626 83308 28632 83320
rect 28684 83308 28690 83360
rect 29196 83348 29224 83456
rect 29270 83444 29276 83496
rect 29328 83484 29334 83496
rect 31128 83493 31156 83524
rect 31113 83487 31171 83493
rect 29328 83456 29373 83484
rect 29328 83444 29334 83456
rect 31113 83453 31125 83487
rect 31159 83453 31171 83487
rect 31113 83447 31171 83453
rect 31202 83444 31208 83496
rect 31260 83484 31266 83496
rect 31496 83493 31524 83524
rect 31481 83487 31539 83493
rect 31260 83456 31305 83484
rect 31260 83444 31266 83456
rect 31481 83453 31493 83487
rect 31527 83453 31539 83487
rect 31481 83447 31539 83453
rect 31665 83487 31723 83493
rect 31665 83453 31677 83487
rect 31711 83484 31723 83487
rect 34238 83484 34244 83496
rect 31711 83456 34244 83484
rect 31711 83453 31723 83456
rect 31665 83447 31723 83453
rect 34238 83444 34244 83456
rect 34296 83444 34302 83496
rect 37274 83484 37280 83496
rect 37235 83456 37280 83484
rect 37274 83444 37280 83456
rect 37332 83444 37338 83496
rect 37918 83484 37924 83496
rect 37879 83456 37924 83484
rect 37918 83444 37924 83456
rect 37976 83444 37982 83496
rect 30098 83376 30104 83428
rect 30156 83416 30162 83428
rect 37642 83416 37648 83428
rect 30156 83388 37648 83416
rect 30156 83376 30162 83388
rect 37642 83376 37648 83388
rect 37700 83376 37706 83428
rect 35802 83348 35808 83360
rect 29196 83320 35808 83348
rect 35802 83308 35808 83320
rect 35860 83308 35866 83360
rect 37458 83348 37464 83360
rect 37419 83320 37464 83348
rect 37458 83308 37464 83320
rect 37516 83308 37522 83360
rect 38102 83348 38108 83360
rect 38063 83320 38108 83348
rect 38102 83308 38108 83320
rect 38160 83308 38166 83360
rect 1104 83258 38824 83280
rect 1104 83206 19606 83258
rect 19658 83206 19670 83258
rect 19722 83206 19734 83258
rect 19786 83206 19798 83258
rect 19850 83206 38824 83258
rect 1104 83184 38824 83206
rect 27246 83104 27252 83156
rect 27304 83144 27310 83156
rect 28166 83144 28172 83156
rect 27304 83116 28172 83144
rect 27304 83104 27310 83116
rect 3510 83036 3516 83088
rect 3568 83076 3574 83088
rect 28092 83085 28120 83116
rect 28166 83104 28172 83116
rect 28224 83104 28230 83156
rect 36170 83144 36176 83156
rect 28283 83116 36176 83144
rect 28077 83079 28135 83085
rect 3568 83048 27937 83076
rect 3568 83036 3574 83048
rect 1394 83008 1400 83020
rect 1355 82980 1400 83008
rect 1394 82968 1400 82980
rect 1452 82968 1458 83020
rect 26970 82968 26976 83020
rect 27028 83008 27034 83020
rect 27909 83017 27937 83048
rect 28077 83045 28089 83079
rect 28123 83045 28135 83079
rect 28077 83039 28135 83045
rect 28283 83017 28311 83116
rect 36170 83104 36176 83116
rect 36228 83104 36234 83156
rect 30374 83036 30380 83088
rect 30432 83076 30438 83088
rect 30432 83048 31064 83076
rect 30432 83036 30438 83048
rect 27801 83011 27859 83017
rect 27801 83008 27813 83011
rect 27028 82980 27813 83008
rect 27028 82968 27034 82980
rect 27801 82977 27813 82980
rect 27847 82977 27859 83011
rect 27801 82971 27859 82977
rect 27894 83011 27952 83017
rect 27894 82977 27906 83011
rect 27940 82977 27952 83011
rect 27894 82971 27952 82977
rect 28169 83011 28227 83017
rect 28169 82977 28181 83011
rect 28215 82977 28227 83011
rect 28169 82971 28227 82977
rect 28266 83011 28324 83017
rect 28266 82977 28278 83011
rect 28312 82977 28324 83011
rect 30650 83008 30656 83020
rect 30611 82980 30656 83008
rect 28266 82971 28324 82977
rect 1673 82943 1731 82949
rect 1673 82909 1685 82943
rect 1719 82940 1731 82943
rect 8846 82940 8852 82952
rect 1719 82912 8852 82940
rect 1719 82909 1731 82912
rect 1673 82903 1731 82909
rect 8846 82900 8852 82912
rect 8904 82900 8910 82952
rect 28184 82804 28212 82971
rect 30650 82968 30656 82980
rect 30708 82968 30714 83020
rect 31036 83017 31064 83048
rect 31021 83011 31079 83017
rect 31021 82977 31033 83011
rect 31067 82977 31079 83011
rect 31021 82971 31079 82977
rect 31110 82968 31116 83020
rect 31168 83008 31174 83020
rect 31168 82980 31213 83008
rect 31168 82968 31174 82980
rect 30009 82943 30067 82949
rect 30009 82940 30021 82943
rect 28276 82912 30021 82940
rect 28276 82884 28304 82912
rect 30009 82909 30021 82912
rect 30055 82909 30067 82943
rect 30009 82903 30067 82909
rect 30745 82943 30803 82949
rect 30745 82909 30757 82943
rect 30791 82940 30803 82943
rect 31202 82940 31208 82952
rect 30791 82912 31208 82940
rect 30791 82909 30803 82912
rect 30745 82903 30803 82909
rect 31202 82900 31208 82912
rect 31260 82900 31266 82952
rect 28258 82832 28264 82884
rect 28316 82832 28322 82884
rect 28445 82875 28503 82881
rect 28445 82841 28457 82875
rect 28491 82872 28503 82875
rect 29822 82872 29828 82884
rect 28491 82844 29828 82872
rect 28491 82841 28503 82844
rect 28445 82835 28503 82841
rect 29822 82832 29828 82844
rect 29880 82832 29886 82884
rect 29086 82804 29092 82816
rect 28184 82776 29092 82804
rect 29086 82764 29092 82776
rect 29144 82764 29150 82816
rect 1104 82714 38824 82736
rect 1104 82662 4246 82714
rect 4298 82662 4310 82714
rect 4362 82662 4374 82714
rect 4426 82662 4438 82714
rect 4490 82662 34966 82714
rect 35018 82662 35030 82714
rect 35082 82662 35094 82714
rect 35146 82662 35158 82714
rect 35210 82662 38824 82714
rect 1104 82640 38824 82662
rect 27985 82603 28043 82609
rect 27985 82569 27997 82603
rect 28031 82600 28043 82603
rect 28994 82600 29000 82612
rect 28031 82572 29000 82600
rect 28031 82569 28043 82572
rect 27985 82563 28043 82569
rect 28994 82560 29000 82572
rect 29052 82560 29058 82612
rect 29089 82603 29147 82609
rect 29089 82569 29101 82603
rect 29135 82600 29147 82603
rect 30650 82600 30656 82612
rect 29135 82572 30656 82600
rect 29135 82569 29147 82572
rect 29089 82563 29147 82569
rect 30650 82560 30656 82572
rect 30708 82560 30714 82612
rect 2038 82492 2044 82544
rect 2096 82532 2102 82544
rect 2096 82504 28580 82532
rect 2096 82492 2102 82504
rect 1946 82424 1952 82476
rect 2004 82464 2010 82476
rect 2004 82436 27476 82464
rect 2004 82424 2010 82436
rect 26694 82356 26700 82408
rect 26752 82396 26758 82408
rect 27448 82405 27476 82436
rect 27522 82424 27528 82476
rect 27580 82464 27586 82476
rect 27580 82436 28488 82464
rect 27580 82424 27586 82436
rect 27341 82399 27399 82405
rect 27341 82396 27353 82399
rect 26752 82368 27353 82396
rect 26752 82356 26758 82368
rect 27341 82365 27353 82368
rect 27387 82365 27399 82399
rect 27341 82359 27399 82365
rect 27434 82399 27492 82405
rect 27434 82365 27446 82399
rect 27480 82365 27492 82399
rect 27434 82359 27492 82365
rect 27847 82399 27905 82405
rect 27847 82365 27859 82399
rect 27893 82396 27905 82399
rect 28166 82396 28172 82408
rect 27893 82368 28172 82396
rect 27893 82365 27905 82368
rect 27847 82359 27905 82365
rect 28166 82356 28172 82368
rect 28224 82356 28230 82408
rect 28460 82405 28488 82436
rect 28552 82405 28580 82504
rect 29822 82492 29828 82544
rect 29880 82532 29886 82544
rect 30282 82532 30288 82544
rect 29880 82504 30288 82532
rect 29880 82492 29886 82504
rect 30282 82492 30288 82504
rect 30340 82492 30346 82544
rect 37366 82532 37372 82544
rect 30392 82504 37372 82532
rect 28445 82399 28503 82405
rect 28445 82365 28457 82399
rect 28491 82365 28503 82399
rect 28445 82359 28503 82365
rect 28538 82399 28596 82405
rect 28538 82365 28550 82399
rect 28584 82365 28596 82399
rect 28718 82396 28724 82408
rect 28679 82368 28724 82396
rect 28538 82359 28596 82365
rect 28718 82356 28724 82368
rect 28776 82356 28782 82408
rect 28951 82399 29009 82405
rect 28951 82365 28963 82399
rect 28997 82396 29009 82399
rect 30392 82396 30420 82504
rect 37366 82492 37372 82504
rect 37424 82492 37430 82544
rect 37461 82535 37519 82541
rect 37461 82501 37473 82535
rect 37507 82532 37519 82535
rect 39206 82532 39212 82544
rect 37507 82504 39212 82532
rect 37507 82501 37519 82504
rect 37461 82495 37519 82501
rect 39206 82492 39212 82504
rect 39264 82492 39270 82544
rect 31570 82464 31576 82476
rect 31531 82436 31576 82464
rect 31570 82424 31576 82436
rect 31628 82424 31634 82476
rect 31110 82396 31116 82408
rect 28997 82368 30420 82396
rect 31071 82368 31116 82396
rect 28997 82365 29009 82368
rect 28951 82359 29009 82365
rect 31110 82356 31116 82368
rect 31168 82356 31174 82408
rect 31202 82356 31208 82408
rect 31260 82396 31266 82408
rect 31481 82399 31539 82405
rect 31260 82368 31305 82396
rect 31260 82356 31266 82368
rect 31481 82365 31493 82399
rect 31527 82396 31539 82399
rect 34146 82396 34152 82408
rect 31527 82368 34152 82396
rect 31527 82365 31539 82368
rect 31481 82359 31539 82365
rect 31588 82340 31616 82368
rect 34146 82356 34152 82368
rect 34204 82356 34210 82408
rect 37274 82396 37280 82408
rect 37235 82368 37280 82396
rect 37274 82356 37280 82368
rect 37332 82356 37338 82408
rect 37918 82396 37924 82408
rect 37879 82368 37924 82396
rect 37918 82356 37924 82368
rect 37976 82356 37982 82408
rect 1854 82328 1860 82340
rect 1815 82300 1860 82328
rect 1854 82288 1860 82300
rect 1912 82288 1918 82340
rect 27246 82288 27252 82340
rect 27304 82328 27310 82340
rect 27617 82331 27675 82337
rect 27617 82328 27629 82331
rect 27304 82300 27629 82328
rect 27304 82288 27310 82300
rect 27617 82297 27629 82300
rect 27663 82297 27675 82331
rect 27617 82291 27675 82297
rect 27709 82331 27767 82337
rect 27709 82297 27721 82331
rect 27755 82328 27767 82331
rect 28813 82331 28871 82337
rect 28813 82328 28825 82331
rect 27755 82300 28825 82328
rect 27755 82297 27767 82300
rect 27709 82291 27767 82297
rect 28813 82297 28825 82300
rect 28859 82328 28871 82331
rect 29086 82328 29092 82340
rect 28859 82300 29092 82328
rect 28859 82297 28871 82300
rect 28813 82291 28871 82297
rect 29086 82288 29092 82300
rect 29144 82328 29150 82340
rect 30006 82328 30012 82340
rect 29144 82300 30012 82328
rect 29144 82288 29150 82300
rect 30006 82288 30012 82300
rect 30064 82288 30070 82340
rect 30466 82328 30472 82340
rect 30427 82300 30472 82328
rect 30466 82288 30472 82300
rect 30524 82288 30530 82340
rect 31570 82288 31576 82340
rect 31628 82288 31634 82340
rect 37550 82328 37556 82340
rect 31726 82300 37556 82328
rect 1949 82263 2007 82269
rect 1949 82229 1961 82263
rect 1995 82260 2007 82263
rect 22094 82260 22100 82272
rect 1995 82232 22100 82260
rect 1995 82229 2007 82232
rect 1949 82223 2007 82229
rect 22094 82220 22100 82232
rect 22152 82220 22158 82272
rect 28718 82220 28724 82272
rect 28776 82260 28782 82272
rect 31726 82260 31754 82300
rect 37550 82288 37556 82300
rect 37608 82288 37614 82340
rect 28776 82232 31754 82260
rect 28776 82220 28782 82232
rect 37274 82220 37280 82272
rect 37332 82260 37338 82272
rect 38105 82263 38163 82269
rect 38105 82260 38117 82263
rect 37332 82232 38117 82260
rect 37332 82220 37338 82232
rect 38105 82229 38117 82232
rect 38151 82229 38163 82263
rect 38105 82223 38163 82229
rect 1104 82170 38824 82192
rect 1104 82118 19606 82170
rect 19658 82118 19670 82170
rect 19722 82118 19734 82170
rect 19786 82118 19798 82170
rect 19850 82118 38824 82170
rect 1104 82096 38824 82118
rect 28626 82016 28632 82068
rect 28684 82056 28690 82068
rect 28684 82028 28994 82056
rect 28684 82016 28690 82028
rect 28718 81920 28724 81932
rect 28679 81892 28724 81920
rect 28718 81880 28724 81892
rect 28776 81880 28782 81932
rect 28626 81852 28632 81864
rect 28587 81824 28632 81852
rect 28626 81812 28632 81824
rect 28684 81812 28690 81864
rect 28966 81852 28994 82028
rect 30282 82016 30288 82068
rect 30340 82056 30346 82068
rect 33870 82056 33876 82068
rect 30340 82028 33876 82056
rect 30340 82016 30346 82028
rect 33870 82016 33876 82028
rect 33928 82016 33934 82068
rect 33042 81988 33048 82000
rect 29104 81960 33048 81988
rect 29104 81929 29132 81960
rect 33042 81948 33048 81960
rect 33100 81948 33106 82000
rect 29089 81923 29147 81929
rect 29089 81889 29101 81923
rect 29135 81889 29147 81923
rect 29089 81883 29147 81889
rect 29178 81880 29184 81932
rect 29236 81920 29242 81932
rect 30377 81923 30435 81929
rect 29236 81892 29281 81920
rect 29236 81880 29242 81892
rect 30377 81889 30389 81923
rect 30423 81920 30435 81923
rect 30650 81920 30656 81932
rect 30423 81892 30656 81920
rect 30423 81889 30435 81892
rect 30377 81883 30435 81889
rect 30650 81880 30656 81892
rect 30708 81880 30714 81932
rect 30745 81923 30803 81929
rect 30745 81889 30757 81923
rect 30791 81920 30803 81923
rect 31570 81920 31576 81932
rect 30791 81892 31576 81920
rect 30791 81889 30803 81892
rect 30745 81883 30803 81889
rect 31570 81880 31576 81892
rect 31628 81880 31634 81932
rect 37182 81920 37188 81932
rect 37143 81892 37188 81920
rect 37182 81880 37188 81892
rect 37240 81880 37246 81932
rect 30469 81855 30527 81861
rect 28966 81824 29960 81852
rect 23842 81744 23848 81796
rect 23900 81784 23906 81796
rect 29825 81787 29883 81793
rect 29825 81784 29837 81787
rect 23900 81756 29837 81784
rect 23900 81744 23906 81756
rect 29825 81753 29837 81756
rect 29871 81753 29883 81787
rect 29825 81747 29883 81753
rect 27246 81676 27252 81728
rect 27304 81716 27310 81728
rect 28169 81719 28227 81725
rect 28169 81716 28181 81719
rect 27304 81688 28181 81716
rect 27304 81676 27310 81688
rect 28169 81685 28181 81688
rect 28215 81685 28227 81719
rect 29932 81716 29960 81824
rect 30469 81821 30481 81855
rect 30515 81821 30527 81855
rect 30469 81815 30527 81821
rect 30837 81855 30895 81861
rect 30837 81821 30849 81855
rect 30883 81852 30895 81855
rect 38378 81852 38384 81864
rect 30883 81824 38384 81852
rect 30883 81821 30895 81824
rect 30837 81815 30895 81821
rect 30484 81784 30512 81815
rect 38378 81812 38384 81824
rect 38436 81812 38442 81864
rect 31202 81784 31208 81796
rect 30484 81756 31208 81784
rect 31202 81744 31208 81756
rect 31260 81744 31266 81796
rect 32858 81716 32864 81728
rect 29932 81688 32864 81716
rect 28169 81679 28227 81685
rect 32858 81676 32864 81688
rect 32916 81676 32922 81728
rect 37369 81719 37427 81725
rect 37369 81685 37381 81719
rect 37415 81716 37427 81719
rect 37550 81716 37556 81728
rect 37415 81688 37556 81716
rect 37415 81685 37427 81688
rect 37369 81679 37427 81685
rect 37550 81676 37556 81688
rect 37608 81676 37614 81728
rect 1104 81626 38824 81648
rect 1104 81574 4246 81626
rect 4298 81574 4310 81626
rect 4362 81574 4374 81626
rect 4426 81574 4438 81626
rect 4490 81574 34966 81626
rect 35018 81574 35030 81626
rect 35082 81574 35094 81626
rect 35146 81574 35158 81626
rect 35210 81574 38824 81626
rect 1104 81552 38824 81574
rect 31570 81472 31576 81524
rect 31628 81472 31634 81524
rect 31588 81444 31616 81472
rect 31496 81416 31616 81444
rect 28166 81336 28172 81388
rect 28224 81376 28230 81388
rect 29178 81376 29184 81388
rect 28224 81348 29184 81376
rect 28224 81336 28230 81348
rect 29178 81336 29184 81348
rect 29236 81336 29242 81388
rect 29454 81376 29460 81388
rect 29415 81348 29460 81376
rect 29454 81336 29460 81348
rect 29512 81336 29518 81388
rect 31496 81376 31524 81416
rect 29564 81348 31524 81376
rect 1854 81308 1860 81320
rect 1815 81280 1860 81308
rect 1854 81268 1860 81280
rect 1912 81268 1918 81320
rect 28994 81308 29000 81320
rect 28955 81280 29000 81308
rect 28994 81268 29000 81280
rect 29052 81268 29058 81320
rect 29089 81311 29147 81317
rect 29089 81277 29101 81311
rect 29135 81308 29147 81311
rect 29365 81311 29423 81317
rect 29135 81280 29316 81308
rect 29135 81277 29147 81280
rect 29089 81271 29147 81277
rect 2038 81240 2044 81252
rect 1999 81212 2044 81240
rect 2038 81200 2044 81212
rect 2096 81200 2102 81252
rect 24578 81200 24584 81252
rect 24636 81240 24642 81252
rect 28353 81243 28411 81249
rect 28353 81240 28365 81243
rect 24636 81212 28365 81240
rect 24636 81200 24642 81212
rect 28353 81209 28365 81212
rect 28399 81209 28411 81243
rect 28353 81203 28411 81209
rect 28626 81200 28632 81252
rect 28684 81240 28690 81252
rect 29288 81240 29316 81280
rect 29365 81277 29377 81311
rect 29411 81308 29423 81311
rect 29564 81308 29592 81348
rect 31110 81308 31116 81320
rect 29411 81280 29592 81308
rect 31071 81280 31116 81308
rect 29411 81277 29423 81280
rect 29365 81271 29423 81277
rect 29472 81252 29500 81280
rect 31110 81268 31116 81280
rect 31168 81268 31174 81320
rect 31202 81268 31208 81320
rect 31260 81308 31266 81320
rect 31496 81317 31524 81348
rect 31573 81379 31631 81385
rect 31573 81345 31585 81379
rect 31619 81376 31631 81379
rect 38194 81376 38200 81388
rect 31619 81348 38200 81376
rect 31619 81345 31631 81348
rect 31573 81339 31631 81345
rect 38194 81336 38200 81348
rect 38252 81336 38258 81388
rect 31481 81311 31539 81317
rect 31260 81280 31353 81308
rect 31260 81268 31266 81280
rect 31481 81277 31493 81311
rect 31527 81277 31539 81311
rect 31481 81271 31539 81277
rect 32398 81268 32404 81320
rect 32456 81308 32462 81320
rect 32769 81311 32827 81317
rect 32769 81308 32781 81311
rect 32456 81280 32781 81308
rect 32456 81268 32462 81280
rect 32769 81277 32781 81280
rect 32815 81277 32827 81311
rect 32769 81271 32827 81277
rect 32861 81311 32919 81317
rect 32861 81277 32873 81311
rect 32907 81277 32919 81311
rect 32861 81271 32919 81277
rect 28684 81212 29316 81240
rect 28684 81200 28690 81212
rect 27338 81132 27344 81184
rect 27396 81172 27402 81184
rect 27522 81172 27528 81184
rect 27396 81144 27528 81172
rect 27396 81132 27402 81144
rect 27522 81132 27528 81144
rect 27580 81132 27586 81184
rect 29288 81172 29316 81212
rect 29454 81200 29460 81252
rect 29512 81200 29518 81252
rect 30374 81200 30380 81252
rect 30432 81240 30438 81252
rect 30469 81243 30527 81249
rect 30469 81240 30481 81243
rect 30432 81212 30481 81240
rect 30432 81200 30438 81212
rect 30469 81209 30481 81212
rect 30515 81209 30527 81243
rect 31220 81240 31248 81268
rect 31570 81240 31576 81252
rect 31220 81212 31576 81240
rect 30469 81203 30527 81209
rect 31570 81200 31576 81212
rect 31628 81200 31634 81252
rect 32125 81243 32183 81249
rect 32125 81209 32137 81243
rect 32171 81240 32183 81243
rect 32674 81240 32680 81252
rect 32171 81212 32680 81240
rect 32171 81209 32183 81212
rect 32125 81203 32183 81209
rect 32674 81200 32680 81212
rect 32732 81200 32738 81252
rect 29638 81172 29644 81184
rect 29288 81144 29644 81172
rect 29638 81132 29644 81144
rect 29696 81172 29702 81184
rect 32876 81172 32904 81271
rect 33042 81268 33048 81320
rect 33100 81308 33106 81320
rect 33137 81311 33195 81317
rect 33137 81308 33149 81311
rect 33100 81280 33149 81308
rect 33100 81268 33106 81280
rect 33137 81277 33149 81280
rect 33183 81277 33195 81311
rect 33137 81271 33195 81277
rect 33321 81311 33379 81317
rect 33321 81277 33333 81311
rect 33367 81308 33379 81311
rect 33502 81308 33508 81320
rect 33367 81280 33508 81308
rect 33367 81277 33379 81280
rect 33321 81271 33379 81277
rect 33502 81268 33508 81280
rect 33560 81268 33566 81320
rect 37274 81308 37280 81320
rect 37235 81280 37280 81308
rect 37274 81268 37280 81280
rect 37332 81268 37338 81320
rect 37918 81308 37924 81320
rect 37879 81280 37924 81308
rect 37918 81268 37924 81280
rect 37976 81268 37982 81320
rect 39390 81240 39396 81252
rect 37476 81212 39396 81240
rect 37476 81181 37504 81212
rect 39390 81200 39396 81212
rect 39448 81200 39454 81252
rect 29696 81144 32904 81172
rect 37461 81175 37519 81181
rect 29696 81132 29702 81144
rect 37461 81141 37473 81175
rect 37507 81141 37519 81175
rect 37461 81135 37519 81141
rect 38105 81175 38163 81181
rect 38105 81141 38117 81175
rect 38151 81172 38163 81175
rect 39298 81172 39304 81184
rect 38151 81144 39304 81172
rect 38151 81141 38163 81144
rect 38105 81135 38163 81141
rect 39298 81132 39304 81144
rect 39356 81132 39362 81184
rect 1104 81082 38824 81104
rect 1104 81030 19606 81082
rect 19658 81030 19670 81082
rect 19722 81030 19734 81082
rect 19786 81030 19798 81082
rect 19850 81030 38824 81082
rect 1104 81008 38824 81030
rect 30098 80968 30104 80980
rect 28322 80940 30104 80968
rect 2682 80860 2688 80912
rect 2740 80900 2746 80912
rect 2740 80872 27937 80900
rect 2740 80860 2746 80872
rect 1394 80832 1400 80844
rect 1355 80804 1400 80832
rect 1394 80792 1400 80804
rect 1452 80792 1458 80844
rect 25774 80792 25780 80844
rect 25832 80832 25838 80844
rect 27909 80841 27937 80872
rect 28322 80841 28350 80940
rect 30098 80928 30104 80940
rect 30156 80928 30162 80980
rect 31202 80928 31208 80980
rect 31260 80928 31266 80980
rect 29454 80860 29460 80912
rect 29512 80900 29518 80912
rect 31220 80900 31248 80928
rect 29512 80872 30604 80900
rect 29512 80860 29518 80872
rect 27801 80835 27859 80841
rect 27801 80832 27813 80835
rect 25832 80804 27813 80832
rect 25832 80792 25838 80804
rect 27801 80801 27813 80804
rect 27847 80801 27859 80835
rect 27801 80795 27859 80801
rect 27894 80835 27952 80841
rect 27894 80801 27906 80835
rect 27940 80801 27952 80835
rect 27894 80795 27952 80801
rect 28077 80835 28135 80841
rect 28077 80801 28089 80835
rect 28123 80801 28135 80835
rect 28077 80795 28135 80801
rect 28169 80835 28227 80841
rect 28169 80801 28181 80835
rect 28215 80801 28227 80835
rect 28169 80795 28227 80801
rect 28307 80835 28365 80841
rect 28307 80801 28319 80835
rect 28353 80801 28365 80835
rect 28307 80795 28365 80801
rect 25866 80724 25872 80776
rect 25924 80764 25930 80776
rect 28092 80764 28120 80795
rect 25924 80736 28120 80764
rect 28184 80764 28212 80795
rect 29178 80792 29184 80844
rect 29236 80832 29242 80844
rect 30576 80841 30604 80872
rect 30760 80872 31248 80900
rect 30760 80841 30788 80872
rect 30193 80835 30251 80841
rect 30193 80832 30205 80835
rect 29236 80804 30205 80832
rect 29236 80792 29242 80804
rect 30193 80801 30205 80804
rect 30239 80801 30251 80835
rect 30193 80795 30251 80801
rect 30561 80835 30619 80841
rect 30561 80801 30573 80835
rect 30607 80801 30619 80835
rect 30561 80795 30619 80801
rect 30745 80835 30803 80841
rect 30745 80801 30757 80835
rect 30791 80801 30803 80835
rect 30745 80795 30803 80801
rect 31202 80792 31208 80844
rect 31260 80832 31266 80844
rect 31297 80835 31355 80841
rect 31297 80832 31309 80835
rect 31260 80804 31309 80832
rect 31260 80792 31266 80804
rect 31297 80801 31309 80804
rect 31343 80801 31355 80835
rect 31297 80795 31355 80801
rect 31481 80835 31539 80841
rect 31481 80801 31493 80835
rect 31527 80801 31539 80835
rect 31481 80795 31539 80801
rect 31573 80835 31631 80841
rect 31573 80801 31585 80835
rect 31619 80801 31631 80835
rect 31573 80795 31631 80801
rect 31757 80835 31815 80841
rect 31757 80801 31769 80835
rect 31803 80801 31815 80835
rect 31757 80795 31815 80801
rect 31844 80835 31902 80841
rect 31844 80801 31856 80835
rect 31890 80832 31902 80835
rect 32858 80832 32864 80844
rect 31890 80804 32864 80832
rect 31890 80801 31902 80804
rect 31844 80795 31902 80801
rect 29454 80764 29460 80776
rect 28184 80736 29460 80764
rect 25924 80724 25930 80736
rect 1581 80631 1639 80637
rect 1581 80597 1593 80631
rect 1627 80628 1639 80631
rect 2682 80628 2688 80640
rect 1627 80600 2688 80628
rect 1627 80597 1639 80600
rect 1581 80591 1639 80597
rect 2682 80588 2688 80600
rect 2740 80588 2746 80640
rect 28092 80628 28120 80736
rect 29454 80724 29460 80736
rect 29512 80724 29518 80776
rect 29638 80724 29644 80776
rect 29696 80764 29702 80776
rect 30098 80764 30104 80776
rect 29696 80736 30104 80764
rect 29696 80724 29702 80736
rect 30098 80724 30104 80736
rect 30156 80724 30162 80776
rect 28445 80699 28503 80705
rect 28445 80665 28457 80699
rect 28491 80696 28503 80699
rect 28491 80668 29776 80696
rect 28491 80665 28503 80668
rect 28445 80659 28503 80665
rect 28626 80628 28632 80640
rect 28092 80600 28632 80628
rect 28626 80588 28632 80600
rect 28684 80588 28690 80640
rect 29638 80628 29644 80640
rect 29599 80600 29644 80628
rect 29638 80588 29644 80600
rect 29696 80588 29702 80640
rect 29748 80628 29776 80668
rect 30650 80628 30656 80640
rect 29748 80600 30656 80628
rect 30650 80588 30656 80600
rect 30708 80588 30714 80640
rect 31496 80628 31524 80795
rect 31588 80696 31616 80795
rect 31772 80764 31800 80795
rect 32858 80792 32864 80804
rect 32916 80792 32922 80844
rect 31938 80764 31944 80776
rect 31772 80736 31944 80764
rect 31938 80724 31944 80736
rect 31996 80724 32002 80776
rect 32582 80696 32588 80708
rect 31588 80668 32588 80696
rect 32582 80656 32588 80668
rect 32640 80656 32646 80708
rect 38010 80628 38016 80640
rect 31496 80600 38016 80628
rect 38010 80588 38016 80600
rect 38068 80588 38074 80640
rect 1104 80538 38824 80560
rect 1104 80486 4246 80538
rect 4298 80486 4310 80538
rect 4362 80486 4374 80538
rect 4426 80486 4438 80538
rect 4490 80486 34966 80538
rect 35018 80486 35030 80538
rect 35082 80486 35094 80538
rect 35146 80486 35158 80538
rect 35210 80486 38824 80538
rect 1104 80464 38824 80486
rect 27801 80427 27859 80433
rect 27801 80393 27813 80427
rect 27847 80424 27859 80427
rect 28166 80424 28172 80436
rect 27847 80396 28172 80424
rect 27847 80393 27859 80396
rect 27801 80387 27859 80393
rect 28166 80384 28172 80396
rect 28224 80384 28230 80436
rect 30837 80427 30895 80433
rect 30837 80424 30849 80427
rect 28460 80396 30849 80424
rect 24118 80316 24124 80368
rect 24176 80356 24182 80368
rect 28258 80356 28264 80368
rect 24176 80328 28264 80356
rect 24176 80316 24182 80328
rect 28258 80316 28264 80328
rect 28316 80316 28322 80368
rect 4062 80248 4068 80300
rect 4120 80288 4126 80300
rect 4120 80260 28396 80288
rect 4120 80248 4126 80260
rect 2590 80180 2596 80232
rect 2648 80220 2654 80232
rect 2648 80192 6914 80220
rect 2648 80180 2654 80192
rect 6886 80152 6914 80192
rect 25682 80180 25688 80232
rect 25740 80220 25746 80232
rect 27157 80223 27215 80229
rect 27157 80220 27169 80223
rect 25740 80192 27169 80220
rect 25740 80180 25746 80192
rect 27157 80189 27169 80192
rect 27203 80189 27215 80223
rect 27157 80183 27215 80189
rect 27250 80223 27308 80229
rect 27250 80189 27262 80223
rect 27296 80189 27308 80223
rect 27250 80183 27308 80189
rect 27663 80223 27721 80229
rect 27663 80189 27675 80223
rect 27709 80189 27721 80223
rect 28258 80220 28264 80232
rect 28219 80192 28264 80220
rect 27663 80183 27721 80189
rect 27264 80152 27292 80183
rect 6886 80124 27292 80152
rect 27433 80155 27491 80161
rect 27433 80121 27445 80155
rect 27479 80121 27491 80155
rect 27433 80115 27491 80121
rect 27525 80155 27583 80161
rect 27525 80121 27537 80155
rect 27571 80121 27583 80155
rect 27678 80152 27706 80183
rect 28258 80180 28264 80192
rect 28316 80180 28322 80232
rect 28368 80229 28396 80260
rect 28354 80223 28412 80229
rect 28354 80189 28366 80223
rect 28400 80189 28412 80223
rect 28354 80183 28412 80189
rect 28460 80152 28488 80396
rect 30837 80393 30849 80396
rect 30883 80393 30895 80427
rect 31938 80424 31944 80436
rect 30837 80387 30895 80393
rect 31220 80396 31944 80424
rect 28905 80359 28963 80365
rect 28905 80325 28917 80359
rect 28951 80356 28963 80359
rect 30929 80359 30987 80365
rect 28951 80328 30880 80356
rect 28951 80325 28963 80328
rect 28905 80319 28963 80325
rect 28626 80288 28632 80300
rect 28552 80260 28632 80288
rect 28552 80229 28580 80260
rect 28626 80248 28632 80260
rect 28684 80288 28690 80300
rect 28994 80288 29000 80300
rect 28684 80260 29000 80288
rect 28684 80248 28690 80260
rect 28994 80248 29000 80260
rect 29052 80248 29058 80300
rect 30852 80288 30880 80328
rect 30929 80325 30941 80359
rect 30975 80356 30987 80359
rect 31220 80356 31248 80396
rect 31386 80356 31392 80368
rect 30975 80328 31248 80356
rect 31312 80328 31392 80356
rect 30975 80325 30987 80328
rect 30929 80319 30987 80325
rect 31110 80288 31116 80300
rect 30852 80260 31116 80288
rect 31110 80248 31116 80260
rect 31168 80248 31174 80300
rect 28537 80223 28595 80229
rect 28537 80189 28549 80223
rect 28583 80189 28595 80223
rect 28537 80183 28595 80189
rect 28767 80223 28825 80229
rect 28767 80189 28779 80223
rect 28813 80220 28825 80223
rect 30282 80220 30288 80232
rect 28813 80192 30288 80220
rect 28813 80189 28825 80192
rect 28767 80183 28825 80189
rect 30282 80180 30288 80192
rect 30340 80180 30346 80232
rect 31312 80229 31340 80328
rect 31386 80316 31392 80328
rect 31444 80316 31450 80368
rect 31297 80223 31355 80229
rect 31297 80189 31309 80223
rect 31343 80189 31355 80223
rect 31297 80183 31355 80189
rect 31389 80223 31447 80229
rect 31389 80189 31401 80223
rect 31435 80189 31447 80223
rect 31496 80220 31524 80396
rect 31938 80384 31944 80396
rect 31996 80384 32002 80436
rect 37461 80359 37519 80365
rect 37461 80325 37473 80359
rect 37507 80356 37519 80359
rect 39022 80356 39028 80368
rect 37507 80328 39028 80356
rect 37507 80325 37519 80328
rect 37461 80319 37519 80325
rect 39022 80316 39028 80328
rect 39080 80316 39086 80368
rect 31573 80223 31631 80229
rect 31573 80220 31585 80223
rect 31496 80192 31585 80220
rect 31389 80183 31447 80189
rect 31573 80189 31585 80192
rect 31619 80189 31631 80223
rect 31573 80183 31631 80189
rect 31665 80223 31723 80229
rect 31665 80189 31677 80223
rect 31711 80220 31723 80223
rect 32950 80220 32956 80232
rect 31711 80192 32956 80220
rect 31711 80189 31723 80192
rect 31665 80183 31723 80189
rect 27678 80124 28488 80152
rect 27525 80115 27583 80121
rect 25866 80044 25872 80096
rect 25924 80084 25930 80096
rect 27448 80084 27476 80115
rect 25924 80056 27476 80084
rect 27540 80084 27568 80115
rect 28626 80112 28632 80164
rect 28684 80152 28690 80164
rect 29454 80152 29460 80164
rect 28684 80124 29460 80152
rect 28684 80112 28690 80124
rect 29454 80112 29460 80124
rect 29512 80112 29518 80164
rect 30837 80155 30895 80161
rect 30837 80121 30849 80155
rect 30883 80152 30895 80155
rect 31404 80152 31432 80183
rect 32950 80180 32956 80192
rect 33008 80180 33014 80232
rect 37274 80220 37280 80232
rect 37235 80192 37280 80220
rect 37274 80180 37280 80192
rect 37332 80180 37338 80232
rect 37918 80220 37924 80232
rect 37879 80192 37924 80220
rect 37918 80180 37924 80192
rect 37976 80180 37982 80232
rect 32582 80152 32588 80164
rect 30883 80124 31248 80152
rect 31404 80124 32588 80152
rect 30883 80121 30895 80124
rect 30837 80115 30895 80121
rect 28166 80084 28172 80096
rect 27540 80056 28172 80084
rect 25924 80044 25930 80056
rect 28166 80044 28172 80056
rect 28224 80044 28230 80096
rect 29270 80044 29276 80096
rect 29328 80084 29334 80096
rect 30929 80087 30987 80093
rect 30929 80084 30941 80087
rect 29328 80056 30941 80084
rect 29328 80044 29334 80056
rect 30929 80053 30941 80056
rect 30975 80053 30987 80087
rect 31110 80084 31116 80096
rect 31071 80056 31116 80084
rect 30929 80047 30987 80053
rect 31110 80044 31116 80056
rect 31168 80044 31174 80096
rect 31220 80084 31248 80124
rect 32582 80112 32588 80124
rect 32640 80112 32646 80164
rect 36906 80152 36912 80164
rect 32692 80124 36912 80152
rect 32692 80084 32720 80124
rect 36906 80112 36912 80124
rect 36964 80112 36970 80164
rect 31220 80056 32720 80084
rect 36722 80044 36728 80096
rect 36780 80084 36786 80096
rect 38105 80087 38163 80093
rect 38105 80084 38117 80087
rect 36780 80056 38117 80084
rect 36780 80044 36786 80056
rect 38105 80053 38117 80056
rect 38151 80053 38163 80087
rect 38105 80047 38163 80053
rect 1104 79994 38824 80016
rect 1104 79942 19606 79994
rect 19658 79942 19670 79994
rect 19722 79942 19734 79994
rect 19786 79942 19798 79994
rect 19850 79942 38824 79994
rect 1104 79920 38824 79942
rect 8846 79840 8852 79892
rect 8904 79880 8910 79892
rect 8904 79852 27936 79880
rect 8904 79840 8910 79852
rect 19306 79784 26372 79812
rect 1394 79744 1400 79756
rect 1355 79716 1400 79744
rect 1394 79704 1400 79716
rect 1452 79704 1458 79756
rect 2038 79636 2044 79688
rect 2096 79676 2102 79688
rect 19306 79676 19334 79784
rect 25590 79704 25596 79756
rect 25648 79744 25654 79756
rect 26344 79753 26372 79784
rect 26418 79772 26424 79824
rect 26476 79812 26482 79824
rect 26513 79815 26571 79821
rect 26513 79812 26525 79815
rect 26476 79784 26525 79812
rect 26476 79772 26482 79784
rect 26513 79781 26525 79784
rect 26559 79781 26571 79815
rect 26513 79775 26571 79781
rect 27908 79753 27936 79852
rect 28092 79852 28350 79880
rect 28092 79821 28120 79852
rect 28077 79815 28135 79821
rect 28077 79781 28089 79815
rect 28123 79781 28135 79815
rect 28077 79775 28135 79781
rect 28166 79772 28172 79824
rect 28224 79812 28230 79824
rect 28322 79812 28350 79852
rect 28626 79840 28632 79892
rect 28684 79880 28690 79892
rect 29178 79880 29184 79892
rect 28684 79852 29184 79880
rect 28684 79840 28690 79852
rect 29178 79840 29184 79852
rect 29236 79840 29242 79892
rect 37734 79880 37740 79892
rect 30024 79852 37740 79880
rect 28994 79812 29000 79824
rect 28224 79784 28269 79812
rect 28322 79784 29000 79812
rect 28224 79772 28230 79784
rect 28994 79772 29000 79784
rect 29052 79772 29058 79824
rect 26237 79747 26295 79753
rect 26237 79744 26249 79747
rect 25648 79716 26249 79744
rect 25648 79704 25654 79716
rect 26237 79713 26249 79716
rect 26283 79713 26295 79747
rect 26237 79707 26295 79713
rect 26330 79747 26388 79753
rect 26330 79713 26342 79747
rect 26376 79713 26388 79747
rect 26605 79747 26663 79753
rect 26605 79744 26617 79747
rect 26330 79707 26388 79713
rect 26528 79716 26617 79744
rect 2096 79648 19334 79676
rect 2096 79636 2102 79648
rect 26050 79636 26056 79688
rect 26108 79676 26114 79688
rect 26528 79676 26556 79716
rect 26605 79713 26617 79716
rect 26651 79713 26663 79747
rect 26605 79707 26663 79713
rect 26702 79747 26760 79753
rect 26702 79713 26714 79747
rect 26748 79713 26760 79747
rect 26702 79707 26760 79713
rect 27801 79747 27859 79753
rect 27801 79713 27813 79747
rect 27847 79713 27859 79747
rect 27908 79747 27979 79753
rect 27908 79716 27933 79747
rect 27801 79707 27859 79713
rect 27921 79713 27933 79716
rect 27967 79713 27979 79747
rect 27921 79707 27979 79713
rect 28307 79747 28365 79753
rect 28307 79713 28319 79747
rect 28353 79744 28365 79747
rect 30024 79744 30052 79852
rect 37734 79840 37740 79852
rect 37792 79840 37798 79892
rect 28353 79716 30052 79744
rect 28353 79713 28365 79716
rect 28307 79707 28365 79713
rect 26717 79676 26745 79707
rect 26108 79648 26556 79676
rect 26628 79648 26745 79676
rect 26108 79636 26114 79648
rect 25498 79568 25504 79620
rect 25556 79608 25562 79620
rect 26628 79608 26656 79648
rect 27816 79608 27844 79707
rect 30098 79704 30104 79756
rect 30156 79744 30162 79756
rect 30193 79747 30251 79753
rect 30193 79744 30205 79747
rect 30156 79716 30205 79744
rect 30156 79704 30162 79716
rect 30193 79713 30205 79716
rect 30239 79713 30251 79747
rect 30193 79707 30251 79713
rect 30561 79747 30619 79753
rect 30561 79713 30573 79747
rect 30607 79744 30619 79747
rect 36814 79744 36820 79756
rect 30607 79716 36820 79744
rect 30607 79713 30619 79716
rect 30561 79707 30619 79713
rect 36814 79704 36820 79716
rect 36872 79704 36878 79756
rect 37182 79744 37188 79756
rect 37143 79716 37188 79744
rect 37182 79704 37188 79716
rect 37240 79704 37246 79756
rect 28994 79636 29000 79688
rect 29052 79676 29058 79688
rect 30285 79679 30343 79685
rect 30285 79676 30297 79679
rect 29052 79648 30297 79676
rect 29052 79636 29058 79648
rect 30285 79645 30297 79648
rect 30331 79645 30343 79679
rect 30285 79639 30343 79645
rect 30653 79679 30711 79685
rect 30653 79645 30665 79679
rect 30699 79676 30711 79679
rect 33042 79676 33048 79688
rect 30699 79648 33048 79676
rect 30699 79645 30711 79648
rect 30653 79639 30711 79645
rect 33042 79636 33048 79648
rect 33100 79636 33106 79688
rect 25556 79580 26656 79608
rect 26712 79580 27844 79608
rect 28445 79611 28503 79617
rect 25556 79568 25562 79580
rect 1578 79540 1584 79552
rect 1539 79512 1584 79540
rect 1578 79500 1584 79512
rect 1636 79500 1642 79552
rect 26050 79500 26056 79552
rect 26108 79540 26114 79552
rect 26712 79540 26740 79580
rect 28445 79577 28457 79611
rect 28491 79608 28503 79611
rect 28626 79608 28632 79620
rect 28491 79580 28632 79608
rect 28491 79577 28503 79580
rect 28445 79571 28503 79577
rect 28626 79568 28632 79580
rect 28684 79568 28690 79620
rect 31386 79568 31392 79620
rect 31444 79608 31450 79620
rect 37369 79611 37427 79617
rect 37369 79608 37381 79611
rect 31444 79580 37381 79608
rect 31444 79568 31450 79580
rect 37369 79577 37381 79580
rect 37415 79577 37427 79611
rect 37369 79571 37427 79577
rect 26108 79512 26740 79540
rect 26881 79543 26939 79549
rect 26108 79500 26114 79512
rect 26881 79509 26893 79543
rect 26927 79540 26939 79543
rect 28166 79540 28172 79552
rect 26927 79512 28172 79540
rect 26927 79509 26939 79512
rect 26881 79503 26939 79509
rect 28166 79500 28172 79512
rect 28224 79500 28230 79552
rect 29641 79543 29699 79549
rect 29641 79509 29653 79543
rect 29687 79540 29699 79543
rect 30374 79540 30380 79552
rect 29687 79512 30380 79540
rect 29687 79509 29699 79512
rect 29641 79503 29699 79509
rect 30374 79500 30380 79512
rect 30432 79500 30438 79552
rect 1104 79450 38824 79472
rect 1104 79398 4246 79450
rect 4298 79398 4310 79450
rect 4362 79398 4374 79450
rect 4426 79398 4438 79450
rect 4490 79398 34966 79450
rect 35018 79398 35030 79450
rect 35082 79398 35094 79450
rect 35146 79398 35158 79450
rect 35210 79398 38824 79450
rect 1104 79376 38824 79398
rect 25498 79336 25504 79348
rect 22066 79308 25504 79336
rect 21726 79228 21732 79280
rect 21784 79268 21790 79280
rect 22066 79268 22094 79308
rect 25498 79296 25504 79308
rect 25556 79296 25562 79348
rect 28626 79296 28632 79348
rect 28684 79336 28690 79348
rect 38105 79339 38163 79345
rect 38105 79336 38117 79339
rect 28684 79308 38117 79336
rect 28684 79296 28690 79308
rect 38105 79305 38117 79308
rect 38151 79305 38163 79339
rect 38105 79299 38163 79305
rect 21784 79240 22094 79268
rect 27586 79240 28534 79268
rect 21784 79228 21790 79240
rect 2682 79160 2688 79212
rect 2740 79200 2746 79212
rect 2740 79172 6914 79200
rect 2740 79160 2746 79172
rect 1854 79064 1860 79076
rect 1815 79036 1860 79064
rect 1854 79024 1860 79036
rect 1912 79024 1918 79076
rect 2038 79064 2044 79076
rect 1999 79036 2044 79064
rect 2038 79024 2044 79036
rect 2096 79024 2102 79076
rect 6886 78996 6914 79172
rect 22094 79160 22100 79212
rect 22152 79200 22158 79212
rect 22152 79172 27200 79200
rect 22152 79160 22158 79172
rect 25038 79092 25044 79144
rect 25096 79132 25102 79144
rect 27172 79141 27200 79172
rect 27065 79135 27123 79141
rect 27065 79132 27077 79135
rect 25096 79104 27077 79132
rect 25096 79092 25102 79104
rect 27065 79101 27077 79104
rect 27111 79101 27123 79135
rect 27065 79095 27123 79101
rect 27158 79135 27216 79141
rect 27158 79101 27170 79135
rect 27204 79101 27216 79135
rect 27430 79132 27436 79144
rect 27391 79104 27436 79132
rect 27158 79095 27216 79101
rect 27430 79092 27436 79104
rect 27488 79092 27494 79144
rect 27586 79141 27614 79240
rect 28506 79200 28534 79240
rect 28718 79228 28724 79280
rect 28776 79268 28782 79280
rect 28813 79271 28871 79277
rect 28813 79268 28825 79271
rect 28776 79240 28825 79268
rect 28776 79228 28782 79240
rect 28813 79237 28825 79240
rect 28859 79237 28871 79271
rect 28813 79231 28871 79237
rect 29549 79271 29607 79277
rect 29549 79237 29561 79271
rect 29595 79268 29607 79271
rect 30282 79268 30288 79280
rect 29595 79240 30288 79268
rect 29595 79237 29607 79240
rect 29549 79231 29607 79237
rect 30282 79228 30288 79240
rect 30340 79228 30346 79280
rect 36354 79200 36360 79212
rect 27678 79172 28304 79200
rect 28506 79172 36360 79200
rect 27571 79135 27629 79141
rect 27571 79101 27583 79135
rect 27617 79101 27629 79135
rect 27571 79095 27629 79101
rect 25866 79024 25872 79076
rect 25924 79064 25930 79076
rect 27341 79067 27399 79073
rect 27341 79064 27353 79067
rect 25924 79036 27353 79064
rect 25924 79024 25930 79036
rect 27341 79033 27353 79036
rect 27387 79033 27399 79067
rect 27678 79064 27706 79172
rect 28276 79141 28304 79172
rect 36354 79160 36360 79172
rect 36412 79160 36418 79212
rect 28169 79135 28227 79141
rect 28169 79101 28181 79135
rect 28215 79101 28227 79135
rect 28169 79095 28227 79101
rect 28262 79135 28320 79141
rect 28262 79101 28274 79135
rect 28308 79101 28320 79135
rect 28262 79095 28320 79101
rect 27341 79027 27399 79033
rect 27540 79036 27706 79064
rect 28184 79064 28212 79095
rect 28350 79092 28356 79144
rect 28408 79132 28414 79144
rect 28537 79135 28595 79141
rect 28537 79132 28549 79135
rect 28408 79104 28549 79132
rect 28408 79092 28414 79104
rect 28537 79101 28549 79104
rect 28583 79101 28595 79135
rect 28537 79095 28595 79101
rect 28675 79135 28733 79141
rect 28675 79101 28687 79135
rect 28721 79132 28733 79135
rect 37458 79132 37464 79144
rect 28721 79104 37464 79132
rect 28721 79101 28733 79104
rect 28675 79095 28733 79101
rect 37458 79092 37464 79104
rect 37516 79092 37522 79144
rect 37918 79132 37924 79144
rect 37879 79104 37924 79132
rect 37918 79092 37924 79104
rect 37976 79092 37982 79144
rect 28445 79067 28503 79073
rect 28184 79036 28350 79064
rect 27540 78996 27568 79036
rect 28322 79008 28350 79036
rect 28445 79033 28457 79067
rect 28491 79033 28503 79067
rect 28445 79027 28503 79033
rect 6886 78968 27568 78996
rect 27709 78999 27767 79005
rect 27709 78965 27721 78999
rect 27755 78996 27767 78999
rect 28166 78996 28172 79008
rect 27755 78968 28172 78996
rect 27755 78965 27767 78968
rect 27709 78959 27767 78965
rect 28166 78956 28172 78968
rect 28224 78956 28230 79008
rect 28322 78968 28356 79008
rect 28350 78956 28356 78968
rect 28408 78956 28414 79008
rect 28460 78996 28488 79027
rect 29270 79024 29276 79076
rect 29328 79064 29334 79076
rect 29365 79067 29423 79073
rect 29365 79064 29377 79067
rect 29328 79036 29377 79064
rect 29328 79024 29334 79036
rect 29365 79033 29377 79036
rect 29411 79033 29423 79067
rect 29365 79027 29423 79033
rect 28718 78996 28724 79008
rect 28460 78968 28724 78996
rect 28718 78956 28724 78968
rect 28776 78956 28782 79008
rect 1104 78906 38824 78928
rect 1104 78854 19606 78906
rect 19658 78854 19670 78906
rect 19722 78854 19734 78906
rect 19786 78854 19798 78906
rect 19850 78854 38824 78906
rect 1104 78832 38824 78854
rect 19306 78764 28120 78792
rect 1578 78480 1584 78532
rect 1636 78520 1642 78532
rect 19306 78520 19334 78764
rect 26418 78684 26424 78736
rect 26476 78724 26482 78736
rect 28092 78733 28120 78764
rect 28166 78752 28172 78804
rect 28224 78792 28230 78804
rect 38102 78792 38108 78804
rect 28224 78764 38108 78792
rect 28224 78752 28230 78764
rect 38102 78752 38108 78764
rect 38160 78752 38166 78804
rect 28077 78727 28135 78733
rect 26476 78696 27937 78724
rect 26476 78684 26482 78696
rect 27909 78665 27937 78696
rect 28077 78693 28089 78727
rect 28123 78693 28135 78727
rect 30098 78724 30104 78736
rect 28077 78687 28135 78693
rect 28828 78696 30104 78724
rect 27801 78659 27859 78665
rect 27801 78625 27813 78659
rect 27847 78625 27859 78659
rect 27801 78619 27859 78625
rect 27894 78659 27952 78665
rect 27894 78625 27906 78659
rect 27940 78625 27952 78659
rect 27894 78619 27952 78625
rect 1636 78492 19334 78520
rect 1636 78480 1642 78492
rect 25590 78412 25596 78464
rect 25648 78452 25654 78464
rect 27430 78452 27436 78464
rect 25648 78424 27436 78452
rect 25648 78412 25654 78424
rect 27430 78412 27436 78424
rect 27488 78412 27494 78464
rect 27816 78452 27844 78619
rect 27909 78588 27937 78619
rect 28166 78616 28172 78668
rect 28224 78656 28230 78668
rect 28307 78659 28365 78665
rect 28224 78628 28269 78656
rect 28224 78616 28230 78628
rect 28307 78625 28319 78659
rect 28353 78656 28365 78659
rect 28442 78656 28448 78668
rect 28353 78628 28448 78656
rect 28353 78625 28365 78628
rect 28307 78619 28365 78625
rect 28442 78616 28448 78628
rect 28500 78616 28506 78668
rect 28718 78588 28724 78600
rect 27909 78560 28724 78588
rect 28718 78548 28724 78560
rect 28776 78548 28782 78600
rect 28445 78523 28503 78529
rect 28445 78489 28457 78523
rect 28491 78520 28503 78523
rect 28828 78520 28856 78696
rect 30098 78684 30104 78696
rect 30156 78684 30162 78736
rect 37182 78724 37188 78736
rect 37143 78696 37188 78724
rect 37182 78684 37188 78696
rect 37240 78684 37246 78736
rect 29457 78659 29515 78665
rect 29457 78625 29469 78659
rect 29503 78656 29515 78659
rect 30006 78656 30012 78668
rect 29503 78628 30012 78656
rect 29503 78625 29515 78628
rect 29457 78619 29515 78625
rect 30006 78616 30012 78628
rect 30064 78616 30070 78668
rect 29181 78591 29239 78597
rect 29181 78557 29193 78591
rect 29227 78588 29239 78591
rect 29270 78588 29276 78600
rect 29227 78560 29276 78588
rect 29227 78557 29239 78560
rect 29181 78551 29239 78557
rect 29270 78548 29276 78560
rect 29328 78548 29334 78600
rect 28491 78492 28856 78520
rect 28491 78489 28503 78492
rect 28445 78483 28503 78489
rect 28718 78452 28724 78464
rect 27816 78424 28724 78452
rect 28718 78412 28724 78424
rect 28776 78412 28782 78464
rect 29178 78412 29184 78464
rect 29236 78452 29242 78464
rect 32582 78452 32588 78464
rect 29236 78424 32588 78452
rect 29236 78412 29242 78424
rect 32582 78412 32588 78424
rect 32640 78412 32646 78464
rect 35894 78412 35900 78464
rect 35952 78452 35958 78464
rect 37277 78455 37335 78461
rect 37277 78452 37289 78455
rect 35952 78424 37289 78452
rect 35952 78412 35958 78424
rect 37277 78421 37289 78424
rect 37323 78421 37335 78455
rect 37277 78415 37335 78421
rect 1104 78362 38824 78384
rect 1104 78310 4246 78362
rect 4298 78310 4310 78362
rect 4362 78310 4374 78362
rect 4426 78310 4438 78362
rect 4490 78310 34966 78362
rect 35018 78310 35030 78362
rect 35082 78310 35094 78362
rect 35146 78310 35158 78362
rect 35210 78310 38824 78362
rect 1104 78288 38824 78310
rect 28442 78208 28448 78260
rect 28500 78248 28506 78260
rect 29365 78251 29423 78257
rect 29365 78248 29377 78251
rect 28500 78220 29377 78248
rect 28500 78208 28506 78220
rect 29365 78217 29377 78220
rect 29411 78217 29423 78251
rect 29365 78211 29423 78217
rect 24210 78140 24216 78192
rect 24268 78180 24274 78192
rect 31386 78180 31392 78192
rect 24268 78152 31392 78180
rect 24268 78140 24274 78152
rect 31386 78140 31392 78152
rect 31444 78140 31450 78192
rect 1854 78044 1860 78056
rect 1815 78016 1860 78044
rect 1854 78004 1860 78016
rect 1912 78004 1918 78056
rect 28077 78047 28135 78053
rect 28077 78013 28089 78047
rect 28123 78044 28135 78047
rect 28994 78044 29000 78056
rect 28123 78016 29000 78044
rect 28123 78013 28135 78016
rect 28077 78007 28135 78013
rect 28994 78004 29000 78016
rect 29052 78004 29058 78056
rect 37182 78044 37188 78056
rect 37143 78016 37188 78044
rect 37182 78004 37188 78016
rect 37240 78004 37246 78056
rect 29270 77976 29276 77988
rect 29231 77948 29276 77976
rect 29270 77936 29276 77948
rect 29328 77936 29334 77988
rect 35986 77936 35992 77988
rect 36044 77976 36050 77988
rect 37918 77976 37924 77988
rect 36044 77948 37412 77976
rect 37879 77948 37924 77976
rect 36044 77936 36050 77948
rect 1946 77908 1952 77920
rect 1907 77880 1952 77908
rect 1946 77868 1952 77880
rect 2004 77868 2010 77920
rect 25498 77868 25504 77920
rect 25556 77908 25562 77920
rect 28169 77911 28227 77917
rect 28169 77908 28181 77911
rect 25556 77880 28181 77908
rect 25556 77868 25562 77880
rect 28169 77877 28181 77880
rect 28215 77908 28227 77911
rect 29086 77908 29092 77920
rect 28215 77880 29092 77908
rect 28215 77877 28227 77880
rect 28169 77871 28227 77877
rect 29086 77868 29092 77880
rect 29144 77868 29150 77920
rect 37274 77908 37280 77920
rect 37235 77880 37280 77908
rect 37274 77868 37280 77880
rect 37332 77868 37338 77920
rect 37384 77908 37412 77948
rect 37918 77936 37924 77948
rect 37976 77936 37982 77988
rect 38013 77911 38071 77917
rect 38013 77908 38025 77911
rect 37384 77880 38025 77908
rect 38013 77877 38025 77880
rect 38059 77877 38071 77911
rect 38013 77871 38071 77877
rect 1104 77818 38824 77840
rect 1104 77766 19606 77818
rect 19658 77766 19670 77818
rect 19722 77766 19734 77818
rect 19786 77766 19798 77818
rect 19850 77766 38824 77818
rect 1104 77744 38824 77766
rect 20162 77664 20168 77716
rect 20220 77704 20226 77716
rect 37274 77704 37280 77716
rect 20220 77676 37280 77704
rect 20220 77664 20226 77676
rect 37274 77664 37280 77676
rect 37332 77664 37338 77716
rect 1394 77568 1400 77580
rect 1355 77540 1400 77568
rect 1394 77528 1400 77540
rect 1452 77528 1458 77580
rect 37182 77568 37188 77580
rect 37143 77540 37188 77568
rect 37182 77528 37188 77540
rect 37240 77528 37246 77580
rect 23750 77460 23756 77512
rect 23808 77500 23814 77512
rect 30374 77500 30380 77512
rect 23808 77472 30380 77500
rect 23808 77460 23814 77472
rect 30374 77460 30380 77472
rect 30432 77460 30438 77512
rect 22922 77392 22928 77444
rect 22980 77432 22986 77444
rect 30282 77432 30288 77444
rect 22980 77404 30288 77432
rect 22980 77392 22986 77404
rect 30282 77392 30288 77404
rect 30340 77392 30346 77444
rect 1581 77367 1639 77373
rect 1581 77333 1593 77367
rect 1627 77364 1639 77367
rect 12250 77364 12256 77376
rect 1627 77336 12256 77364
rect 1627 77333 1639 77336
rect 1581 77327 1639 77333
rect 12250 77324 12256 77336
rect 12308 77324 12314 77376
rect 30006 77324 30012 77376
rect 30064 77364 30070 77376
rect 31202 77364 31208 77376
rect 30064 77336 31208 77364
rect 30064 77324 30070 77336
rect 31202 77324 31208 77336
rect 31260 77324 31266 77376
rect 36814 77324 36820 77376
rect 36872 77364 36878 77376
rect 37277 77367 37335 77373
rect 37277 77364 37289 77367
rect 36872 77336 37289 77364
rect 36872 77324 36878 77336
rect 37277 77333 37289 77336
rect 37323 77333 37335 77367
rect 37277 77327 37335 77333
rect 1104 77274 38824 77296
rect 1104 77222 4246 77274
rect 4298 77222 4310 77274
rect 4362 77222 4374 77274
rect 4426 77222 4438 77274
rect 4490 77222 34966 77274
rect 35018 77222 35030 77274
rect 35082 77222 35094 77274
rect 35146 77222 35158 77274
rect 35210 77222 38824 77274
rect 1104 77200 38824 77222
rect 25501 77095 25559 77101
rect 25501 77061 25513 77095
rect 25547 77092 25559 77095
rect 28994 77092 29000 77104
rect 25547 77064 29000 77092
rect 25547 77061 25559 77064
rect 25501 77055 25559 77061
rect 28994 77052 29000 77064
rect 29052 77052 29058 77104
rect 29273 77095 29331 77101
rect 29273 77061 29285 77095
rect 29319 77092 29331 77095
rect 29454 77092 29460 77104
rect 29319 77064 29460 77092
rect 29319 77061 29331 77064
rect 29273 77055 29331 77061
rect 29454 77052 29460 77064
rect 29512 77052 29518 77104
rect 24854 76848 24860 76900
rect 24912 76888 24918 76900
rect 25317 76891 25375 76897
rect 25317 76888 25329 76891
rect 24912 76860 25329 76888
rect 24912 76848 24918 76860
rect 25317 76857 25329 76860
rect 25363 76857 25375 76891
rect 25317 76851 25375 76857
rect 29089 76891 29147 76897
rect 29089 76857 29101 76891
rect 29135 76888 29147 76891
rect 29270 76888 29276 76900
rect 29135 76860 29276 76888
rect 29135 76857 29147 76860
rect 29089 76851 29147 76857
rect 29270 76848 29276 76860
rect 29328 76848 29334 76900
rect 37918 76888 37924 76900
rect 37879 76860 37924 76888
rect 37918 76848 37924 76860
rect 37976 76848 37982 76900
rect 38010 76820 38016 76832
rect 37971 76792 38016 76820
rect 38010 76780 38016 76792
rect 38068 76780 38074 76832
rect 1104 76730 38824 76752
rect 1104 76678 19606 76730
rect 19658 76678 19670 76730
rect 19722 76678 19734 76730
rect 19786 76678 19798 76730
rect 19850 76678 38824 76730
rect 1104 76656 38824 76678
rect 23014 76576 23020 76628
rect 23072 76616 23078 76628
rect 38010 76616 38016 76628
rect 23072 76588 38016 76616
rect 23072 76576 23078 76588
rect 38010 76576 38016 76588
rect 38068 76576 38074 76628
rect 1394 76480 1400 76492
rect 1355 76452 1400 76480
rect 1394 76440 1400 76452
rect 1452 76440 1458 76492
rect 24765 76483 24823 76489
rect 24765 76449 24777 76483
rect 24811 76480 24823 76483
rect 24854 76480 24860 76492
rect 24811 76452 24860 76480
rect 24811 76449 24823 76452
rect 24765 76443 24823 76449
rect 24854 76440 24860 76452
rect 24912 76440 24918 76492
rect 37182 76480 37188 76492
rect 37143 76452 37188 76480
rect 37182 76440 37188 76452
rect 37240 76440 37246 76492
rect 22066 76316 31754 76344
rect 1581 76279 1639 76285
rect 1581 76245 1593 76279
rect 1627 76276 1639 76279
rect 8294 76276 8300 76288
rect 1627 76248 8300 76276
rect 1627 76245 1639 76248
rect 1581 76239 1639 76245
rect 8294 76236 8300 76248
rect 8352 76236 8358 76288
rect 19242 76236 19248 76288
rect 19300 76276 19306 76288
rect 22066 76276 22094 76316
rect 19300 76248 22094 76276
rect 24949 76279 25007 76285
rect 19300 76236 19306 76248
rect 24949 76245 24961 76279
rect 24995 76276 25007 76279
rect 31570 76276 31576 76288
rect 24995 76248 31576 76276
rect 24995 76245 25007 76248
rect 24949 76239 25007 76245
rect 31570 76236 31576 76248
rect 31628 76236 31634 76288
rect 31726 76276 31754 76316
rect 37277 76279 37335 76285
rect 37277 76276 37289 76279
rect 31726 76248 37289 76276
rect 37277 76245 37289 76248
rect 37323 76245 37335 76279
rect 37277 76239 37335 76245
rect 1104 76186 38824 76208
rect 1104 76134 4246 76186
rect 4298 76134 4310 76186
rect 4362 76134 4374 76186
rect 4426 76134 4438 76186
rect 4490 76134 34966 76186
rect 35018 76134 35030 76186
rect 35082 76134 35094 76186
rect 35146 76134 35158 76186
rect 35210 76134 38824 76186
rect 1104 76112 38824 76134
rect 32582 75896 32588 75948
rect 32640 75936 32646 75948
rect 38286 75936 38292 75948
rect 32640 75908 38292 75936
rect 32640 75896 32646 75908
rect 38286 75896 38292 75908
rect 38344 75896 38350 75948
rect 22738 75828 22744 75880
rect 22796 75868 22802 75880
rect 24854 75868 24860 75880
rect 22796 75840 24860 75868
rect 22796 75828 22802 75840
rect 24854 75828 24860 75840
rect 24912 75868 24918 75880
rect 25225 75871 25283 75877
rect 25225 75868 25237 75871
rect 24912 75840 25237 75868
rect 24912 75828 24918 75840
rect 25225 75837 25237 75840
rect 25271 75837 25283 75871
rect 37182 75868 37188 75880
rect 37143 75840 37188 75868
rect 25225 75831 25283 75837
rect 37182 75828 37188 75840
rect 37240 75828 37246 75880
rect 1854 75800 1860 75812
rect 1815 75772 1860 75800
rect 1854 75760 1860 75772
rect 1912 75760 1918 75812
rect 36078 75760 36084 75812
rect 36136 75800 36142 75812
rect 37918 75800 37924 75812
rect 36136 75772 37412 75800
rect 37879 75772 37924 75800
rect 36136 75760 36142 75772
rect 1949 75735 2007 75741
rect 1949 75701 1961 75735
rect 1995 75732 2007 75735
rect 9674 75732 9680 75744
rect 1995 75704 9680 75732
rect 1995 75701 2007 75704
rect 1949 75695 2007 75701
rect 9674 75692 9680 75704
rect 9732 75692 9738 75744
rect 25409 75735 25467 75741
rect 25409 75701 25421 75735
rect 25455 75732 25467 75735
rect 26418 75732 26424 75744
rect 25455 75704 26424 75732
rect 25455 75701 25467 75704
rect 25409 75695 25467 75701
rect 26418 75692 26424 75704
rect 26476 75692 26482 75744
rect 33962 75692 33968 75744
rect 34020 75732 34026 75744
rect 36170 75732 36176 75744
rect 34020 75704 36176 75732
rect 34020 75692 34026 75704
rect 36170 75692 36176 75704
rect 36228 75692 36234 75744
rect 37274 75732 37280 75744
rect 37235 75704 37280 75732
rect 37274 75692 37280 75704
rect 37332 75692 37338 75744
rect 37384 75732 37412 75772
rect 37918 75760 37924 75772
rect 37976 75760 37982 75812
rect 38013 75735 38071 75741
rect 38013 75732 38025 75735
rect 37384 75704 38025 75732
rect 38013 75701 38025 75704
rect 38059 75701 38071 75735
rect 38013 75695 38071 75701
rect 1104 75642 38824 75664
rect 1104 75590 19606 75642
rect 19658 75590 19670 75642
rect 19722 75590 19734 75642
rect 19786 75590 19798 75642
rect 19850 75590 38824 75642
rect 1104 75568 38824 75590
rect 19150 75488 19156 75540
rect 19208 75528 19214 75540
rect 37274 75528 37280 75540
rect 19208 75500 37280 75528
rect 19208 75488 19214 75500
rect 37274 75488 37280 75500
rect 37332 75488 37338 75540
rect 26418 75352 26424 75404
rect 26476 75392 26482 75404
rect 26878 75392 26884 75404
rect 26476 75364 26884 75392
rect 26476 75352 26482 75364
rect 26878 75352 26884 75364
rect 26936 75352 26942 75404
rect 29546 75352 29552 75404
rect 29604 75392 29610 75404
rect 30282 75392 30288 75404
rect 29604 75364 30288 75392
rect 29604 75352 29610 75364
rect 30282 75352 30288 75364
rect 30340 75352 30346 75404
rect 37182 75392 37188 75404
rect 37143 75364 37188 75392
rect 37182 75352 37188 75364
rect 37240 75352 37246 75404
rect 29178 75216 29184 75268
rect 29236 75256 29242 75268
rect 29546 75256 29552 75268
rect 29236 75228 29552 75256
rect 29236 75216 29242 75228
rect 29546 75216 29552 75228
rect 29604 75216 29610 75268
rect 26510 75148 26516 75200
rect 26568 75188 26574 75200
rect 26970 75188 26976 75200
rect 26568 75160 26976 75188
rect 26568 75148 26574 75160
rect 26970 75148 26976 75160
rect 27028 75148 27034 75200
rect 36354 75148 36360 75200
rect 36412 75188 36418 75200
rect 37277 75191 37335 75197
rect 37277 75188 37289 75191
rect 36412 75160 37289 75188
rect 36412 75148 36418 75160
rect 37277 75157 37289 75160
rect 37323 75157 37335 75191
rect 37277 75151 37335 75157
rect 1104 75098 38824 75120
rect 1104 75046 4246 75098
rect 4298 75046 4310 75098
rect 4362 75046 4374 75098
rect 4426 75046 4438 75098
rect 4490 75046 34966 75098
rect 35018 75046 35030 75098
rect 35082 75046 35094 75098
rect 35146 75046 35158 75098
rect 35210 75046 38824 75098
rect 1104 75024 38824 75046
rect 1854 74780 1860 74792
rect 1815 74752 1860 74780
rect 1854 74740 1860 74752
rect 1912 74740 1918 74792
rect 2041 74715 2099 74721
rect 2041 74681 2053 74715
rect 2087 74712 2099 74715
rect 9214 74712 9220 74724
rect 2087 74684 9220 74712
rect 2087 74681 2099 74684
rect 2041 74675 2099 74681
rect 9214 74672 9220 74684
rect 9272 74672 9278 74724
rect 37918 74712 37924 74724
rect 37879 74684 37924 74712
rect 37918 74672 37924 74684
rect 37976 74672 37982 74724
rect 20254 74604 20260 74656
rect 20312 74644 20318 74656
rect 38013 74647 38071 74653
rect 38013 74644 38025 74647
rect 20312 74616 38025 74644
rect 20312 74604 20318 74616
rect 38013 74613 38025 74616
rect 38059 74613 38071 74647
rect 38013 74607 38071 74613
rect 1104 74554 38824 74576
rect 1104 74502 19606 74554
rect 19658 74502 19670 74554
rect 19722 74502 19734 74554
rect 19786 74502 19798 74554
rect 19850 74502 38824 74554
rect 1104 74480 38824 74502
rect 1854 74304 1860 74316
rect 1815 74276 1860 74304
rect 1854 74264 1860 74276
rect 1912 74264 1918 74316
rect 37182 74304 37188 74316
rect 37143 74276 37188 74304
rect 37182 74264 37188 74276
rect 37240 74264 37246 74316
rect 27430 74196 27436 74248
rect 27488 74236 27494 74248
rect 28166 74236 28172 74248
rect 27488 74208 28172 74236
rect 27488 74196 27494 74208
rect 28166 74196 28172 74208
rect 28224 74196 28230 74248
rect 2041 74171 2099 74177
rect 2041 74137 2053 74171
rect 2087 74168 2099 74171
rect 8938 74168 8944 74180
rect 2087 74140 8944 74168
rect 2087 74137 2099 74140
rect 2041 74131 2099 74137
rect 8938 74128 8944 74140
rect 8996 74128 9002 74180
rect 22186 74060 22192 74112
rect 22244 74100 22250 74112
rect 37277 74103 37335 74109
rect 37277 74100 37289 74103
rect 22244 74072 37289 74100
rect 22244 74060 22250 74072
rect 37277 74069 37289 74072
rect 37323 74069 37335 74103
rect 37277 74063 37335 74069
rect 1104 74010 38824 74032
rect 1104 73958 4246 74010
rect 4298 73958 4310 74010
rect 4362 73958 4374 74010
rect 4426 73958 4438 74010
rect 4490 73958 34966 74010
rect 35018 73958 35030 74010
rect 35082 73958 35094 74010
rect 35146 73958 35158 74010
rect 35210 73958 38824 74010
rect 1104 73936 38824 73958
rect 28626 73856 28632 73908
rect 28684 73896 28690 73908
rect 29365 73899 29423 73905
rect 29365 73896 29377 73899
rect 28684 73868 29377 73896
rect 28684 73856 28690 73868
rect 29365 73865 29377 73868
rect 29411 73865 29423 73899
rect 29365 73859 29423 73865
rect 29181 73695 29239 73701
rect 29181 73661 29193 73695
rect 29227 73692 29239 73695
rect 29270 73692 29276 73704
rect 29227 73664 29276 73692
rect 29227 73661 29239 73664
rect 29181 73655 29239 73661
rect 29270 73652 29276 73664
rect 29328 73652 29334 73704
rect 37182 73692 37188 73704
rect 37143 73664 37188 73692
rect 37182 73652 37188 73664
rect 37240 73652 37246 73704
rect 37918 73624 37924 73636
rect 37879 73596 37924 73624
rect 37918 73584 37924 73596
rect 37976 73584 37982 73636
rect 37274 73556 37280 73568
rect 37235 73528 37280 73556
rect 37274 73516 37280 73528
rect 37332 73516 37338 73568
rect 38010 73556 38016 73568
rect 37971 73528 38016 73556
rect 38010 73516 38016 73528
rect 38068 73516 38074 73568
rect 1104 73466 38824 73488
rect 1104 73414 19606 73466
rect 19658 73414 19670 73466
rect 19722 73414 19734 73466
rect 19786 73414 19798 73466
rect 19850 73414 38824 73466
rect 1104 73392 38824 73414
rect 20346 73312 20352 73364
rect 20404 73352 20410 73364
rect 37274 73352 37280 73364
rect 20404 73324 37280 73352
rect 20404 73312 20410 73324
rect 37274 73312 37280 73324
rect 37332 73312 37338 73364
rect 17862 73244 17868 73296
rect 17920 73284 17926 73296
rect 38010 73284 38016 73296
rect 17920 73256 38016 73284
rect 17920 73244 17926 73256
rect 38010 73244 38016 73256
rect 38068 73244 38074 73296
rect 1854 73216 1860 73228
rect 1815 73188 1860 73216
rect 1854 73176 1860 73188
rect 1912 73176 1918 73228
rect 2041 73219 2099 73225
rect 2041 73185 2053 73219
rect 2087 73216 2099 73219
rect 6270 73216 6276 73228
rect 2087 73188 6276 73216
rect 2087 73185 2099 73188
rect 2041 73179 2099 73185
rect 6270 73176 6276 73188
rect 6328 73176 6334 73228
rect 8294 73176 8300 73228
rect 8352 73216 8358 73228
rect 12158 73216 12164 73228
rect 8352 73188 12164 73216
rect 8352 73176 8358 73188
rect 12158 73176 12164 73188
rect 12216 73176 12222 73228
rect 37182 73216 37188 73228
rect 37143 73188 37188 73216
rect 37182 73176 37188 73188
rect 37240 73176 37246 73228
rect 37090 72972 37096 73024
rect 37148 73012 37154 73024
rect 37277 73015 37335 73021
rect 37277 73012 37289 73015
rect 37148 72984 37289 73012
rect 37148 72972 37154 72984
rect 37277 72981 37289 72984
rect 37323 72981 37335 73015
rect 37277 72975 37335 72981
rect 1104 72922 38824 72944
rect 1104 72870 4246 72922
rect 4298 72870 4310 72922
rect 4362 72870 4374 72922
rect 4426 72870 4438 72922
rect 4490 72870 34966 72922
rect 35018 72870 35030 72922
rect 35082 72870 35094 72922
rect 35146 72870 35158 72922
rect 35210 72870 38824 72922
rect 1104 72848 38824 72870
rect 37918 72604 37924 72616
rect 37879 72576 37924 72604
rect 37918 72564 37924 72576
rect 37976 72564 37982 72616
rect 1854 72536 1860 72548
rect 1815 72508 1860 72536
rect 1854 72496 1860 72508
rect 1912 72496 1918 72548
rect 2041 72539 2099 72545
rect 2041 72505 2053 72539
rect 2087 72536 2099 72539
rect 4798 72536 4804 72548
rect 2087 72508 4804 72536
rect 2087 72505 2099 72508
rect 2041 72499 2099 72505
rect 4798 72496 4804 72508
rect 4856 72496 4862 72548
rect 37642 72428 37648 72480
rect 37700 72468 37706 72480
rect 38013 72471 38071 72477
rect 38013 72468 38025 72471
rect 37700 72440 38025 72468
rect 37700 72428 37706 72440
rect 38013 72437 38025 72440
rect 38059 72437 38071 72471
rect 38013 72431 38071 72437
rect 1104 72378 38824 72400
rect 1104 72326 19606 72378
rect 19658 72326 19670 72378
rect 19722 72326 19734 72378
rect 19786 72326 19798 72378
rect 19850 72326 38824 72378
rect 1104 72304 38824 72326
rect 37182 72128 37188 72140
rect 37143 72100 37188 72128
rect 37182 72088 37188 72100
rect 37240 72088 37246 72140
rect 37369 71995 37427 72001
rect 37369 71961 37381 71995
rect 37415 71992 37427 71995
rect 38378 71992 38384 72004
rect 37415 71964 38384 71992
rect 37415 71961 37427 71964
rect 37369 71955 37427 71961
rect 38378 71952 38384 71964
rect 38436 71952 38442 72004
rect 1104 71834 38824 71856
rect 1104 71782 4246 71834
rect 4298 71782 4310 71834
rect 4362 71782 4374 71834
rect 4426 71782 4438 71834
rect 4490 71782 34966 71834
rect 35018 71782 35030 71834
rect 35082 71782 35094 71834
rect 35146 71782 35158 71834
rect 35210 71782 38824 71834
rect 1104 71760 38824 71782
rect 33962 71720 33968 71732
rect 33923 71692 33968 71720
rect 33962 71680 33968 71692
rect 34020 71680 34026 71732
rect 1854 71516 1860 71528
rect 1815 71488 1860 71516
rect 1854 71476 1860 71488
rect 1912 71476 1918 71528
rect 33686 71476 33692 71528
rect 33744 71516 33750 71528
rect 33781 71519 33839 71525
rect 33781 71516 33793 71519
rect 33744 71488 33793 71516
rect 33744 71476 33750 71488
rect 33781 71485 33793 71488
rect 33827 71485 33839 71519
rect 37182 71516 37188 71528
rect 37143 71488 37188 71516
rect 33781 71479 33839 71485
rect 37182 71476 37188 71488
rect 37240 71476 37246 71528
rect 37369 71519 37427 71525
rect 37369 71485 37381 71519
rect 37415 71516 37427 71519
rect 39114 71516 39120 71528
rect 37415 71488 39120 71516
rect 37415 71485 37427 71488
rect 37369 71479 37427 71485
rect 39114 71476 39120 71488
rect 39172 71476 39178 71528
rect 2041 71451 2099 71457
rect 2041 71417 2053 71451
rect 2087 71448 2099 71451
rect 3510 71448 3516 71460
rect 2087 71420 3516 71448
rect 2087 71417 2099 71420
rect 2041 71411 2099 71417
rect 3510 71408 3516 71420
rect 3568 71408 3574 71460
rect 37918 71448 37924 71460
rect 37879 71420 37924 71448
rect 37918 71408 37924 71420
rect 37976 71408 37982 71460
rect 38105 71451 38163 71457
rect 38105 71417 38117 71451
rect 38151 71448 38163 71451
rect 39482 71448 39488 71460
rect 38151 71420 39488 71448
rect 38151 71417 38163 71420
rect 38105 71411 38163 71417
rect 39482 71408 39488 71420
rect 39540 71408 39546 71460
rect 1104 71290 38824 71312
rect 1104 71238 19606 71290
rect 19658 71238 19670 71290
rect 19722 71238 19734 71290
rect 19786 71238 19798 71290
rect 19850 71238 38824 71290
rect 1104 71216 38824 71238
rect 1854 71040 1860 71052
rect 1815 71012 1860 71040
rect 1854 71000 1860 71012
rect 1912 71000 1918 71052
rect 3694 71000 3700 71052
rect 3752 71040 3758 71052
rect 15286 71040 15292 71052
rect 3752 71012 15292 71040
rect 3752 71000 3758 71012
rect 15286 71000 15292 71012
rect 15344 71000 15350 71052
rect 37182 71040 37188 71052
rect 37143 71012 37188 71040
rect 37182 71000 37188 71012
rect 37240 71000 37246 71052
rect 2041 70907 2099 70913
rect 2041 70873 2053 70907
rect 2087 70904 2099 70907
rect 6362 70904 6368 70916
rect 2087 70876 6368 70904
rect 2087 70873 2099 70876
rect 2041 70867 2099 70873
rect 6362 70864 6368 70876
rect 6420 70864 6426 70916
rect 37369 70907 37427 70913
rect 37369 70873 37381 70907
rect 37415 70904 37427 70907
rect 38286 70904 38292 70916
rect 37415 70876 38292 70904
rect 37415 70873 37427 70876
rect 37369 70867 37427 70873
rect 38286 70864 38292 70876
rect 38344 70864 38350 70916
rect 1104 70746 38824 70768
rect 1104 70694 4246 70746
rect 4298 70694 4310 70746
rect 4362 70694 4374 70746
rect 4426 70694 4438 70746
rect 4490 70694 34966 70746
rect 35018 70694 35030 70746
rect 35082 70694 35094 70746
rect 35146 70694 35158 70746
rect 35210 70694 38824 70746
rect 1104 70672 38824 70694
rect 38105 70499 38163 70505
rect 38105 70496 38117 70499
rect 22066 70468 38117 70496
rect 21634 70388 21640 70440
rect 21692 70428 21698 70440
rect 22066 70428 22094 70468
rect 38105 70465 38117 70468
rect 38151 70465 38163 70499
rect 38105 70459 38163 70465
rect 37918 70428 37924 70440
rect 21692 70400 22094 70428
rect 37879 70400 37924 70428
rect 21692 70388 21698 70400
rect 37918 70388 37924 70400
rect 37976 70388 37982 70440
rect 1104 70202 38824 70224
rect 1104 70150 19606 70202
rect 19658 70150 19670 70202
rect 19722 70150 19734 70202
rect 19786 70150 19798 70202
rect 19850 70150 38824 70202
rect 1104 70128 38824 70150
rect 1854 69952 1860 69964
rect 1815 69924 1860 69952
rect 1854 69912 1860 69924
rect 1912 69912 1918 69964
rect 37182 69952 37188 69964
rect 37143 69924 37188 69952
rect 37182 69912 37188 69924
rect 37240 69912 37246 69964
rect 2041 69819 2099 69825
rect 2041 69785 2053 69819
rect 2087 69816 2099 69819
rect 3418 69816 3424 69828
rect 2087 69788 3424 69816
rect 2087 69785 2099 69788
rect 2041 69779 2099 69785
rect 3418 69776 3424 69788
rect 3476 69776 3482 69828
rect 23198 69708 23204 69760
rect 23256 69748 23262 69760
rect 37277 69751 37335 69757
rect 37277 69748 37289 69751
rect 23256 69720 37289 69748
rect 23256 69708 23262 69720
rect 37277 69717 37289 69720
rect 37323 69717 37335 69751
rect 37277 69711 37335 69717
rect 1104 69658 38824 69680
rect 1104 69606 4246 69658
rect 4298 69606 4310 69658
rect 4362 69606 4374 69658
rect 4426 69606 4438 69658
rect 4490 69606 34966 69658
rect 35018 69606 35030 69658
rect 35082 69606 35094 69658
rect 35146 69606 35158 69658
rect 35210 69606 38824 69658
rect 1104 69584 38824 69606
rect 37369 69411 37427 69417
rect 37369 69408 37381 69411
rect 22066 69380 37381 69408
rect 18966 69300 18972 69352
rect 19024 69340 19030 69352
rect 22066 69340 22094 69380
rect 37369 69377 37381 69380
rect 37415 69377 37427 69411
rect 37369 69371 37427 69377
rect 38105 69343 38163 69349
rect 38105 69340 38117 69343
rect 19024 69312 22094 69340
rect 31726 69312 38117 69340
rect 19024 69300 19030 69312
rect 17770 69164 17776 69216
rect 17828 69204 17834 69216
rect 31726 69204 31754 69312
rect 38105 69309 38117 69312
rect 38151 69309 38163 69343
rect 38105 69303 38163 69309
rect 37182 69272 37188 69284
rect 37143 69244 37188 69272
rect 37182 69232 37188 69244
rect 37240 69232 37246 69284
rect 37918 69272 37924 69284
rect 37879 69244 37924 69272
rect 37918 69232 37924 69244
rect 37976 69232 37982 69284
rect 17828 69176 31754 69204
rect 17828 69164 17834 69176
rect 1104 69114 38824 69136
rect 1104 69062 19606 69114
rect 19658 69062 19670 69114
rect 19722 69062 19734 69114
rect 19786 69062 19798 69114
rect 19850 69062 38824 69114
rect 1104 69040 38824 69062
rect 1854 68932 1860 68944
rect 1815 68904 1860 68932
rect 1854 68892 1860 68904
rect 1912 68892 1918 68944
rect 29178 68892 29184 68944
rect 29236 68932 29242 68944
rect 34054 68932 34060 68944
rect 29236 68904 34060 68932
rect 29236 68892 29242 68904
rect 34054 68892 34060 68904
rect 34112 68892 34118 68944
rect 37182 68864 37188 68876
rect 37143 68836 37188 68864
rect 37182 68824 37188 68836
rect 37240 68824 37246 68876
rect 2041 68731 2099 68737
rect 2041 68697 2053 68731
rect 2087 68728 2099 68731
rect 2130 68728 2136 68740
rect 2087 68700 2136 68728
rect 2087 68697 2099 68700
rect 2041 68691 2099 68697
rect 2130 68688 2136 68700
rect 2188 68688 2194 68740
rect 37369 68663 37427 68669
rect 37369 68629 37381 68663
rect 37415 68660 37427 68663
rect 38838 68660 38844 68672
rect 37415 68632 38844 68660
rect 37415 68629 37427 68632
rect 37369 68623 37427 68629
rect 38838 68620 38844 68632
rect 38896 68620 38902 68672
rect 1104 68570 38824 68592
rect 1104 68518 4246 68570
rect 4298 68518 4310 68570
rect 4362 68518 4374 68570
rect 4426 68518 4438 68570
rect 4490 68518 34966 68570
rect 35018 68518 35030 68570
rect 35082 68518 35094 68570
rect 35146 68518 35158 68570
rect 35210 68518 38824 68570
rect 1104 68496 38824 68518
rect 3142 68280 3148 68332
rect 3200 68320 3206 68332
rect 22002 68320 22008 68332
rect 3200 68292 22008 68320
rect 3200 68280 3206 68292
rect 22002 68280 22008 68292
rect 22060 68280 22066 68332
rect 1854 68252 1860 68264
rect 1815 68224 1860 68252
rect 1854 68212 1860 68224
rect 1912 68212 1918 68264
rect 37274 68252 37280 68264
rect 37235 68224 37280 68252
rect 37274 68212 37280 68224
rect 37332 68212 37338 68264
rect 37921 68255 37979 68261
rect 37921 68221 37933 68255
rect 37967 68252 37979 68255
rect 38933 68255 38991 68261
rect 38933 68252 38945 68255
rect 37967 68224 38945 68252
rect 37967 68221 37979 68224
rect 37921 68215 37979 68221
rect 38933 68221 38945 68224
rect 38979 68221 38991 68255
rect 38933 68215 38991 68221
rect 2041 68187 2099 68193
rect 2041 68153 2053 68187
rect 2087 68184 2099 68187
rect 9030 68184 9036 68196
rect 2087 68156 9036 68184
rect 2087 68153 2099 68156
rect 2041 68147 2099 68153
rect 9030 68144 9036 68156
rect 9088 68144 9094 68196
rect 37461 68119 37519 68125
rect 37461 68085 37473 68119
rect 37507 68116 37519 68119
rect 37826 68116 37832 68128
rect 37507 68088 37832 68116
rect 37507 68085 37519 68088
rect 37461 68079 37519 68085
rect 37826 68076 37832 68088
rect 37884 68076 37890 68128
rect 38105 68119 38163 68125
rect 38105 68085 38117 68119
rect 38151 68116 38163 68119
rect 38194 68116 38200 68128
rect 38151 68088 38200 68116
rect 38151 68085 38163 68088
rect 38105 68079 38163 68085
rect 38194 68076 38200 68088
rect 38252 68076 38258 68128
rect 1104 68026 38824 68048
rect 1104 67974 19606 68026
rect 19658 67974 19670 68026
rect 19722 67974 19734 68026
rect 19786 67974 19798 68026
rect 19850 67974 38824 68026
rect 1104 67952 38824 67974
rect 37182 67776 37188 67788
rect 37143 67748 37188 67776
rect 37182 67736 37188 67748
rect 37240 67736 37246 67788
rect 33502 67600 33508 67652
rect 33560 67640 33566 67652
rect 34698 67640 34704 67652
rect 33560 67612 34704 67640
rect 33560 67600 33566 67612
rect 34698 67600 34704 67612
rect 34756 67600 34762 67652
rect 37366 67640 37372 67652
rect 37327 67612 37372 67640
rect 37366 67600 37372 67612
rect 37424 67600 37430 67652
rect 38930 67640 38936 67652
rect 38891 67612 38936 67640
rect 38930 67600 38936 67612
rect 38988 67600 38994 67652
rect 1104 67482 38824 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 34966 67482
rect 35018 67430 35030 67482
rect 35082 67430 35094 67482
rect 35146 67430 35158 67482
rect 35210 67430 38824 67482
rect 1104 67408 38824 67430
rect 37461 67303 37519 67309
rect 37461 67269 37473 67303
rect 37507 67300 37519 67303
rect 38746 67300 38752 67312
rect 37507 67272 38752 67300
rect 37507 67269 37519 67272
rect 37461 67263 37519 67269
rect 38746 67260 38752 67272
rect 38804 67260 38810 67312
rect 1394 67164 1400 67176
rect 1355 67136 1400 67164
rect 1394 67124 1400 67136
rect 1452 67124 1458 67176
rect 37274 67164 37280 67176
rect 37235 67136 37280 67164
rect 37274 67124 37280 67136
rect 37332 67124 37338 67176
rect 37918 67164 37924 67176
rect 37879 67136 37924 67164
rect 37918 67124 37924 67136
rect 37976 67124 37982 67176
rect 1581 67031 1639 67037
rect 1581 66997 1593 67031
rect 1627 67028 1639 67031
rect 7742 67028 7748 67040
rect 1627 67000 7748 67028
rect 1627 66997 1639 67000
rect 1581 66991 1639 66997
rect 7742 66988 7748 67000
rect 7800 66988 7806 67040
rect 38105 67031 38163 67037
rect 38105 66997 38117 67031
rect 38151 67028 38163 67031
rect 38654 67028 38660 67040
rect 38151 67000 38660 67028
rect 38151 66997 38163 67000
rect 38105 66991 38163 66997
rect 38654 66988 38660 67000
rect 38712 66988 38718 67040
rect 1104 66938 38824 66960
rect 1104 66886 19606 66938
rect 19658 66886 19670 66938
rect 19722 66886 19734 66938
rect 19786 66886 19798 66938
rect 19850 66886 38824 66938
rect 1104 66864 38824 66886
rect 1394 66688 1400 66700
rect 1355 66660 1400 66688
rect 1394 66648 1400 66660
rect 1452 66648 1458 66700
rect 1581 66487 1639 66493
rect 1581 66453 1593 66487
rect 1627 66484 1639 66487
rect 2222 66484 2228 66496
rect 1627 66456 2228 66484
rect 1627 66453 1639 66456
rect 1581 66447 1639 66453
rect 2222 66444 2228 66456
rect 2280 66444 2286 66496
rect 1104 66394 38824 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 34966 66394
rect 35018 66342 35030 66394
rect 35082 66342 35094 66394
rect 35146 66342 35158 66394
rect 35210 66342 38824 66394
rect 1104 66320 38824 66342
rect 37461 66215 37519 66221
rect 37461 66181 37473 66215
rect 37507 66212 37519 66215
rect 38562 66212 38568 66224
rect 37507 66184 38568 66212
rect 37507 66181 37519 66184
rect 37461 66175 37519 66181
rect 38562 66172 38568 66184
rect 38620 66172 38626 66224
rect 37274 66076 37280 66088
rect 37235 66048 37280 66076
rect 37274 66036 37280 66048
rect 37332 66036 37338 66088
rect 37918 66076 37924 66088
rect 37879 66048 37924 66076
rect 37918 66036 37924 66048
rect 37976 66036 37982 66088
rect 38105 65943 38163 65949
rect 38105 65909 38117 65943
rect 38151 65940 38163 65943
rect 38838 65940 38844 65952
rect 38151 65912 38844 65940
rect 38151 65909 38163 65912
rect 38105 65903 38163 65909
rect 38838 65900 38844 65912
rect 38896 65900 38902 65952
rect 1104 65850 38824 65872
rect 1104 65798 19606 65850
rect 19658 65798 19670 65850
rect 19722 65798 19734 65850
rect 19786 65798 19798 65850
rect 19850 65798 38824 65850
rect 1104 65776 38824 65798
rect 1394 65600 1400 65612
rect 1355 65572 1400 65600
rect 1394 65560 1400 65572
rect 1452 65560 1458 65612
rect 34698 65560 34704 65612
rect 34756 65600 34762 65612
rect 35526 65600 35532 65612
rect 34756 65572 35532 65600
rect 34756 65560 34762 65572
rect 35526 65560 35532 65572
rect 35584 65560 35590 65612
rect 37182 65600 37188 65612
rect 37143 65572 37188 65600
rect 37182 65560 37188 65572
rect 37240 65560 37246 65612
rect 1946 65492 1952 65544
rect 2004 65532 2010 65544
rect 12986 65532 12992 65544
rect 2004 65504 12992 65532
rect 2004 65492 2010 65504
rect 12986 65492 12992 65504
rect 13044 65492 13050 65544
rect 33318 65492 33324 65544
rect 33376 65532 33382 65544
rect 34054 65532 34060 65544
rect 33376 65504 34060 65532
rect 33376 65492 33382 65504
rect 34054 65492 34060 65504
rect 34112 65492 34118 65544
rect 32858 65424 32864 65476
rect 32916 65464 32922 65476
rect 34790 65464 34796 65476
rect 32916 65436 34796 65464
rect 32916 65424 32922 65436
rect 34790 65424 34796 65436
rect 34848 65424 34854 65476
rect 1581 65399 1639 65405
rect 1581 65365 1593 65399
rect 1627 65396 1639 65399
rect 1670 65396 1676 65408
rect 1627 65368 1676 65396
rect 1627 65365 1639 65368
rect 1581 65359 1639 65365
rect 1670 65356 1676 65368
rect 1728 65356 1734 65408
rect 37369 65399 37427 65405
rect 37369 65365 37381 65399
rect 37415 65396 37427 65399
rect 39574 65396 39580 65408
rect 37415 65368 39580 65396
rect 37415 65365 37427 65368
rect 37369 65359 37427 65365
rect 39574 65356 39580 65368
rect 39632 65356 39638 65408
rect 1104 65306 38824 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 34966 65306
rect 35018 65254 35030 65306
rect 35082 65254 35094 65306
rect 35146 65254 35158 65306
rect 35210 65254 38824 65306
rect 1104 65232 38824 65254
rect 1581 65127 1639 65133
rect 1581 65093 1593 65127
rect 1627 65124 1639 65127
rect 9122 65124 9128 65136
rect 1627 65096 9128 65124
rect 1627 65093 1639 65096
rect 1581 65087 1639 65093
rect 9122 65084 9128 65096
rect 9180 65084 9186 65136
rect 33870 65084 33876 65136
rect 33928 65124 33934 65136
rect 37461 65127 37519 65133
rect 37461 65124 37473 65127
rect 33928 65096 37473 65124
rect 33928 65084 33934 65096
rect 37461 65093 37473 65096
rect 37507 65093 37519 65127
rect 37461 65087 37519 65093
rect 1394 64988 1400 65000
rect 1355 64960 1400 64988
rect 1394 64948 1400 64960
rect 1452 64948 1458 65000
rect 34146 64948 34152 65000
rect 34204 64988 34210 65000
rect 35250 64988 35256 65000
rect 34204 64960 35256 64988
rect 34204 64948 34210 64960
rect 35250 64948 35256 64960
rect 35308 64948 35314 65000
rect 37182 64948 37188 65000
rect 37240 64988 37246 65000
rect 37277 64991 37335 64997
rect 37277 64988 37289 64991
rect 37240 64960 37289 64988
rect 37240 64948 37246 64960
rect 37277 64957 37289 64960
rect 37323 64957 37335 64991
rect 37918 64988 37924 65000
rect 37879 64960 37924 64988
rect 37277 64951 37335 64957
rect 37918 64948 37924 64960
rect 37976 64948 37982 65000
rect 19978 64880 19984 64932
rect 20036 64920 20042 64932
rect 20036 64892 38148 64920
rect 20036 64880 20042 64892
rect 38120 64861 38148 64892
rect 38105 64855 38163 64861
rect 38105 64821 38117 64855
rect 38151 64821 38163 64855
rect 38105 64815 38163 64821
rect 1104 64762 38824 64784
rect 1104 64710 19606 64762
rect 19658 64710 19670 64762
rect 19722 64710 19734 64762
rect 19786 64710 19798 64762
rect 19850 64710 38824 64762
rect 1104 64688 38824 64710
rect 34606 64648 34612 64660
rect 34567 64620 34612 64648
rect 34606 64608 34612 64620
rect 34664 64608 34670 64660
rect 34238 64472 34244 64524
rect 34296 64512 34302 64524
rect 34333 64515 34391 64521
rect 34333 64512 34345 64515
rect 34296 64484 34345 64512
rect 34296 64472 34302 64484
rect 34333 64481 34345 64484
rect 34379 64481 34391 64515
rect 34333 64475 34391 64481
rect 34517 64515 34575 64521
rect 34517 64481 34529 64515
rect 34563 64481 34575 64515
rect 34517 64475 34575 64481
rect 33962 64404 33968 64456
rect 34020 64444 34026 64456
rect 34532 64444 34560 64475
rect 34020 64416 34560 64444
rect 34020 64404 34026 64416
rect 1104 64218 38824 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 34966 64218
rect 35018 64166 35030 64218
rect 35082 64166 35094 64218
rect 35146 64166 35158 64218
rect 35210 64166 38824 64218
rect 1104 64144 38824 64166
rect 15286 64104 15292 64116
rect 15247 64076 15292 64104
rect 15286 64064 15292 64076
rect 15344 64064 15350 64116
rect 34146 64064 34152 64116
rect 34204 64104 34210 64116
rect 34241 64107 34299 64113
rect 34241 64104 34253 64107
rect 34204 64076 34253 64104
rect 34204 64064 34210 64076
rect 34241 64073 34253 64076
rect 34287 64073 34299 64107
rect 34241 64067 34299 64073
rect 33962 63928 33968 63980
rect 34020 63928 34026 63980
rect 1394 63900 1400 63912
rect 1355 63872 1400 63900
rect 1394 63860 1400 63872
rect 1452 63860 1458 63912
rect 33980 63900 34008 63928
rect 34146 63900 34152 63912
rect 33980 63872 34152 63900
rect 34146 63860 34152 63872
rect 34204 63860 34210 63912
rect 37274 63900 37280 63912
rect 37235 63872 37280 63900
rect 37274 63860 37280 63872
rect 37332 63860 37338 63912
rect 37918 63900 37924 63912
rect 37879 63872 37924 63900
rect 37918 63860 37924 63872
rect 37976 63860 37982 63912
rect 15194 63832 15200 63844
rect 15155 63804 15200 63832
rect 15194 63792 15200 63804
rect 15252 63792 15258 63844
rect 33318 63792 33324 63844
rect 33376 63832 33382 63844
rect 33965 63835 34023 63841
rect 33965 63832 33977 63835
rect 33376 63804 33977 63832
rect 33376 63792 33382 63804
rect 33965 63801 33977 63804
rect 34011 63801 34023 63835
rect 33965 63795 34023 63801
rect 34882 63792 34888 63844
rect 34940 63832 34946 63844
rect 34940 63804 38148 63832
rect 34940 63792 34946 63804
rect 1581 63767 1639 63773
rect 1581 63733 1593 63767
rect 1627 63764 1639 63767
rect 7558 63764 7564 63776
rect 1627 63736 7564 63764
rect 1627 63733 1639 63736
rect 1581 63727 1639 63733
rect 7558 63724 7564 63736
rect 7616 63724 7622 63776
rect 34606 63724 34612 63776
rect 34664 63764 34670 63776
rect 38120 63773 38148 63804
rect 37461 63767 37519 63773
rect 37461 63764 37473 63767
rect 34664 63736 37473 63764
rect 34664 63724 34670 63736
rect 37461 63733 37473 63736
rect 37507 63733 37519 63767
rect 37461 63727 37519 63733
rect 38105 63767 38163 63773
rect 38105 63733 38117 63767
rect 38151 63733 38163 63767
rect 38105 63727 38163 63733
rect 1104 63674 38824 63696
rect 1104 63622 19606 63674
rect 19658 63622 19670 63674
rect 19722 63622 19734 63674
rect 19786 63622 19798 63674
rect 19850 63622 38824 63674
rect 1104 63600 38824 63622
rect 22002 63520 22008 63572
rect 22060 63560 22066 63572
rect 34882 63560 34888 63572
rect 22060 63532 34888 63560
rect 22060 63520 22066 63532
rect 34882 63520 34888 63532
rect 34940 63520 34946 63572
rect 35434 63560 35440 63572
rect 35395 63532 35440 63560
rect 35434 63520 35440 63532
rect 35492 63520 35498 63572
rect 36446 63560 36452 63572
rect 36407 63532 36452 63560
rect 36446 63520 36452 63532
rect 36504 63520 36510 63572
rect 32950 63452 32956 63504
rect 33008 63492 33014 63504
rect 33008 63464 34376 63492
rect 33008 63452 33014 63464
rect 1394 63424 1400 63436
rect 1355 63396 1400 63424
rect 1394 63384 1400 63396
rect 1452 63384 1458 63436
rect 33134 63424 33140 63436
rect 33095 63396 33140 63424
rect 33134 63384 33140 63396
rect 33192 63384 33198 63436
rect 33336 63433 33364 63464
rect 33321 63427 33379 63433
rect 33321 63393 33333 63427
rect 33367 63393 33379 63427
rect 33321 63387 33379 63393
rect 33502 63384 33508 63436
rect 33560 63424 33566 63436
rect 33689 63427 33747 63433
rect 33689 63424 33701 63427
rect 33560 63396 33701 63424
rect 33560 63384 33566 63396
rect 33689 63393 33701 63396
rect 33735 63393 33747 63427
rect 33689 63387 33747 63393
rect 33870 63384 33876 63436
rect 33928 63424 33934 63436
rect 34348 63433 34376 63464
rect 34514 63452 34520 63504
rect 34572 63492 34578 63504
rect 34701 63495 34759 63501
rect 34701 63492 34713 63495
rect 34572 63464 34713 63492
rect 34572 63452 34578 63464
rect 34701 63461 34713 63464
rect 34747 63461 34759 63495
rect 36173 63495 36231 63501
rect 36173 63492 36185 63495
rect 34701 63455 34759 63461
rect 34808 63464 36185 63492
rect 34149 63427 34207 63433
rect 34149 63424 34161 63427
rect 33928 63396 34161 63424
rect 33928 63384 33934 63396
rect 34149 63393 34161 63396
rect 34195 63393 34207 63427
rect 34149 63387 34207 63393
rect 34333 63427 34391 63433
rect 34333 63393 34345 63427
rect 34379 63393 34391 63427
rect 34333 63387 34391 63393
rect 20898 63316 20904 63368
rect 20956 63356 20962 63368
rect 34808 63356 34836 63464
rect 36173 63461 36185 63464
rect 36219 63461 36231 63495
rect 36173 63455 36231 63461
rect 35161 63427 35219 63433
rect 35161 63393 35173 63427
rect 35207 63393 35219 63427
rect 35161 63387 35219 63393
rect 20956 63328 34836 63356
rect 20956 63316 20962 63328
rect 20530 63248 20536 63300
rect 20588 63288 20594 63300
rect 35176 63288 35204 63387
rect 35250 63384 35256 63436
rect 35308 63424 35314 63436
rect 35345 63427 35403 63433
rect 35345 63424 35357 63427
rect 35308 63396 35357 63424
rect 35308 63384 35314 63396
rect 35345 63393 35357 63396
rect 35391 63424 35403 63427
rect 36357 63427 36415 63433
rect 36357 63424 36369 63427
rect 35391 63396 36369 63424
rect 35391 63393 35403 63396
rect 35345 63387 35403 63393
rect 36357 63393 36369 63396
rect 36403 63393 36415 63427
rect 37182 63424 37188 63436
rect 37143 63396 37188 63424
rect 36357 63387 36415 63393
rect 37182 63384 37188 63396
rect 37240 63384 37246 63436
rect 20588 63260 35204 63288
rect 20588 63248 20594 63260
rect 1581 63223 1639 63229
rect 1581 63189 1593 63223
rect 1627 63220 1639 63223
rect 9490 63220 9496 63232
rect 1627 63192 9496 63220
rect 1627 63189 1639 63192
rect 1581 63183 1639 63189
rect 9490 63180 9496 63192
rect 9548 63180 9554 63232
rect 32398 63180 32404 63232
rect 32456 63220 32462 63232
rect 34698 63220 34704 63232
rect 32456 63192 34704 63220
rect 32456 63180 32462 63192
rect 34698 63180 34704 63192
rect 34756 63180 34762 63232
rect 37369 63223 37427 63229
rect 37369 63189 37381 63223
rect 37415 63220 37427 63223
rect 38470 63220 38476 63232
rect 37415 63192 38476 63220
rect 37415 63189 37427 63192
rect 37369 63183 37427 63189
rect 38470 63180 38476 63192
rect 38528 63180 38534 63232
rect 1104 63130 38824 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 34966 63130
rect 35018 63078 35030 63130
rect 35082 63078 35094 63130
rect 35146 63078 35158 63130
rect 35210 63078 38824 63130
rect 1104 63056 38824 63078
rect 29086 62976 29092 63028
rect 29144 63016 29150 63028
rect 32398 63016 32404 63028
rect 29144 62988 32404 63016
rect 29144 62976 29150 62988
rect 32398 62976 32404 62988
rect 32456 62976 32462 63028
rect 33042 63016 33048 63028
rect 33003 62988 33048 63016
rect 33042 62976 33048 62988
rect 33100 62976 33106 63028
rect 34057 63019 34115 63025
rect 34057 62985 34069 63019
rect 34103 62985 34115 63019
rect 34057 62979 34115 62985
rect 31754 62908 31760 62960
rect 31812 62948 31818 62960
rect 34072 62948 34100 62979
rect 31812 62920 34100 62948
rect 31812 62908 31818 62920
rect 8938 62840 8944 62892
rect 8996 62880 9002 62892
rect 10042 62880 10048 62892
rect 8996 62852 10048 62880
rect 8996 62840 9002 62852
rect 10042 62840 10048 62852
rect 10100 62840 10106 62892
rect 33042 62840 33048 62892
rect 33100 62880 33106 62892
rect 34146 62880 34152 62892
rect 33100 62852 34152 62880
rect 33100 62840 33106 62852
rect 34146 62840 34152 62852
rect 34204 62880 34210 62892
rect 34974 62880 34980 62892
rect 34204 62852 34980 62880
rect 34204 62840 34210 62852
rect 34974 62840 34980 62852
rect 35032 62880 35038 62892
rect 35250 62880 35256 62892
rect 35032 62852 35256 62880
rect 35032 62840 35038 62852
rect 35250 62840 35256 62852
rect 35308 62840 35314 62892
rect 8018 62772 8024 62824
rect 8076 62812 8082 62824
rect 21450 62812 21456 62824
rect 8076 62784 21456 62812
rect 8076 62772 8082 62784
rect 21450 62772 21456 62784
rect 21508 62772 21514 62824
rect 24578 62772 24584 62824
rect 24636 62812 24642 62824
rect 24762 62812 24768 62824
rect 24636 62784 24768 62812
rect 24636 62772 24642 62784
rect 24762 62772 24768 62784
rect 24820 62772 24826 62824
rect 32950 62812 32956 62824
rect 32911 62784 32956 62812
rect 32950 62772 32956 62784
rect 33008 62812 33014 62824
rect 33965 62815 34023 62821
rect 33965 62812 33977 62815
rect 33008 62784 33977 62812
rect 33008 62772 33014 62784
rect 33965 62781 33977 62784
rect 34011 62781 34023 62815
rect 37274 62812 37280 62824
rect 37235 62784 37280 62812
rect 33965 62775 34023 62781
rect 37274 62772 37280 62784
rect 37332 62772 37338 62824
rect 37918 62812 37924 62824
rect 37879 62784 37924 62812
rect 37918 62772 37924 62784
rect 37976 62772 37982 62824
rect 32122 62704 32128 62756
rect 32180 62744 32186 62756
rect 32769 62747 32827 62753
rect 32769 62744 32781 62747
rect 32180 62716 32781 62744
rect 32180 62704 32186 62716
rect 32769 62713 32781 62716
rect 32815 62713 32827 62747
rect 32769 62707 32827 62713
rect 33781 62747 33839 62753
rect 33781 62713 33793 62747
rect 33827 62713 33839 62747
rect 33781 62707 33839 62713
rect 32398 62636 32404 62688
rect 32456 62676 32462 62688
rect 33796 62676 33824 62707
rect 32456 62648 33824 62676
rect 32456 62636 32462 62648
rect 33962 62636 33968 62688
rect 34020 62676 34026 62688
rect 34146 62676 34152 62688
rect 34020 62648 34152 62676
rect 34020 62636 34026 62648
rect 34146 62636 34152 62648
rect 34204 62636 34210 62688
rect 37458 62676 37464 62688
rect 37419 62648 37464 62676
rect 37458 62636 37464 62648
rect 37516 62636 37522 62688
rect 38102 62676 38108 62688
rect 38063 62648 38108 62676
rect 38102 62636 38108 62648
rect 38160 62636 38166 62688
rect 1104 62586 38824 62608
rect 1104 62534 19606 62586
rect 19658 62534 19670 62586
rect 19722 62534 19734 62586
rect 19786 62534 19798 62586
rect 19850 62534 38824 62586
rect 1104 62512 38824 62534
rect 30009 62475 30067 62481
rect 30009 62441 30021 62475
rect 30055 62472 30067 62475
rect 32950 62472 32956 62484
rect 30055 62444 32956 62472
rect 30055 62441 30067 62444
rect 30009 62435 30067 62441
rect 32950 62432 32956 62444
rect 33008 62472 33014 62484
rect 33008 62444 33733 62472
rect 33008 62432 33014 62444
rect 22830 62364 22836 62416
rect 22888 62404 22894 62416
rect 31754 62404 31760 62416
rect 22888 62376 31760 62404
rect 22888 62364 22894 62376
rect 31754 62364 31760 62376
rect 31812 62364 31818 62416
rect 1394 62336 1400 62348
rect 1355 62308 1400 62336
rect 1394 62296 1400 62308
rect 1452 62296 1458 62348
rect 24302 62296 24308 62348
rect 24360 62336 24366 62348
rect 29914 62336 29920 62348
rect 24360 62308 29920 62336
rect 24360 62296 24366 62308
rect 29914 62296 29920 62308
rect 29972 62336 29978 62348
rect 30745 62339 30803 62345
rect 30745 62336 30757 62339
rect 29972 62308 30757 62336
rect 29972 62296 29978 62308
rect 30745 62305 30757 62308
rect 30791 62305 30803 62339
rect 30745 62299 30803 62305
rect 30929 62339 30987 62345
rect 30929 62305 30941 62339
rect 30975 62336 30987 62339
rect 33042 62336 33048 62348
rect 30975 62308 33048 62336
rect 30975 62305 30987 62308
rect 30929 62299 30987 62305
rect 33042 62296 33048 62308
rect 33100 62296 33106 62348
rect 33705 62345 33733 62444
rect 33778 62364 33784 62416
rect 33836 62404 33842 62416
rect 34057 62407 34115 62413
rect 34057 62404 34069 62407
rect 33836 62376 34069 62404
rect 33836 62364 33842 62376
rect 34057 62373 34069 62376
rect 34103 62373 34115 62407
rect 34057 62367 34115 62373
rect 33413 62339 33471 62345
rect 33413 62305 33425 62339
rect 33459 62336 33471 62339
rect 33505 62339 33563 62345
rect 33505 62336 33517 62339
rect 33459 62308 33517 62336
rect 33459 62305 33471 62308
rect 33413 62299 33471 62305
rect 33505 62305 33517 62308
rect 33551 62305 33563 62339
rect 33505 62299 33563 62305
rect 33689 62339 33747 62345
rect 33689 62305 33701 62339
rect 33735 62305 33747 62339
rect 33689 62299 33747 62305
rect 34793 62339 34851 62345
rect 34793 62305 34805 62339
rect 34839 62305 34851 62339
rect 34974 62336 34980 62348
rect 34935 62308 34980 62336
rect 34793 62299 34851 62305
rect 21174 62228 21180 62280
rect 21232 62268 21238 62280
rect 34808 62268 34836 62299
rect 34974 62296 34980 62308
rect 35032 62296 35038 62348
rect 35342 62336 35348 62348
rect 35303 62308 35348 62336
rect 35342 62296 35348 62308
rect 35400 62296 35406 62348
rect 21232 62240 34836 62268
rect 21232 62228 21238 62240
rect 23106 62160 23112 62212
rect 23164 62200 23170 62212
rect 38102 62200 38108 62212
rect 23164 62172 38108 62200
rect 23164 62160 23170 62172
rect 38102 62160 38108 62172
rect 38160 62160 38166 62212
rect 1581 62135 1639 62141
rect 1581 62101 1593 62135
rect 1627 62132 1639 62135
rect 7834 62132 7840 62144
rect 1627 62104 7840 62132
rect 1627 62101 1639 62104
rect 1581 62095 1639 62101
rect 7834 62092 7840 62104
rect 7892 62092 7898 62144
rect 33413 62135 33471 62141
rect 33413 62101 33425 62135
rect 33459 62132 33471 62135
rect 33870 62132 33876 62144
rect 33459 62104 33876 62132
rect 33459 62101 33471 62104
rect 33413 62095 33471 62101
rect 33870 62092 33876 62104
rect 33928 62092 33934 62144
rect 1104 62042 38824 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 34966 62042
rect 35018 61990 35030 62042
rect 35082 61990 35094 62042
rect 35146 61990 35158 62042
rect 35210 61990 38824 62042
rect 1104 61968 38824 61990
rect 1394 61724 1400 61736
rect 1355 61696 1400 61724
rect 1394 61684 1400 61696
rect 1452 61684 1458 61736
rect 37274 61724 37280 61736
rect 37235 61696 37280 61724
rect 37274 61684 37280 61696
rect 37332 61684 37338 61736
rect 37918 61724 37924 61736
rect 37879 61696 37924 61724
rect 37918 61684 37924 61696
rect 37976 61684 37982 61736
rect 1581 61591 1639 61597
rect 1581 61557 1593 61591
rect 1627 61588 1639 61591
rect 8478 61588 8484 61600
rect 1627 61560 8484 61588
rect 1627 61557 1639 61560
rect 1581 61551 1639 61557
rect 8478 61548 8484 61560
rect 8536 61548 8542 61600
rect 35342 61548 35348 61600
rect 35400 61588 35406 61600
rect 37461 61591 37519 61597
rect 37461 61588 37473 61591
rect 35400 61560 37473 61588
rect 35400 61548 35406 61560
rect 37461 61557 37473 61560
rect 37507 61557 37519 61591
rect 38102 61588 38108 61600
rect 38063 61560 38108 61588
rect 37461 61551 37519 61557
rect 38102 61548 38108 61560
rect 38160 61548 38166 61600
rect 1104 61498 38824 61520
rect 1104 61446 19606 61498
rect 19658 61446 19670 61498
rect 19722 61446 19734 61498
rect 19786 61446 19798 61498
rect 19850 61446 38824 61498
rect 1104 61424 38824 61446
rect 23382 61276 23388 61328
rect 23440 61316 23446 61328
rect 38102 61316 38108 61328
rect 23440 61288 38108 61316
rect 23440 61276 23446 61288
rect 38102 61276 38108 61288
rect 38160 61276 38166 61328
rect 37182 61248 37188 61260
rect 37143 61220 37188 61248
rect 37182 61208 37188 61220
rect 37240 61208 37246 61260
rect 34790 61004 34796 61056
rect 34848 61044 34854 61056
rect 37369 61047 37427 61053
rect 37369 61044 37381 61047
rect 34848 61016 37381 61044
rect 34848 61004 34854 61016
rect 37369 61013 37381 61016
rect 37415 61013 37427 61047
rect 37369 61007 37427 61013
rect 1104 60954 38824 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 34966 60954
rect 35018 60902 35030 60954
rect 35082 60902 35094 60954
rect 35146 60902 35158 60954
rect 35210 60902 38824 60954
rect 1104 60880 38824 60902
rect 28626 60840 28632 60852
rect 26068 60812 28632 60840
rect 1394 60636 1400 60648
rect 1355 60608 1400 60636
rect 1394 60596 1400 60608
rect 1452 60596 1458 60648
rect 25961 60639 26019 60645
rect 25961 60605 25973 60639
rect 26007 60636 26019 60639
rect 26068 60636 26096 60812
rect 28626 60800 28632 60812
rect 28684 60800 28690 60852
rect 34425 60843 34483 60849
rect 34425 60809 34437 60843
rect 34471 60840 34483 60843
rect 35710 60840 35716 60852
rect 34471 60812 35716 60840
rect 34471 60809 34483 60812
rect 34425 60803 34483 60809
rect 35710 60800 35716 60812
rect 35768 60800 35774 60852
rect 26160 60744 28994 60772
rect 26160 60645 26188 60744
rect 26007 60608 26096 60636
rect 26145 60639 26203 60645
rect 26007 60605 26019 60608
rect 25961 60599 26019 60605
rect 26145 60605 26157 60639
rect 26191 60605 26203 60639
rect 26145 60599 26203 60605
rect 26329 60639 26387 60645
rect 26329 60605 26341 60639
rect 26375 60605 26387 60639
rect 26510 60636 26516 60648
rect 26471 60608 26516 60636
rect 26329 60599 26387 60605
rect 24394 60528 24400 60580
rect 24452 60568 24458 60580
rect 24452 60540 26096 60568
rect 24452 60528 24458 60540
rect 1581 60503 1639 60509
rect 1581 60469 1593 60503
rect 1627 60500 1639 60503
rect 6546 60500 6552 60512
rect 1627 60472 6552 60500
rect 1627 60469 1639 60472
rect 1581 60463 1639 60469
rect 6546 60460 6552 60472
rect 6604 60460 6610 60512
rect 25866 60460 25872 60512
rect 25924 60500 25930 60512
rect 25961 60503 26019 60509
rect 25961 60500 25973 60503
rect 25924 60472 25973 60500
rect 25924 60460 25930 60472
rect 25961 60469 25973 60472
rect 26007 60469 26019 60503
rect 26068 60500 26096 60540
rect 26344 60500 26372 60599
rect 26510 60596 26516 60608
rect 26568 60596 26574 60648
rect 28966 60568 28994 60744
rect 30098 60596 30104 60648
rect 30156 60636 30162 60648
rect 34241 60639 34299 60645
rect 34241 60636 34253 60639
rect 30156 60608 34253 60636
rect 30156 60596 30162 60608
rect 34241 60605 34253 60608
rect 34287 60605 34299 60639
rect 37274 60636 37280 60648
rect 37235 60608 37280 60636
rect 34241 60599 34299 60605
rect 37274 60596 37280 60608
rect 37332 60596 37338 60648
rect 37918 60636 37924 60648
rect 37879 60608 37924 60636
rect 37918 60596 37924 60608
rect 37976 60596 37982 60648
rect 29546 60568 29552 60580
rect 28966 60540 29552 60568
rect 29546 60528 29552 60540
rect 29604 60528 29610 60580
rect 37458 60500 37464 60512
rect 26068 60472 26372 60500
rect 37419 60472 37464 60500
rect 25961 60463 26019 60469
rect 37458 60460 37464 60472
rect 37516 60460 37522 60512
rect 38102 60500 38108 60512
rect 38063 60472 38108 60500
rect 38102 60460 38108 60472
rect 38160 60460 38166 60512
rect 1104 60410 38824 60432
rect 1104 60358 19606 60410
rect 19658 60358 19670 60410
rect 19722 60358 19734 60410
rect 19786 60358 19798 60410
rect 19850 60358 38824 60410
rect 1104 60336 38824 60358
rect 18322 60256 18328 60308
rect 18380 60296 18386 60308
rect 38102 60296 38108 60308
rect 18380 60268 38108 60296
rect 18380 60256 18386 60268
rect 38102 60256 38108 60268
rect 38160 60256 38166 60308
rect 18506 60188 18512 60240
rect 18564 60228 18570 60240
rect 37458 60228 37464 60240
rect 18564 60200 37464 60228
rect 18564 60188 18570 60200
rect 37458 60188 37464 60200
rect 37516 60188 37522 60240
rect 1394 60160 1400 60172
rect 1355 60132 1400 60160
rect 1394 60120 1400 60132
rect 1452 60120 1458 60172
rect 37182 60160 37188 60172
rect 37143 60132 37188 60160
rect 37182 60120 37188 60132
rect 37240 60120 37246 60172
rect 26326 59984 26332 60036
rect 26384 60024 26390 60036
rect 27430 60024 27436 60036
rect 26384 59996 27436 60024
rect 26384 59984 26390 59996
rect 27430 59984 27436 59996
rect 27488 59984 27494 60036
rect 37274 59984 37280 60036
rect 37332 60024 37338 60036
rect 39206 60024 39212 60036
rect 37332 59996 39212 60024
rect 37332 59984 37338 59996
rect 39206 59984 39212 59996
rect 39264 59984 39270 60036
rect 1581 59959 1639 59965
rect 1581 59925 1593 59959
rect 1627 59956 1639 59959
rect 8938 59956 8944 59968
rect 1627 59928 8944 59956
rect 1627 59925 1639 59928
rect 1581 59919 1639 59925
rect 8938 59916 8944 59928
rect 8996 59916 9002 59968
rect 19978 59916 19984 59968
rect 20036 59956 20042 59968
rect 37369 59959 37427 59965
rect 37369 59956 37381 59959
rect 20036 59928 37381 59956
rect 20036 59916 20042 59928
rect 37369 59925 37381 59928
rect 37415 59925 37427 59959
rect 37369 59919 37427 59925
rect 1104 59866 38824 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 34966 59866
rect 35018 59814 35030 59866
rect 35082 59814 35094 59866
rect 35146 59814 35158 59866
rect 35210 59814 38824 59866
rect 1104 59792 38824 59814
rect 36722 59752 36728 59764
rect 26804 59724 36728 59752
rect 18782 59576 18788 59628
rect 18840 59616 18846 59628
rect 18840 59588 22094 59616
rect 18840 59576 18846 59588
rect 22066 59480 22094 59588
rect 23290 59576 23296 59628
rect 23348 59616 23354 59628
rect 23348 59588 26556 59616
rect 23348 59576 23354 59588
rect 26234 59548 26240 59560
rect 26195 59520 26240 59548
rect 26234 59508 26240 59520
rect 26292 59508 26298 59560
rect 26528 59557 26556 59588
rect 26804 59557 26832 59724
rect 36722 59712 36728 59724
rect 36780 59712 36786 59764
rect 37093 59687 37151 59693
rect 37093 59684 37105 59687
rect 31726 59656 37105 59684
rect 31726 59616 31754 59656
rect 37093 59653 37105 59656
rect 37139 59653 37151 59687
rect 37093 59647 37151 59653
rect 26896 59588 31754 59616
rect 26513 59551 26571 59557
rect 26513 59517 26525 59551
rect 26559 59517 26571 59551
rect 26513 59511 26571 59517
rect 26789 59551 26847 59557
rect 26789 59517 26801 59551
rect 26835 59517 26847 59551
rect 26789 59511 26847 59517
rect 26896 59480 26924 59588
rect 36538 59576 36544 59628
rect 36596 59616 36602 59628
rect 36814 59616 36820 59628
rect 36596 59588 36820 59616
rect 36596 59576 36602 59588
rect 36814 59576 36820 59588
rect 36872 59576 36878 59628
rect 26973 59551 27031 59557
rect 26973 59517 26985 59551
rect 27019 59548 27031 59551
rect 36906 59548 36912 59560
rect 27019 59520 31754 59548
rect 36867 59520 36912 59548
rect 27019 59517 27031 59520
rect 26973 59511 27031 59517
rect 22066 59452 26924 59480
rect 24486 59372 24492 59424
rect 24544 59412 24550 59424
rect 26329 59415 26387 59421
rect 26329 59412 26341 59415
rect 24544 59384 26341 59412
rect 24544 59372 24550 59384
rect 26329 59381 26341 59384
rect 26375 59381 26387 59415
rect 31726 59412 31754 59520
rect 36906 59508 36912 59520
rect 36964 59508 36970 59560
rect 37274 59508 37280 59560
rect 37332 59548 37338 59560
rect 37553 59551 37611 59557
rect 37553 59548 37565 59551
rect 37332 59520 37565 59548
rect 37332 59508 37338 59520
rect 37553 59517 37565 59520
rect 37599 59517 37611 59551
rect 37734 59548 37740 59560
rect 37695 59520 37740 59548
rect 37553 59511 37611 59517
rect 37734 59508 37740 59520
rect 37792 59508 37798 59560
rect 38010 59557 38016 59560
rect 37967 59551 38016 59557
rect 37967 59517 37979 59551
rect 38013 59517 38016 59551
rect 37967 59511 38016 59517
rect 38010 59508 38016 59511
rect 38068 59508 38074 59560
rect 36722 59440 36728 59492
rect 36780 59480 36786 59492
rect 37825 59483 37883 59489
rect 37825 59480 37837 59483
rect 36780 59452 37837 59480
rect 36780 59440 36786 59452
rect 37825 59449 37837 59452
rect 37871 59449 37883 59483
rect 37825 59443 37883 59449
rect 36262 59412 36268 59424
rect 31726 59384 36268 59412
rect 26329 59375 26387 59381
rect 36262 59372 36268 59384
rect 36320 59372 36326 59424
rect 36814 59372 36820 59424
rect 36872 59412 36878 59424
rect 38105 59415 38163 59421
rect 38105 59412 38117 59415
rect 36872 59384 38117 59412
rect 36872 59372 36878 59384
rect 38105 59381 38117 59384
rect 38151 59381 38163 59415
rect 38105 59375 38163 59381
rect 1104 59322 38824 59344
rect 1104 59270 19606 59322
rect 19658 59270 19670 59322
rect 19722 59270 19734 59322
rect 19786 59270 19798 59322
rect 19850 59270 38824 59322
rect 1104 59248 38824 59270
rect 7282 59100 7288 59152
rect 7340 59140 7346 59152
rect 7650 59140 7656 59152
rect 7340 59112 7656 59140
rect 7340 59100 7346 59112
rect 7650 59100 7656 59112
rect 7708 59140 7714 59152
rect 10229 59143 10287 59149
rect 10229 59140 10241 59143
rect 7708 59112 10241 59140
rect 7708 59100 7714 59112
rect 10229 59109 10241 59112
rect 10275 59109 10287 59143
rect 10229 59103 10287 59109
rect 1394 59072 1400 59084
rect 1355 59044 1400 59072
rect 1394 59032 1400 59044
rect 1452 59032 1458 59084
rect 12250 59072 12256 59084
rect 12211 59044 12256 59072
rect 12250 59032 12256 59044
rect 12308 59032 12314 59084
rect 36446 59072 36452 59084
rect 36407 59044 36452 59072
rect 36446 59032 36452 59044
rect 36504 59032 36510 59084
rect 37182 59072 37188 59084
rect 37143 59044 37188 59072
rect 37182 59032 37188 59044
rect 37240 59032 37246 59084
rect 10413 59007 10471 59013
rect 10413 58973 10425 59007
rect 10459 59004 10471 59007
rect 11974 59004 11980 59016
rect 10459 58976 11980 59004
rect 10459 58973 10471 58976
rect 10413 58967 10471 58973
rect 11974 58964 11980 58976
rect 12032 59004 12038 59016
rect 12069 59007 12127 59013
rect 12069 59004 12081 59007
rect 12032 58976 12081 59004
rect 12032 58964 12038 58976
rect 12069 58973 12081 58976
rect 12115 58973 12127 59007
rect 12069 58967 12127 58973
rect 36354 58964 36360 59016
rect 36412 59004 36418 59016
rect 36998 59004 37004 59016
rect 36412 58976 37004 59004
rect 36412 58964 36418 58976
rect 36998 58964 37004 58976
rect 37056 58964 37062 59016
rect 33962 58896 33968 58948
rect 34020 58936 34026 58948
rect 34330 58936 34336 58948
rect 34020 58908 34336 58936
rect 34020 58896 34026 58908
rect 34330 58896 34336 58908
rect 34388 58896 34394 58948
rect 35250 58896 35256 58948
rect 35308 58936 35314 58948
rect 37369 58939 37427 58945
rect 37369 58936 37381 58939
rect 35308 58908 37381 58936
rect 35308 58896 35314 58908
rect 37369 58905 37381 58908
rect 37415 58905 37427 58939
rect 37369 58899 37427 58905
rect 1578 58868 1584 58880
rect 1539 58840 1584 58868
rect 1578 58828 1584 58840
rect 1636 58828 1642 58880
rect 12437 58871 12495 58877
rect 12437 58837 12449 58871
rect 12483 58868 12495 58871
rect 17310 58868 17316 58880
rect 12483 58840 17316 58868
rect 12483 58837 12495 58840
rect 12437 58831 12495 58837
rect 17310 58828 17316 58840
rect 17368 58828 17374 58880
rect 20806 58828 20812 58880
rect 20864 58868 20870 58880
rect 36633 58871 36691 58877
rect 36633 58868 36645 58871
rect 20864 58840 36645 58868
rect 20864 58828 20870 58840
rect 36633 58837 36645 58840
rect 36679 58837 36691 58871
rect 36633 58831 36691 58837
rect 1104 58778 38824 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 34966 58778
rect 35018 58726 35030 58778
rect 35082 58726 35094 58778
rect 35146 58726 35158 58778
rect 35210 58726 38824 58778
rect 1104 58704 38824 58726
rect 27154 58664 27160 58676
rect 26436 58636 27016 58664
rect 27115 58636 27160 58664
rect 2038 58488 2044 58540
rect 2096 58528 2102 58540
rect 12805 58531 12863 58537
rect 12805 58528 12817 58531
rect 2096 58500 12204 58528
rect 2096 58488 2102 58500
rect 1394 58460 1400 58472
rect 1355 58432 1400 58460
rect 1394 58420 1400 58432
rect 1452 58420 1458 58472
rect 12176 58469 12204 58500
rect 12406 58500 12817 58528
rect 12069 58463 12127 58469
rect 12069 58429 12081 58463
rect 12115 58429 12127 58463
rect 12069 58423 12127 58429
rect 12161 58463 12219 58469
rect 12161 58429 12173 58463
rect 12207 58429 12219 58463
rect 12161 58423 12219 58429
rect 11974 58352 11980 58404
rect 12032 58392 12038 58404
rect 12084 58392 12112 58423
rect 12406 58392 12434 58500
rect 12805 58497 12817 58500
rect 12851 58528 12863 58531
rect 26234 58528 26240 58540
rect 12851 58500 26240 58528
rect 12851 58497 12863 58500
rect 12805 58491 12863 58497
rect 26234 58488 26240 58500
rect 26292 58488 26298 58540
rect 12986 58460 12992 58472
rect 12947 58432 12992 58460
rect 12986 58420 12992 58432
rect 13044 58420 13050 58472
rect 26436 58460 26464 58636
rect 26988 58596 27016 58636
rect 27154 58624 27160 58636
rect 27212 58624 27218 58676
rect 35894 58624 35900 58676
rect 35952 58664 35958 58676
rect 38010 58664 38016 58676
rect 35952 58636 38016 58664
rect 35952 58624 35958 58636
rect 38010 58624 38016 58636
rect 38068 58624 38074 58676
rect 34330 58596 34336 58608
rect 26988 58568 34336 58596
rect 34330 58556 34336 58568
rect 34388 58556 34394 58608
rect 36998 58556 37004 58608
rect 37056 58596 37062 58608
rect 37056 58568 37964 58596
rect 37056 58556 37062 58568
rect 26510 58488 26516 58540
rect 26568 58528 26574 58540
rect 26568 58500 26924 58528
rect 26568 58488 26574 58500
rect 26896 58469 26924 58500
rect 36722 58488 36728 58540
rect 36780 58528 36786 58540
rect 36780 58500 37872 58528
rect 36780 58488 36786 58500
rect 26605 58463 26663 58469
rect 26605 58460 26617 58463
rect 26436 58432 26617 58460
rect 26605 58429 26617 58432
rect 26651 58429 26663 58463
rect 26605 58423 26663 58429
rect 26881 58463 26939 58469
rect 26881 58429 26893 58463
rect 26927 58429 26939 58463
rect 26881 58423 26939 58429
rect 26973 58463 27031 58469
rect 26973 58429 26985 58463
rect 27019 58429 27031 58463
rect 26973 58423 27031 58429
rect 12032 58364 12434 58392
rect 12032 58352 12038 58364
rect 26234 58352 26240 58404
rect 26292 58392 26298 58404
rect 26789 58395 26847 58401
rect 26789 58392 26801 58395
rect 26292 58364 26801 58392
rect 26292 58352 26298 58364
rect 26789 58361 26801 58364
rect 26835 58361 26847 58395
rect 26789 58355 26847 58361
rect 1581 58327 1639 58333
rect 1581 58293 1593 58327
rect 1627 58324 1639 58327
rect 1762 58324 1768 58336
rect 1627 58296 1768 58324
rect 1627 58293 1639 58296
rect 1581 58287 1639 58293
rect 1762 58284 1768 58296
rect 1820 58284 1826 58336
rect 12342 58324 12348 58336
rect 12303 58296 12348 58324
rect 12342 58284 12348 58296
rect 12400 58284 12406 58336
rect 13173 58327 13231 58333
rect 13173 58293 13185 58327
rect 13219 58324 13231 58327
rect 17494 58324 17500 58336
rect 13219 58296 17500 58324
rect 13219 58293 13231 58296
rect 13173 58287 13231 58293
rect 17494 58284 17500 58296
rect 17552 58284 17558 58336
rect 18046 58284 18052 58336
rect 18104 58324 18110 58336
rect 26988 58324 27016 58423
rect 35986 58420 35992 58472
rect 36044 58460 36050 58472
rect 36354 58460 36360 58472
rect 36044 58432 36360 58460
rect 36044 58420 36050 58432
rect 36354 58420 36360 58432
rect 36412 58420 36418 58472
rect 36446 58420 36452 58472
rect 36504 58460 36510 58472
rect 36832 58469 36860 58500
rect 36541 58463 36599 58469
rect 36541 58460 36553 58463
rect 36504 58432 36553 58460
rect 36504 58420 36510 58432
rect 36541 58429 36553 58432
rect 36587 58429 36599 58463
rect 36541 58423 36599 58429
rect 36817 58463 36875 58469
rect 36817 58429 36829 58463
rect 36863 58429 36875 58463
rect 36817 58423 36875 58429
rect 36906 58420 36912 58472
rect 36964 58460 36970 58472
rect 37550 58460 37556 58472
rect 36964 58432 37009 58460
rect 37511 58432 37556 58460
rect 36964 58420 36970 58432
rect 37550 58420 37556 58432
rect 37608 58420 37614 58472
rect 37844 58469 37872 58500
rect 37936 58469 37964 58568
rect 37829 58463 37887 58469
rect 37829 58429 37841 58463
rect 37875 58429 37887 58463
rect 37829 58423 37887 58429
rect 37921 58463 37979 58469
rect 37921 58429 37933 58463
rect 37967 58429 37979 58463
rect 37921 58423 37979 58429
rect 36725 58395 36783 58401
rect 36725 58361 36737 58395
rect 36771 58392 36783 58395
rect 37734 58392 37740 58404
rect 36771 58364 37740 58392
rect 36771 58361 36783 58364
rect 36725 58355 36783 58361
rect 37734 58352 37740 58364
rect 37792 58352 37798 58404
rect 37844 58392 37872 58423
rect 38933 58395 38991 58401
rect 38933 58392 38945 58395
rect 37844 58364 38945 58392
rect 38933 58361 38945 58364
rect 38979 58361 38991 58395
rect 38933 58355 38991 58361
rect 18104 58296 27016 58324
rect 18104 58284 18110 58296
rect 35986 58284 35992 58336
rect 36044 58324 36050 58336
rect 37093 58327 37151 58333
rect 37093 58324 37105 58327
rect 36044 58296 37105 58324
rect 36044 58284 36050 58296
rect 37093 58293 37105 58296
rect 37139 58293 37151 58327
rect 38102 58324 38108 58336
rect 38063 58296 38108 58324
rect 37093 58287 37151 58293
rect 38102 58284 38108 58296
rect 38160 58284 38166 58336
rect 1104 58234 38824 58256
rect 1104 58182 19606 58234
rect 19658 58182 19670 58234
rect 19722 58182 19734 58234
rect 19786 58182 19798 58234
rect 19850 58182 38824 58234
rect 1104 58160 38824 58182
rect 26786 58080 26792 58132
rect 26844 58120 26850 58132
rect 27154 58120 27160 58132
rect 26844 58092 27160 58120
rect 26844 58080 26850 58092
rect 27154 58080 27160 58092
rect 27212 58080 27218 58132
rect 11974 57944 11980 57996
rect 12032 57984 12038 57996
rect 12069 57987 12127 57993
rect 12069 57984 12081 57987
rect 12032 57956 12081 57984
rect 12032 57944 12038 57956
rect 12069 57953 12081 57956
rect 12115 57953 12127 57987
rect 12069 57947 12127 57953
rect 12158 57944 12164 57996
rect 12216 57984 12222 57996
rect 12253 57987 12311 57993
rect 12253 57984 12265 57987
rect 12216 57956 12265 57984
rect 12216 57944 12222 57956
rect 12253 57953 12265 57956
rect 12299 57953 12311 57987
rect 12253 57947 12311 57953
rect 12434 57944 12440 57996
rect 12492 57984 12498 57996
rect 36446 57984 36452 57996
rect 12492 57956 12537 57984
rect 36407 57956 36452 57984
rect 12492 57944 12498 57956
rect 36446 57944 36452 57956
rect 36504 57944 36510 57996
rect 36722 57944 36728 57996
rect 36780 57984 36786 57996
rect 36998 57984 37004 57996
rect 36780 57956 37004 57984
rect 36780 57944 36786 57956
rect 36998 57944 37004 57956
rect 37056 57944 37062 57996
rect 37182 57984 37188 57996
rect 37143 57956 37188 57984
rect 37182 57944 37188 57956
rect 37240 57944 37246 57996
rect 9030 57876 9036 57928
rect 9088 57916 9094 57928
rect 10502 57916 10508 57928
rect 9088 57888 10508 57916
rect 9088 57876 9094 57888
rect 10502 57876 10508 57888
rect 10560 57876 10566 57928
rect 20162 57876 20168 57928
rect 20220 57916 20226 57928
rect 20622 57916 20628 57928
rect 20220 57888 20628 57916
rect 20220 57876 20226 57888
rect 20622 57876 20628 57888
rect 20680 57876 20686 57928
rect 22278 57876 22284 57928
rect 22336 57916 22342 57928
rect 28534 57916 28540 57928
rect 22336 57888 28540 57916
rect 22336 57876 22342 57888
rect 28534 57876 28540 57888
rect 28592 57876 28598 57928
rect 25222 57808 25228 57860
rect 25280 57848 25286 57860
rect 27430 57848 27436 57860
rect 25280 57820 27436 57848
rect 25280 57808 25286 57820
rect 27430 57808 27436 57820
rect 27488 57808 27494 57860
rect 37369 57851 37427 57857
rect 37369 57848 37381 57851
rect 31726 57820 37381 57848
rect 18874 57740 18880 57792
rect 18932 57780 18938 57792
rect 31726 57780 31754 57820
rect 37369 57817 37381 57820
rect 37415 57817 37427 57851
rect 37369 57811 37427 57817
rect 36538 57780 36544 57792
rect 18932 57752 31754 57780
rect 36499 57752 36544 57780
rect 18932 57740 18938 57752
rect 36538 57740 36544 57752
rect 36596 57740 36602 57792
rect 1104 57690 38824 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 38824 57690
rect 1104 57616 38824 57638
rect 21818 57536 21824 57588
rect 21876 57576 21882 57588
rect 27157 57579 27215 57585
rect 27157 57576 27169 57579
rect 21876 57548 27169 57576
rect 21876 57536 21882 57548
rect 27157 57545 27169 57548
rect 27203 57545 27215 57579
rect 27157 57539 27215 57545
rect 27430 57536 27436 57588
rect 27488 57576 27494 57588
rect 36538 57576 36544 57588
rect 27488 57548 36544 57576
rect 27488 57536 27494 57548
rect 36538 57536 36544 57548
rect 36596 57536 36602 57588
rect 20530 57468 20536 57520
rect 20588 57508 20594 57520
rect 37093 57511 37151 57517
rect 37093 57508 37105 57511
rect 20588 57480 37105 57508
rect 20588 57468 20594 57480
rect 37093 57477 37105 57480
rect 37139 57477 37151 57511
rect 37093 57471 37151 57477
rect 26510 57400 26516 57452
rect 26568 57440 26574 57452
rect 26568 57412 27292 57440
rect 26568 57400 26574 57412
rect 1394 57372 1400 57384
rect 1355 57344 1400 57372
rect 1394 57332 1400 57344
rect 1452 57332 1458 57384
rect 25590 57332 25596 57384
rect 25648 57372 25654 57384
rect 26896 57381 26924 57412
rect 26605 57375 26663 57381
rect 26605 57372 26617 57375
rect 25648 57344 26617 57372
rect 25648 57332 25654 57344
rect 26605 57341 26617 57344
rect 26651 57341 26663 57375
rect 26789 57375 26847 57381
rect 26789 57372 26801 57375
rect 26605 57335 26663 57341
rect 26712 57344 26801 57372
rect 17218 57264 17224 57316
rect 17276 57304 17282 57316
rect 17276 57276 17954 57304
rect 17276 57264 17282 57276
rect 1581 57239 1639 57245
rect 1581 57205 1593 57239
rect 1627 57236 1639 57239
rect 3602 57236 3608 57248
rect 1627 57208 3608 57236
rect 1627 57205 1639 57208
rect 1581 57199 1639 57205
rect 3602 57196 3608 57208
rect 3660 57196 3666 57248
rect 17926 57236 17954 57276
rect 26234 57264 26240 57316
rect 26292 57304 26298 57316
rect 26712 57304 26740 57344
rect 26789 57341 26801 57344
rect 26835 57341 26847 57375
rect 26789 57335 26847 57341
rect 26881 57375 26939 57381
rect 26881 57341 26893 57375
rect 26927 57341 26939 57375
rect 26881 57335 26939 57341
rect 27019 57375 27077 57381
rect 27019 57341 27031 57375
rect 27065 57372 27077 57375
rect 27264 57372 27292 57412
rect 28626 57400 28632 57452
rect 28684 57440 28690 57452
rect 34698 57440 34704 57452
rect 28684 57412 34704 57440
rect 28684 57400 28690 57412
rect 34698 57400 34704 57412
rect 34756 57400 34762 57452
rect 39390 57440 39396 57452
rect 37568 57412 39396 57440
rect 29181 57375 29239 57381
rect 29181 57372 29193 57375
rect 27065 57344 27200 57372
rect 27264 57344 29193 57372
rect 27065 57341 27077 57344
rect 27019 57335 27077 57341
rect 26292 57276 26740 57304
rect 26292 57264 26298 57276
rect 27172 57236 27200 57344
rect 29181 57341 29193 57344
rect 29227 57341 29239 57375
rect 32582 57372 32588 57384
rect 29181 57335 29239 57341
rect 31726 57344 32588 57372
rect 28997 57307 29055 57313
rect 28997 57273 29009 57307
rect 29043 57304 29055 57307
rect 29362 57304 29368 57316
rect 29043 57276 29368 57304
rect 29043 57273 29055 57276
rect 28997 57267 29055 57273
rect 29362 57264 29368 57276
rect 29420 57304 29426 57316
rect 31726 57304 31754 57344
rect 32582 57332 32588 57344
rect 32640 57332 32646 57384
rect 36909 57375 36967 57381
rect 36909 57341 36921 57375
rect 36955 57372 36967 57375
rect 36998 57372 37004 57384
rect 36955 57344 37004 57372
rect 36955 57341 36967 57344
rect 36909 57335 36967 57341
rect 36998 57332 37004 57344
rect 37056 57332 37062 57384
rect 37568 57381 37596 57412
rect 39390 57400 39396 57412
rect 39448 57400 39454 57452
rect 37553 57375 37611 57381
rect 37553 57341 37565 57375
rect 37599 57341 37611 57375
rect 37553 57335 37611 57341
rect 37921 57375 37979 57381
rect 37921 57341 37933 57375
rect 37967 57372 37979 57375
rect 38010 57372 38016 57384
rect 37967 57344 38016 57372
rect 37967 57341 37979 57344
rect 37921 57335 37979 57341
rect 38010 57332 38016 57344
rect 38068 57332 38074 57384
rect 29420 57276 31754 57304
rect 29420 57264 29426 57276
rect 37274 57264 37280 57316
rect 37332 57304 37338 57316
rect 37734 57304 37740 57316
rect 37332 57276 37740 57304
rect 37332 57264 37338 57276
rect 37734 57264 37740 57276
rect 37792 57264 37798 57316
rect 37829 57307 37887 57313
rect 37829 57273 37841 57307
rect 37875 57304 37887 57307
rect 38933 57307 38991 57313
rect 38933 57304 38945 57307
rect 37875 57276 38945 57304
rect 37875 57273 37887 57276
rect 37829 57267 37887 57273
rect 38933 57273 38945 57276
rect 38979 57304 38991 57307
rect 39206 57304 39212 57316
rect 38979 57276 39212 57304
rect 38979 57273 38991 57276
rect 38933 57267 38991 57273
rect 39206 57264 39212 57276
rect 39264 57264 39270 57316
rect 17926 57208 27200 57236
rect 37550 57196 37556 57248
rect 37608 57236 37614 57248
rect 38105 57239 38163 57245
rect 38105 57236 38117 57239
rect 37608 57208 38117 57236
rect 37608 57196 37614 57208
rect 38105 57205 38117 57208
rect 38151 57205 38163 57239
rect 38105 57199 38163 57205
rect 1104 57146 38824 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 38824 57146
rect 1104 57072 38824 57094
rect 1578 56992 1584 57044
rect 1636 57032 1642 57044
rect 5074 57032 5080 57044
rect 1636 57004 5080 57032
rect 1636 56992 1642 57004
rect 5074 56992 5080 57004
rect 5132 56992 5138 57044
rect 7006 56992 7012 57044
rect 7064 57032 7070 57044
rect 7064 57004 17954 57032
rect 7064 56992 7070 57004
rect 8294 56924 8300 56976
rect 8352 56964 8358 56976
rect 17218 56964 17224 56976
rect 8352 56936 17224 56964
rect 8352 56924 8358 56936
rect 17218 56924 17224 56936
rect 17276 56924 17282 56976
rect 1394 56896 1400 56908
rect 1355 56868 1400 56896
rect 1394 56856 1400 56868
rect 1452 56856 1458 56908
rect 17926 56828 17954 57004
rect 26510 56992 26516 57044
rect 26568 57032 26574 57044
rect 26568 57004 26648 57032
rect 26568 56992 26574 57004
rect 26620 56973 26648 57004
rect 27522 56992 27528 57044
rect 27580 56992 27586 57044
rect 35802 56992 35808 57044
rect 35860 57032 35866 57044
rect 38102 57032 38108 57044
rect 35860 57004 38108 57032
rect 35860 56992 35866 57004
rect 38102 56992 38108 57004
rect 38160 56992 38166 57044
rect 26605 56967 26663 56973
rect 26605 56933 26617 56967
rect 26651 56964 26663 56967
rect 26878 56964 26884 56976
rect 26651 56936 26884 56964
rect 26651 56933 26663 56936
rect 26605 56927 26663 56933
rect 26878 56924 26884 56936
rect 26936 56924 26942 56976
rect 27540 56964 27568 56992
rect 34514 56964 34520 56976
rect 27172 56936 27568 56964
rect 28966 56936 34520 56964
rect 26510 56905 26516 56908
rect 26237 56899 26295 56905
rect 26237 56865 26249 56899
rect 26283 56896 26295 56899
rect 26329 56899 26387 56905
rect 26329 56896 26341 56899
rect 26283 56868 26341 56896
rect 26283 56865 26295 56868
rect 26237 56859 26295 56865
rect 26329 56865 26341 56868
rect 26375 56865 26387 56899
rect 26329 56859 26387 56865
rect 26467 56899 26516 56905
rect 26467 56865 26479 56899
rect 26513 56865 26516 56899
rect 26467 56859 26516 56865
rect 26510 56856 26516 56859
rect 26568 56856 26574 56908
rect 26721 56899 26779 56905
rect 26721 56896 26733 56899
rect 26616 56868 26733 56896
rect 26616 56828 26644 56868
rect 26721 56865 26733 56868
rect 26767 56865 26779 56899
rect 26721 56859 26779 56865
rect 17926 56800 26644 56828
rect 18230 56720 18236 56772
rect 18288 56760 18294 56772
rect 26881 56763 26939 56769
rect 18288 56732 26832 56760
rect 18288 56720 18294 56732
rect 1578 56692 1584 56704
rect 1539 56664 1584 56692
rect 1578 56652 1584 56664
rect 1636 56652 1642 56704
rect 26237 56695 26295 56701
rect 26237 56661 26249 56695
rect 26283 56692 26295 56695
rect 26510 56692 26516 56704
rect 26283 56664 26516 56692
rect 26283 56661 26295 56664
rect 26237 56655 26295 56661
rect 26510 56652 26516 56664
rect 26568 56652 26574 56704
rect 26804 56692 26832 56732
rect 26881 56729 26893 56763
rect 26927 56760 26939 56763
rect 27172 56760 27200 56936
rect 27522 56856 27528 56908
rect 27580 56896 27586 56908
rect 28966 56896 28994 56936
rect 34514 56924 34520 56936
rect 34572 56924 34578 56976
rect 36446 56964 36452 56976
rect 36407 56936 36452 56964
rect 36446 56924 36452 56936
rect 36504 56924 36510 56976
rect 37182 56896 37188 56908
rect 27580 56868 28994 56896
rect 37143 56868 37188 56896
rect 27580 56856 27586 56868
rect 37182 56856 37188 56868
rect 37240 56856 37246 56908
rect 28534 56788 28540 56840
rect 28592 56828 28598 56840
rect 36633 56831 36691 56837
rect 36633 56828 36645 56831
rect 28592 56800 36645 56828
rect 28592 56788 28598 56800
rect 36633 56797 36645 56800
rect 36679 56797 36691 56831
rect 36633 56791 36691 56797
rect 37369 56763 37427 56769
rect 37369 56760 37381 56763
rect 26927 56732 27200 56760
rect 28966 56732 37381 56760
rect 26927 56729 26939 56732
rect 26881 56723 26939 56729
rect 28966 56692 28994 56732
rect 37369 56729 37381 56732
rect 37415 56729 37427 56763
rect 37369 56723 37427 56729
rect 26804 56664 28994 56692
rect 1104 56602 38824 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 38824 56602
rect 1104 56528 38824 56550
rect 9122 56448 9128 56500
rect 9180 56488 9186 56500
rect 9766 56488 9772 56500
rect 9180 56460 9772 56488
rect 9180 56448 9186 56460
rect 9766 56448 9772 56460
rect 9824 56448 9830 56500
rect 27249 56491 27307 56497
rect 26625 56460 27108 56488
rect 26625 56284 26653 56460
rect 26878 56312 26884 56364
rect 26936 56312 26942 56364
rect 27080 56352 27108 56460
rect 27249 56457 27261 56491
rect 27295 56488 27307 56491
rect 27614 56488 27620 56500
rect 27295 56460 27620 56488
rect 27295 56457 27307 56460
rect 27249 56451 27307 56457
rect 27614 56448 27620 56460
rect 27672 56448 27678 56500
rect 32950 56448 32956 56500
rect 33008 56488 33014 56500
rect 36817 56491 36875 56497
rect 36817 56488 36829 56491
rect 33008 56460 36829 56488
rect 33008 56448 33014 56460
rect 36817 56457 36829 56460
rect 36863 56457 36875 56491
rect 36817 56451 36875 56457
rect 37274 56448 37280 56500
rect 37332 56488 37338 56500
rect 37461 56491 37519 56497
rect 37461 56488 37473 56491
rect 37332 56460 37473 56488
rect 37332 56448 37338 56460
rect 37461 56457 37473 56460
rect 37507 56457 37519 56491
rect 37461 56451 37519 56457
rect 27522 56380 27528 56432
rect 27580 56420 27586 56432
rect 28810 56420 28816 56432
rect 27580 56392 28816 56420
rect 27580 56380 27586 56392
rect 28810 56380 28816 56392
rect 28868 56380 28874 56432
rect 31726 56392 34192 56420
rect 29914 56352 29920 56364
rect 27080 56324 29920 56352
rect 29914 56312 29920 56324
rect 29972 56312 29978 56364
rect 26697 56287 26755 56293
rect 26697 56284 26709 56287
rect 26625 56256 26709 56284
rect 26697 56253 26709 56256
rect 26743 56253 26755 56287
rect 26896 56284 26924 56312
rect 26973 56287 27031 56293
rect 26973 56284 26985 56287
rect 26896 56256 26985 56284
rect 26697 56247 26755 56253
rect 26973 56253 26985 56256
rect 27019 56253 27031 56287
rect 26973 56247 27031 56253
rect 27065 56287 27123 56293
rect 27065 56253 27077 56287
rect 27111 56253 27123 56287
rect 27065 56247 27123 56253
rect 26234 56176 26240 56228
rect 26292 56216 26298 56228
rect 26878 56216 26884 56228
rect 26292 56188 26884 56216
rect 26292 56176 26298 56188
rect 26878 56176 26884 56188
rect 26936 56176 26942 56228
rect 8386 56108 8392 56160
rect 8444 56148 8450 56160
rect 27080 56148 27108 56247
rect 28626 56244 28632 56296
rect 28684 56284 28690 56296
rect 31726 56284 31754 56392
rect 28684 56256 31754 56284
rect 28684 56244 28690 56256
rect 27614 56176 27620 56228
rect 27672 56216 27678 56228
rect 34054 56216 34060 56228
rect 27672 56188 34060 56216
rect 27672 56176 27678 56188
rect 34054 56176 34060 56188
rect 34112 56176 34118 56228
rect 8444 56120 27108 56148
rect 34164 56148 34192 56392
rect 36538 56380 36544 56432
rect 36596 56420 36602 56432
rect 37182 56420 37188 56432
rect 36596 56392 37188 56420
rect 36596 56380 36602 56392
rect 37182 56380 37188 56392
rect 37240 56380 37246 56432
rect 35802 56244 35808 56296
rect 35860 56284 35866 56296
rect 36173 56287 36231 56293
rect 36173 56284 36185 56287
rect 35860 56256 36185 56284
rect 35860 56244 35866 56256
rect 36173 56253 36185 56256
rect 36219 56253 36231 56287
rect 36173 56247 36231 56253
rect 36266 56287 36324 56293
rect 36266 56253 36278 56287
rect 36312 56253 36324 56287
rect 36266 56247 36324 56253
rect 35710 56176 35716 56228
rect 35768 56216 35774 56228
rect 36281 56216 36309 56247
rect 36354 56244 36360 56296
rect 36412 56284 36418 56296
rect 36449 56287 36507 56293
rect 36449 56284 36461 56287
rect 36412 56256 36461 56284
rect 36412 56244 36418 56256
rect 36449 56253 36461 56256
rect 36495 56253 36507 56287
rect 36449 56247 36507 56253
rect 36679 56287 36737 56293
rect 36679 56253 36691 56287
rect 36725 56284 36737 56287
rect 37826 56284 37832 56296
rect 36725 56256 37832 56284
rect 36725 56253 36737 56256
rect 36679 56247 36737 56253
rect 37826 56244 37832 56256
rect 37884 56244 37890 56296
rect 36538 56216 36544 56228
rect 35768 56188 36309 56216
rect 36499 56188 36544 56216
rect 35768 56176 35774 56188
rect 36538 56176 36544 56188
rect 36596 56176 36602 56228
rect 37369 56219 37427 56225
rect 37369 56185 37381 56219
rect 37415 56185 37427 56219
rect 37369 56179 37427 56185
rect 37384 56148 37412 56179
rect 39390 56148 39396 56160
rect 34164 56120 39396 56148
rect 8444 56108 8450 56120
rect 39390 56108 39396 56120
rect 39448 56108 39454 56160
rect 1104 56058 38824 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 38824 56058
rect 1104 55984 38824 56006
rect 26878 55904 26884 55956
rect 26936 55944 26942 55956
rect 28626 55944 28632 55956
rect 26936 55916 28632 55944
rect 26936 55904 26942 55916
rect 28626 55904 28632 55916
rect 28684 55904 28690 55956
rect 35621 55947 35679 55953
rect 35621 55913 35633 55947
rect 35667 55944 35679 55947
rect 36262 55944 36268 55956
rect 35667 55916 36268 55944
rect 35667 55913 35679 55916
rect 35621 55907 35679 55913
rect 36262 55904 36268 55916
rect 36320 55944 36326 55956
rect 38930 55944 38936 55956
rect 36320 55916 36492 55944
rect 36320 55904 36326 55916
rect 6730 55836 6736 55888
rect 6788 55876 6794 55888
rect 17126 55876 17132 55888
rect 6788 55848 17132 55876
rect 6788 55836 6794 55848
rect 17126 55836 17132 55848
rect 17184 55836 17190 55888
rect 33318 55836 33324 55888
rect 33376 55876 33382 55888
rect 33502 55876 33508 55888
rect 33376 55848 33508 55876
rect 33376 55836 33382 55848
rect 33502 55836 33508 55848
rect 33560 55836 33566 55888
rect 34054 55836 34060 55888
rect 34112 55876 34118 55888
rect 35250 55876 35256 55888
rect 34112 55848 35256 55876
rect 34112 55836 34118 55848
rect 35250 55836 35256 55848
rect 35308 55836 35314 55888
rect 36464 55885 36492 55916
rect 36729 55916 38936 55944
rect 36449 55879 36507 55885
rect 36449 55845 36461 55879
rect 36495 55845 36507 55879
rect 36449 55839 36507 55845
rect 1394 55808 1400 55820
rect 1355 55780 1400 55808
rect 1394 55768 1400 55780
rect 1452 55768 1458 55820
rect 34793 55811 34851 55817
rect 34793 55777 34805 55811
rect 34839 55808 34851 55811
rect 34882 55808 34888 55820
rect 34839 55780 34888 55808
rect 34839 55777 34851 55780
rect 34793 55771 34851 55777
rect 34882 55768 34888 55780
rect 34940 55768 34946 55820
rect 35529 55811 35587 55817
rect 35529 55777 35541 55811
rect 35575 55777 35587 55811
rect 35529 55771 35587 55777
rect 36173 55811 36231 55817
rect 36173 55777 36185 55811
rect 36219 55777 36231 55811
rect 36173 55771 36231 55777
rect 1578 55700 1584 55752
rect 1636 55740 1642 55752
rect 6454 55740 6460 55752
rect 1636 55712 6460 55740
rect 1636 55700 1642 55712
rect 6454 55700 6460 55712
rect 6512 55700 6518 55752
rect 21910 55700 21916 55752
rect 21968 55740 21974 55752
rect 35544 55740 35572 55771
rect 21968 55712 35572 55740
rect 36188 55740 36216 55771
rect 36262 55768 36268 55820
rect 36320 55808 36326 55820
rect 36538 55808 36544 55820
rect 36320 55780 36365 55808
rect 36499 55780 36544 55808
rect 36320 55768 36326 55780
rect 36538 55768 36544 55780
rect 36596 55768 36602 55820
rect 36729 55817 36757 55916
rect 38930 55904 38936 55916
rect 38988 55904 38994 55956
rect 36679 55811 36757 55817
rect 36679 55777 36691 55811
rect 36725 55780 36757 55811
rect 36725 55777 36737 55780
rect 36679 55771 36737 55777
rect 36814 55768 36820 55820
rect 36872 55768 36878 55820
rect 36832 55740 36860 55768
rect 36188 55712 36860 55740
rect 21968 55700 21974 55712
rect 28994 55632 29000 55684
rect 29052 55672 29058 55684
rect 36817 55675 36875 55681
rect 36817 55672 36829 55675
rect 29052 55644 36829 55672
rect 29052 55632 29058 55644
rect 36817 55641 36829 55644
rect 36863 55641 36875 55675
rect 36817 55635 36875 55641
rect 1581 55607 1639 55613
rect 1581 55573 1593 55607
rect 1627 55604 1639 55607
rect 4890 55604 4896 55616
rect 1627 55576 4896 55604
rect 1627 55573 1639 55576
rect 1581 55567 1639 55573
rect 4890 55564 4896 55576
rect 4948 55564 4954 55616
rect 34977 55607 35035 55613
rect 34977 55573 34989 55607
rect 35023 55604 35035 55607
rect 35250 55604 35256 55616
rect 35023 55576 35256 55604
rect 35023 55573 35035 55576
rect 34977 55567 35035 55573
rect 35250 55564 35256 55576
rect 35308 55564 35314 55616
rect 1104 55514 38824 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 38824 55514
rect 1104 55440 38824 55462
rect 28626 55360 28632 55412
rect 28684 55400 28690 55412
rect 29181 55403 29239 55409
rect 29181 55400 29193 55403
rect 28684 55372 29193 55400
rect 28684 55360 28690 55372
rect 29181 55369 29193 55372
rect 29227 55369 29239 55403
rect 29181 55363 29239 55369
rect 36446 55360 36452 55412
rect 36504 55400 36510 55412
rect 36504 55372 36952 55400
rect 36504 55360 36510 55372
rect 36924 55344 36952 55372
rect 20070 55292 20076 55344
rect 20128 55332 20134 55344
rect 22094 55332 22100 55344
rect 20128 55304 22100 55332
rect 20128 55292 20134 55304
rect 22094 55292 22100 55304
rect 22152 55292 22158 55344
rect 36354 55292 36360 55344
rect 36412 55332 36418 55344
rect 36412 55304 36584 55332
rect 36412 55292 36418 55304
rect 35710 55224 35716 55276
rect 35768 55264 35774 55276
rect 36446 55264 36452 55276
rect 35768 55236 36452 55264
rect 35768 55224 35774 55236
rect 36446 55224 36452 55236
rect 36504 55224 36510 55276
rect 36556 55264 36584 55304
rect 36906 55292 36912 55344
rect 36964 55292 36970 55344
rect 37182 55264 37188 55276
rect 36556 55236 37188 55264
rect 1394 55196 1400 55208
rect 1355 55168 1400 55196
rect 1394 55156 1400 55168
rect 1452 55156 1458 55208
rect 29086 55196 29092 55208
rect 29047 55168 29092 55196
rect 29086 55156 29092 55168
rect 29144 55156 29150 55208
rect 34609 55199 34667 55205
rect 34609 55165 34621 55199
rect 34655 55196 34667 55199
rect 35434 55196 35440 55208
rect 34655 55168 35440 55196
rect 34655 55165 34667 55168
rect 34609 55159 34667 55165
rect 35434 55156 35440 55168
rect 35492 55156 35498 55208
rect 35986 55156 35992 55208
rect 36044 55196 36050 55208
rect 36354 55205 36360 55208
rect 36173 55199 36231 55205
rect 36173 55196 36185 55199
rect 36044 55168 36185 55196
rect 36044 55156 36050 55168
rect 36173 55165 36185 55168
rect 36219 55165 36231 55199
rect 36173 55159 36231 55165
rect 36321 55199 36360 55205
rect 36321 55165 36333 55199
rect 36321 55159 36360 55165
rect 36354 55156 36360 55159
rect 36412 55156 36418 55208
rect 36556 55196 36584 55236
rect 37182 55224 37188 55236
rect 37240 55224 37246 55276
rect 37752 55236 38056 55264
rect 36464 55168 36584 55196
rect 36679 55199 36737 55205
rect 20622 55088 20628 55140
rect 20680 55128 20686 55140
rect 22278 55128 22284 55140
rect 20680 55100 22284 55128
rect 20680 55088 20686 55100
rect 22278 55088 22284 55100
rect 22336 55088 22342 55140
rect 36464 55137 36492 55168
rect 36679 55165 36691 55199
rect 36725 55196 36737 55199
rect 37366 55196 37372 55208
rect 36725 55168 37372 55196
rect 36725 55165 36737 55168
rect 36679 55159 36737 55165
rect 37366 55156 37372 55168
rect 37424 55156 37430 55208
rect 37553 55199 37611 55205
rect 37553 55165 37565 55199
rect 37599 55196 37611 55199
rect 37752 55196 37780 55236
rect 37918 55196 37924 55208
rect 37599 55168 37780 55196
rect 37879 55168 37924 55196
rect 37599 55165 37611 55168
rect 37553 55159 37611 55165
rect 37918 55156 37924 55168
rect 37976 55156 37982 55208
rect 38028 55196 38056 55236
rect 39298 55196 39304 55208
rect 38028 55168 39304 55196
rect 39298 55156 39304 55168
rect 39356 55156 39362 55208
rect 36449 55131 36507 55137
rect 36449 55097 36461 55131
rect 36495 55097 36507 55131
rect 36449 55091 36507 55097
rect 36538 55088 36544 55140
rect 36596 55128 36602 55140
rect 37734 55128 37740 55140
rect 36596 55100 36641 55128
rect 37695 55100 37740 55128
rect 36596 55088 36602 55100
rect 37734 55088 37740 55100
rect 37792 55088 37798 55140
rect 37826 55088 37832 55140
rect 37884 55128 37890 55140
rect 37884 55100 37929 55128
rect 37884 55088 37890 55100
rect 1578 55060 1584 55072
rect 1539 55032 1584 55060
rect 1578 55020 1584 55032
rect 1636 55020 1642 55072
rect 34793 55063 34851 55069
rect 34793 55029 34805 55063
rect 34839 55060 34851 55063
rect 35158 55060 35164 55072
rect 34839 55032 35164 55060
rect 34839 55029 34851 55032
rect 34793 55023 34851 55029
rect 35158 55020 35164 55032
rect 35216 55020 35222 55072
rect 35434 55020 35440 55072
rect 35492 55060 35498 55072
rect 36817 55063 36875 55069
rect 36817 55060 36829 55063
rect 35492 55032 36829 55060
rect 35492 55020 35498 55032
rect 36817 55029 36829 55032
rect 36863 55029 36875 55063
rect 36817 55023 36875 55029
rect 37458 55020 37464 55072
rect 37516 55060 37522 55072
rect 38105 55063 38163 55069
rect 38105 55060 38117 55063
rect 37516 55032 38117 55060
rect 37516 55020 37522 55032
rect 38105 55029 38117 55032
rect 38151 55029 38163 55063
rect 38105 55023 38163 55029
rect 1104 54970 38824 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 38824 54970
rect 1104 54896 38824 54918
rect 19978 54816 19984 54868
rect 20036 54856 20042 54868
rect 20622 54856 20628 54868
rect 20036 54828 20628 54856
rect 20036 54816 20042 54828
rect 20622 54816 20628 54828
rect 20680 54816 20686 54868
rect 34330 54816 34336 54868
rect 34388 54856 34394 54868
rect 35713 54859 35771 54865
rect 35713 54856 35725 54859
rect 34388 54828 35725 54856
rect 34388 54816 34394 54828
rect 35713 54825 35725 54828
rect 35759 54825 35771 54859
rect 35713 54819 35771 54825
rect 36449 54791 36507 54797
rect 36188 54760 36400 54788
rect 35529 54723 35587 54729
rect 35529 54689 35541 54723
rect 35575 54720 35587 54723
rect 35710 54720 35716 54732
rect 35575 54692 35716 54720
rect 35575 54689 35587 54692
rect 35529 54683 35587 54689
rect 35710 54680 35716 54692
rect 35768 54680 35774 54732
rect 36188 54729 36216 54760
rect 36173 54723 36231 54729
rect 36173 54689 36185 54723
rect 36219 54689 36231 54723
rect 36173 54683 36231 54689
rect 36266 54723 36324 54729
rect 36266 54689 36278 54723
rect 36312 54689 36324 54723
rect 36266 54683 36324 54689
rect 35986 54612 35992 54664
rect 36044 54652 36050 54664
rect 36280 54652 36308 54683
rect 36044 54624 36308 54652
rect 36372 54652 36400 54760
rect 36449 54757 36461 54791
rect 36495 54788 36507 54791
rect 37182 54788 37188 54800
rect 36495 54760 37188 54788
rect 36495 54757 36507 54760
rect 36449 54751 36507 54757
rect 37182 54748 37188 54760
rect 37240 54748 37246 54800
rect 36538 54720 36544 54732
rect 36499 54692 36544 54720
rect 36538 54680 36544 54692
rect 36596 54680 36602 54732
rect 36679 54723 36737 54729
rect 36679 54689 36691 54723
rect 36725 54720 36737 54723
rect 38194 54720 38200 54732
rect 36725 54692 38200 54720
rect 36725 54689 36737 54692
rect 36679 54683 36737 54689
rect 38194 54680 38200 54692
rect 38252 54680 38258 54732
rect 37550 54652 37556 54664
rect 36372 54624 37556 54652
rect 36044 54612 36050 54624
rect 37550 54612 37556 54624
rect 37608 54612 37614 54664
rect 21266 54584 21272 54596
rect 12406 54556 21272 54584
rect 2866 54476 2872 54528
rect 2924 54516 2930 54528
rect 12406 54516 12434 54556
rect 21266 54544 21272 54556
rect 21324 54544 21330 54596
rect 35158 54544 35164 54596
rect 35216 54584 35222 54596
rect 38930 54584 38936 54596
rect 35216 54556 38936 54584
rect 35216 54544 35222 54556
rect 38930 54544 38936 54556
rect 38988 54544 38994 54596
rect 2924 54488 12434 54516
rect 2924 54476 2930 54488
rect 24578 54476 24584 54528
rect 24636 54516 24642 54528
rect 32674 54516 32680 54528
rect 24636 54488 32680 54516
rect 24636 54476 24642 54488
rect 32674 54476 32680 54488
rect 32732 54476 32738 54528
rect 33042 54476 33048 54528
rect 33100 54516 33106 54528
rect 36817 54519 36875 54525
rect 36817 54516 36829 54519
rect 33100 54488 36829 54516
rect 33100 54476 33106 54488
rect 36817 54485 36829 54488
rect 36863 54485 36875 54519
rect 36817 54479 36875 54485
rect 1104 54426 38824 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 38824 54426
rect 1104 54352 38824 54374
rect 36262 54312 36268 54324
rect 36223 54284 36268 54312
rect 36262 54272 36268 54284
rect 36320 54272 36326 54324
rect 35894 54204 35900 54256
rect 35952 54244 35958 54256
rect 36909 54247 36967 54253
rect 36909 54244 36921 54247
rect 35952 54216 36921 54244
rect 35952 54204 35958 54216
rect 36909 54213 36921 54216
rect 36955 54213 36967 54247
rect 36909 54207 36967 54213
rect 39022 54176 39028 54188
rect 37568 54148 39028 54176
rect 1394 54108 1400 54120
rect 1355 54080 1400 54108
rect 1394 54068 1400 54080
rect 1452 54068 1458 54120
rect 25590 54068 25596 54120
rect 25648 54108 25654 54120
rect 31386 54108 31392 54120
rect 25648 54080 31392 54108
rect 25648 54068 25654 54080
rect 31386 54068 31392 54080
rect 31444 54068 31450 54120
rect 35802 54068 35808 54120
rect 35860 54108 35866 54120
rect 36449 54111 36507 54117
rect 36449 54108 36461 54111
rect 35860 54080 36461 54108
rect 35860 54068 35866 54080
rect 36449 54077 36461 54080
rect 36495 54077 36507 54111
rect 37090 54108 37096 54120
rect 37051 54080 37096 54108
rect 36449 54071 36507 54077
rect 37090 54068 37096 54080
rect 37148 54068 37154 54120
rect 37568 54117 37596 54148
rect 39022 54136 39028 54148
rect 39080 54136 39086 54188
rect 37553 54111 37611 54117
rect 37553 54077 37565 54111
rect 37599 54077 37611 54111
rect 37553 54071 37611 54077
rect 37921 54111 37979 54117
rect 37921 54077 37933 54111
rect 37967 54108 37979 54111
rect 38194 54108 38200 54120
rect 37967 54080 38200 54108
rect 37967 54077 37979 54080
rect 37921 54071 37979 54077
rect 38194 54068 38200 54080
rect 38252 54068 38258 54120
rect 36262 54000 36268 54052
rect 36320 54040 36326 54052
rect 36906 54040 36912 54052
rect 36320 54012 36912 54040
rect 36320 54000 36326 54012
rect 36906 54000 36912 54012
rect 36964 54000 36970 54052
rect 37734 54040 37740 54052
rect 37695 54012 37740 54040
rect 37734 54000 37740 54012
rect 37792 54000 37798 54052
rect 37826 54000 37832 54052
rect 37884 54040 37890 54052
rect 37884 54012 37929 54040
rect 37884 54000 37890 54012
rect 1581 53975 1639 53981
rect 1581 53941 1593 53975
rect 1627 53972 1639 53975
rect 1946 53972 1952 53984
rect 1627 53944 1952 53972
rect 1627 53941 1639 53944
rect 1581 53935 1639 53941
rect 1946 53932 1952 53944
rect 2004 53932 2010 53984
rect 35434 53932 35440 53984
rect 35492 53972 35498 53984
rect 35710 53972 35716 53984
rect 35492 53944 35716 53972
rect 35492 53932 35498 53944
rect 35710 53932 35716 53944
rect 35768 53932 35774 53984
rect 35894 53932 35900 53984
rect 35952 53972 35958 53984
rect 37182 53972 37188 53984
rect 35952 53944 37188 53972
rect 35952 53932 35958 53944
rect 37182 53932 37188 53944
rect 37240 53932 37246 53984
rect 37550 53932 37556 53984
rect 37608 53972 37614 53984
rect 38105 53975 38163 53981
rect 38105 53972 38117 53975
rect 37608 53944 38117 53972
rect 37608 53932 37614 53944
rect 38105 53941 38117 53944
rect 38151 53941 38163 53975
rect 38105 53935 38163 53941
rect 1104 53882 38824 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 38824 53882
rect 1104 53808 38824 53830
rect 31754 53728 31760 53780
rect 31812 53768 31818 53780
rect 33962 53768 33968 53780
rect 31812 53740 33968 53768
rect 31812 53728 31818 53740
rect 33962 53728 33968 53740
rect 34020 53728 34026 53780
rect 36446 53728 36452 53780
rect 36504 53768 36510 53780
rect 36541 53771 36599 53777
rect 36541 53768 36553 53771
rect 36504 53740 36553 53768
rect 36504 53728 36510 53740
rect 36541 53737 36553 53740
rect 36587 53737 36599 53771
rect 36541 53731 36599 53737
rect 36722 53728 36728 53780
rect 36780 53768 36786 53780
rect 37185 53771 37243 53777
rect 37185 53768 37197 53771
rect 36780 53740 37197 53768
rect 36780 53728 36786 53740
rect 37185 53737 37197 53740
rect 37231 53737 37243 53771
rect 37185 53731 37243 53737
rect 1394 53632 1400 53644
rect 1355 53604 1400 53632
rect 1394 53592 1400 53604
rect 1452 53592 1458 53644
rect 36722 53632 36728 53644
rect 36683 53604 36728 53632
rect 36722 53592 36728 53604
rect 36780 53592 36786 53644
rect 37366 53632 37372 53644
rect 37327 53604 37372 53632
rect 37366 53592 37372 53604
rect 37424 53592 37430 53644
rect 1581 53431 1639 53437
rect 1581 53397 1593 53431
rect 1627 53428 1639 53431
rect 7926 53428 7932 53440
rect 1627 53400 7932 53428
rect 1627 53397 1639 53400
rect 1581 53391 1639 53397
rect 7926 53388 7932 53400
rect 7984 53388 7990 53440
rect 1104 53338 38824 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 38824 53338
rect 1104 53264 38824 53286
rect 27065 53227 27123 53233
rect 27065 53193 27077 53227
rect 27111 53224 27123 53227
rect 27154 53224 27160 53236
rect 27111 53196 27160 53224
rect 27111 53193 27123 53196
rect 27065 53187 27123 53193
rect 27154 53184 27160 53196
rect 27212 53184 27218 53236
rect 28966 53196 37596 53224
rect 24210 53116 24216 53168
rect 24268 53156 24274 53168
rect 28966 53156 28994 53196
rect 24268 53128 28994 53156
rect 24268 53116 24274 53128
rect 34698 53116 34704 53168
rect 34756 53156 34762 53168
rect 36081 53159 36139 53165
rect 36081 53156 36093 53159
rect 34756 53128 36093 53156
rect 34756 53116 34762 53128
rect 36081 53125 36093 53128
rect 36127 53125 36139 53159
rect 36081 53119 36139 53125
rect 3418 53048 3424 53100
rect 3476 53088 3482 53100
rect 9950 53088 9956 53100
rect 3476 53060 9956 53088
rect 3476 53048 3482 53060
rect 9950 53048 9956 53060
rect 10008 53048 10014 53100
rect 35434 53088 35440 53100
rect 26528 53060 35440 53088
rect 26528 53029 26556 53060
rect 35434 53048 35440 53060
rect 35492 53048 35498 53100
rect 26513 53023 26571 53029
rect 26513 52989 26525 53023
rect 26559 52989 26571 53023
rect 26886 53023 26944 53029
rect 26886 53020 26898 53023
rect 26513 52983 26571 52989
rect 26620 52992 26898 53020
rect 8018 52912 8024 52964
rect 8076 52952 8082 52964
rect 26620 52952 26648 52992
rect 26886 52989 26898 52992
rect 26932 52989 26944 53023
rect 26886 52983 26944 52989
rect 34054 52980 34060 53032
rect 34112 53020 34118 53032
rect 34698 53020 34704 53032
rect 34112 52992 34704 53020
rect 34112 52980 34118 52992
rect 34698 52980 34704 52992
rect 34756 52980 34762 53032
rect 35802 52980 35808 53032
rect 35860 53020 35866 53032
rect 35897 53023 35955 53029
rect 35897 53020 35909 53023
rect 35860 52992 35909 53020
rect 35860 52980 35866 52992
rect 35897 52989 35909 52992
rect 35943 52989 35955 53023
rect 35897 52983 35955 52989
rect 36541 53023 36599 53029
rect 36541 52989 36553 53023
rect 36587 53020 36599 53023
rect 36630 53020 36636 53032
rect 36587 52992 36636 53020
rect 36587 52989 36599 52992
rect 36541 52983 36599 52989
rect 36630 52980 36636 52992
rect 36688 52980 36694 53032
rect 36906 53020 36912 53032
rect 36867 52992 36912 53020
rect 36906 52980 36912 52992
rect 36964 52980 36970 53032
rect 37568 53029 37596 53196
rect 37553 53023 37611 53029
rect 37553 52989 37565 53023
rect 37599 52989 37611 53023
rect 37734 53020 37740 53032
rect 37695 52992 37740 53020
rect 37553 52983 37611 52989
rect 37734 52980 37740 52992
rect 37792 52980 37798 53032
rect 37921 53023 37979 53029
rect 37921 52989 37933 53023
rect 37967 53020 37979 53023
rect 38102 53020 38108 53032
rect 37967 52992 38108 53020
rect 37967 52989 37979 52992
rect 37921 52983 37979 52989
rect 38102 52980 38108 52992
rect 38160 52980 38166 53032
rect 8076 52924 26648 52952
rect 26697 52955 26755 52961
rect 8076 52912 8082 52924
rect 26697 52921 26709 52955
rect 26743 52921 26755 52955
rect 26697 52915 26755 52921
rect 26326 52844 26332 52896
rect 26384 52884 26390 52896
rect 26712 52884 26740 52915
rect 26786 52912 26792 52964
rect 26844 52952 26850 52964
rect 36722 52952 36728 52964
rect 26844 52924 26889 52952
rect 36683 52924 36728 52952
rect 26844 52912 26850 52924
rect 36722 52912 36728 52924
rect 36780 52912 36786 52964
rect 36817 52955 36875 52961
rect 36817 52921 36829 52955
rect 36863 52952 36875 52955
rect 37826 52952 37832 52964
rect 36863 52924 37832 52952
rect 36863 52921 36875 52924
rect 36817 52915 36875 52921
rect 37826 52912 37832 52924
rect 37884 52912 37890 52964
rect 26384 52856 26740 52884
rect 26384 52844 26390 52856
rect 36630 52844 36636 52896
rect 36688 52884 36694 52896
rect 37093 52887 37151 52893
rect 37093 52884 37105 52887
rect 36688 52856 37105 52884
rect 36688 52844 36694 52856
rect 37093 52853 37105 52856
rect 37139 52853 37151 52887
rect 37093 52847 37151 52853
rect 37182 52844 37188 52896
rect 37240 52884 37246 52896
rect 38105 52887 38163 52893
rect 38105 52884 38117 52887
rect 37240 52856 38117 52884
rect 37240 52844 37246 52856
rect 38105 52853 38117 52856
rect 38151 52853 38163 52887
rect 38105 52847 38163 52853
rect 1104 52794 38824 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 38824 52794
rect 1104 52720 38824 52742
rect 36354 52640 36360 52692
rect 36412 52680 36418 52692
rect 36541 52683 36599 52689
rect 36541 52680 36553 52683
rect 36412 52652 36553 52680
rect 36412 52640 36418 52652
rect 36541 52649 36553 52652
rect 36587 52649 36599 52683
rect 36541 52643 36599 52649
rect 36814 52640 36820 52692
rect 36872 52680 36878 52692
rect 37185 52683 37243 52689
rect 37185 52680 37197 52683
rect 36872 52652 37197 52680
rect 36872 52640 36878 52652
rect 37185 52649 37197 52652
rect 37231 52649 37243 52683
rect 37185 52643 37243 52649
rect 1854 52544 1860 52556
rect 1815 52516 1860 52544
rect 1854 52504 1860 52516
rect 1912 52504 1918 52556
rect 7834 52504 7840 52556
rect 7892 52544 7898 52556
rect 8754 52544 8760 52556
rect 7892 52516 8760 52544
rect 7892 52504 7898 52516
rect 8754 52504 8760 52516
rect 8812 52504 8818 52556
rect 20162 52504 20168 52556
rect 20220 52544 20226 52556
rect 28534 52544 28540 52556
rect 20220 52516 28540 52544
rect 20220 52504 20226 52516
rect 28534 52504 28540 52516
rect 28592 52504 28598 52556
rect 36722 52544 36728 52556
rect 36683 52516 36728 52544
rect 36722 52504 36728 52516
rect 36780 52504 36786 52556
rect 37182 52504 37188 52556
rect 37240 52544 37246 52556
rect 37369 52547 37427 52553
rect 37369 52544 37381 52547
rect 37240 52516 37381 52544
rect 37240 52504 37246 52516
rect 37369 52513 37381 52516
rect 37415 52513 37427 52547
rect 37369 52507 37427 52513
rect 2041 52479 2099 52485
rect 2041 52445 2053 52479
rect 2087 52476 2099 52479
rect 18046 52476 18052 52488
rect 2087 52448 18052 52476
rect 2087 52445 2099 52448
rect 2041 52439 2099 52445
rect 18046 52436 18052 52448
rect 18104 52436 18110 52488
rect 34514 52368 34520 52420
rect 34572 52408 34578 52420
rect 36814 52408 36820 52420
rect 34572 52380 36820 52408
rect 34572 52368 34578 52380
rect 36814 52368 36820 52380
rect 36872 52368 36878 52420
rect 21726 52300 21732 52352
rect 21784 52340 21790 52352
rect 27154 52340 27160 52352
rect 21784 52312 27160 52340
rect 21784 52300 21790 52312
rect 27154 52300 27160 52312
rect 27212 52300 27218 52352
rect 1104 52250 38824 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 38824 52250
rect 1104 52176 38824 52198
rect 21726 52096 21732 52148
rect 21784 52136 21790 52148
rect 28810 52136 28816 52148
rect 21784 52108 28816 52136
rect 21784 52096 21790 52108
rect 28810 52096 28816 52108
rect 28868 52096 28874 52148
rect 2041 52071 2099 52077
rect 2041 52037 2053 52071
rect 2087 52068 2099 52071
rect 8294 52068 8300 52080
rect 2087 52040 8300 52068
rect 2087 52037 2099 52040
rect 2041 52031 2099 52037
rect 8294 52028 8300 52040
rect 8352 52028 8358 52080
rect 27065 52071 27123 52077
rect 27065 52037 27077 52071
rect 27111 52068 27123 52071
rect 27522 52068 27528 52080
rect 27111 52040 27528 52068
rect 27111 52037 27123 52040
rect 27065 52031 27123 52037
rect 27522 52028 27528 52040
rect 27580 52028 27586 52080
rect 34330 52000 34336 52012
rect 26528 51972 34336 52000
rect 26528 51941 26556 51972
rect 34330 51960 34336 51972
rect 34388 51960 34394 52012
rect 26513 51935 26571 51941
rect 26513 51901 26525 51935
rect 26559 51901 26571 51935
rect 26786 51932 26792 51944
rect 26747 51904 26792 51932
rect 26513 51895 26571 51901
rect 26786 51892 26792 51904
rect 26844 51892 26850 51944
rect 26886 51935 26944 51941
rect 26886 51901 26898 51935
rect 26932 51901 26944 51935
rect 26886 51895 26944 51901
rect 1854 51864 1860 51876
rect 1815 51836 1860 51864
rect 1854 51824 1860 51836
rect 1912 51824 1918 51876
rect 26326 51824 26332 51876
rect 26384 51864 26390 51876
rect 26697 51867 26755 51873
rect 26697 51864 26709 51867
rect 26384 51836 26709 51864
rect 26384 51824 26390 51836
rect 26697 51833 26709 51836
rect 26743 51833 26755 51867
rect 26697 51827 26755 51833
rect 22186 51756 22192 51808
rect 22244 51796 22250 51808
rect 26896 51796 26924 51895
rect 27154 51892 27160 51944
rect 27212 51932 27218 51944
rect 37553 51935 37611 51941
rect 37553 51932 37565 51935
rect 27212 51904 37565 51932
rect 27212 51892 27218 51904
rect 37553 51901 37565 51904
rect 37599 51901 37611 51935
rect 37553 51895 37611 51901
rect 37921 51935 37979 51941
rect 37921 51901 37933 51935
rect 37967 51932 37979 51935
rect 39022 51932 39028 51944
rect 37967 51904 39028 51932
rect 37967 51901 37979 51904
rect 37921 51895 37979 51901
rect 39022 51892 39028 51904
rect 39080 51892 39086 51944
rect 37734 51864 37740 51876
rect 37695 51836 37740 51864
rect 37734 51824 37740 51836
rect 37792 51824 37798 51876
rect 37826 51824 37832 51876
rect 37884 51864 37890 51876
rect 37884 51836 37929 51864
rect 37884 51824 37890 51836
rect 22244 51768 26924 51796
rect 22244 51756 22250 51768
rect 36446 51756 36452 51808
rect 36504 51796 36510 51808
rect 38105 51799 38163 51805
rect 38105 51796 38117 51799
rect 36504 51768 38117 51796
rect 36504 51756 36510 51768
rect 38105 51765 38117 51768
rect 38151 51765 38163 51799
rect 38105 51759 38163 51765
rect 1104 51706 38824 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 38824 51706
rect 1104 51632 38824 51654
rect 19797 51595 19855 51601
rect 19797 51561 19809 51595
rect 19843 51592 19855 51595
rect 21542 51592 21548 51604
rect 19843 51564 21548 51592
rect 19843 51561 19855 51564
rect 19797 51555 19855 51561
rect 21542 51552 21548 51564
rect 21600 51552 21606 51604
rect 22462 51552 22468 51604
rect 22520 51592 22526 51604
rect 23109 51595 23167 51601
rect 23109 51592 23121 51595
rect 22520 51564 23121 51592
rect 22520 51552 22526 51564
rect 23109 51561 23121 51564
rect 23155 51561 23167 51595
rect 24946 51592 24952 51604
rect 24907 51564 24952 51592
rect 23109 51555 23167 51561
rect 24946 51552 24952 51564
rect 25004 51552 25010 51604
rect 27522 51592 27528 51604
rect 26436 51564 27528 51592
rect 7650 51484 7656 51536
rect 7708 51524 7714 51536
rect 7708 51496 26372 51524
rect 7708 51484 7714 51496
rect 19521 51459 19579 51465
rect 19521 51456 19533 51459
rect 6886 51428 19533 51456
rect 3418 51348 3424 51400
rect 3476 51388 3482 51400
rect 6886 51388 6914 51428
rect 19521 51425 19533 51428
rect 19567 51425 19579 51459
rect 19521 51419 19579 51425
rect 21266 51416 21272 51468
rect 21324 51456 21330 51468
rect 23017 51459 23075 51465
rect 23017 51456 23029 51459
rect 21324 51428 23029 51456
rect 21324 51416 21330 51428
rect 23017 51425 23029 51428
rect 23063 51425 23075 51459
rect 23017 51419 23075 51425
rect 24673 51459 24731 51465
rect 24673 51425 24685 51459
rect 24719 51425 24731 51459
rect 24673 51419 24731 51425
rect 26237 51459 26295 51465
rect 26237 51425 26249 51459
rect 26283 51425 26295 51459
rect 26237 51419 26295 51425
rect 3476 51360 6914 51388
rect 3476 51348 3482 51360
rect 11054 51280 11060 51332
rect 11112 51320 11118 51332
rect 24688 51320 24716 51419
rect 11112 51292 24716 51320
rect 26252 51320 26280 51419
rect 26344 51388 26372 51496
rect 26436 51465 26464 51564
rect 27522 51552 27528 51564
rect 27580 51552 27586 51604
rect 29086 51552 29092 51604
rect 29144 51552 29150 51604
rect 29178 51552 29184 51604
rect 29236 51592 29242 51604
rect 29825 51595 29883 51601
rect 29825 51592 29837 51595
rect 29236 51564 29837 51592
rect 29236 51552 29242 51564
rect 29825 51561 29837 51564
rect 29871 51561 29883 51595
rect 29825 51555 29883 51561
rect 35986 51552 35992 51604
rect 36044 51592 36050 51604
rect 37185 51595 37243 51601
rect 37185 51592 37197 51595
rect 36044 51564 37197 51592
rect 36044 51552 36050 51564
rect 37185 51561 37197 51564
rect 37231 51561 37243 51595
rect 37185 51555 37243 51561
rect 26513 51527 26571 51533
rect 26513 51493 26525 51527
rect 26559 51524 26571 51527
rect 26786 51524 26792 51536
rect 26559 51496 26792 51524
rect 26559 51493 26571 51496
rect 26513 51487 26571 51493
rect 26786 51484 26792 51496
rect 26844 51484 26850 51536
rect 28810 51524 28816 51536
rect 28771 51496 28816 51524
rect 28810 51484 28816 51496
rect 28868 51484 28874 51536
rect 26421 51459 26479 51465
rect 26421 51425 26433 51459
rect 26467 51425 26479 51459
rect 26610 51459 26668 51465
rect 26610 51456 26622 51459
rect 26421 51419 26479 51425
rect 26528 51428 26622 51456
rect 26528 51388 26556 51428
rect 26610 51425 26622 51428
rect 26656 51425 26668 51459
rect 26610 51419 26668 51425
rect 27893 51459 27951 51465
rect 27893 51425 27905 51459
rect 27939 51456 27951 51459
rect 28534 51456 28540 51468
rect 27939 51428 28540 51456
rect 27939 51425 27951 51428
rect 27893 51419 27951 51425
rect 28534 51416 28540 51428
rect 28592 51416 28598 51468
rect 29104 51400 29132 51552
rect 30190 51524 30196 51536
rect 29196 51496 30196 51524
rect 29196 51465 29224 51496
rect 30190 51484 30196 51496
rect 30248 51484 30254 51536
rect 34977 51527 35035 51533
rect 34977 51493 34989 51527
rect 35023 51524 35035 51527
rect 35526 51524 35532 51536
rect 35023 51496 35532 51524
rect 35023 51493 35035 51496
rect 34977 51487 35035 51493
rect 35526 51484 35532 51496
rect 35584 51484 35590 51536
rect 29181 51459 29239 51465
rect 29181 51425 29193 51459
rect 29227 51425 29239 51459
rect 29181 51419 29239 51425
rect 29362 51416 29368 51468
rect 29420 51456 29426 51468
rect 29733 51459 29791 51465
rect 29733 51456 29745 51459
rect 29420 51428 29745 51456
rect 29420 51416 29426 51428
rect 29733 51425 29745 51428
rect 29779 51425 29791 51459
rect 34609 51459 34667 51465
rect 34609 51456 34621 51459
rect 29733 51419 29791 51425
rect 31726 51428 34621 51456
rect 26344 51360 26556 51388
rect 29086 51348 29092 51400
rect 29144 51348 29150 51400
rect 29546 51348 29552 51400
rect 29604 51388 29610 51400
rect 31726 51388 31754 51428
rect 34609 51425 34621 51428
rect 34655 51425 34667 51459
rect 36538 51456 36544 51468
rect 36499 51428 36544 51456
rect 34609 51419 34667 51425
rect 36538 51416 36544 51428
rect 36596 51416 36602 51468
rect 37366 51456 37372 51468
rect 37327 51428 37372 51456
rect 37366 51416 37372 51428
rect 37424 51416 37430 51468
rect 29604 51360 31754 51388
rect 29604 51348 29610 51360
rect 26252 51292 26556 51320
rect 11112 51280 11118 51292
rect 26528 51252 26556 51292
rect 26712 51292 31754 51320
rect 26712 51252 26740 51292
rect 26528 51224 26740 51252
rect 26789 51255 26847 51261
rect 26789 51221 26801 51255
rect 26835 51252 26847 51255
rect 27982 51252 27988 51264
rect 26835 51224 27988 51252
rect 26835 51221 26847 51224
rect 26789 51215 26847 51221
rect 27982 51212 27988 51224
rect 28040 51212 28046 51264
rect 28169 51255 28227 51261
rect 28169 51221 28181 51255
rect 28215 51252 28227 51255
rect 29730 51252 29736 51264
rect 28215 51224 29736 51252
rect 28215 51221 28227 51224
rect 28169 51215 28227 51221
rect 29730 51212 29736 51224
rect 29788 51212 29794 51264
rect 31726 51252 31754 51292
rect 36262 51280 36268 51332
rect 36320 51320 36326 51332
rect 36538 51320 36544 51332
rect 36320 51292 36544 51320
rect 36320 51280 36326 51292
rect 36538 51280 36544 51292
rect 36596 51280 36602 51332
rect 36725 51323 36783 51329
rect 36725 51289 36737 51323
rect 36771 51320 36783 51323
rect 36814 51320 36820 51332
rect 36771 51292 36820 51320
rect 36771 51289 36783 51292
rect 36725 51283 36783 51289
rect 36814 51280 36820 51292
rect 36872 51280 36878 51332
rect 33318 51252 33324 51264
rect 31726 51224 33324 51252
rect 33318 51212 33324 51224
rect 33376 51212 33382 51264
rect 1104 51162 38824 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 38824 51162
rect 1104 51088 38824 51110
rect 1670 51008 1676 51060
rect 1728 51048 1734 51060
rect 8294 51048 8300 51060
rect 1728 51020 8300 51048
rect 1728 51008 1734 51020
rect 8294 51008 8300 51020
rect 8352 51008 8358 51060
rect 20714 51048 20720 51060
rect 20675 51020 20720 51048
rect 20714 51008 20720 51020
rect 20772 51008 20778 51060
rect 22554 51048 22560 51060
rect 22515 51020 22560 51048
rect 22554 51008 22560 51020
rect 22612 51008 22618 51060
rect 23566 51048 23572 51060
rect 23527 51020 23572 51048
rect 23566 51008 23572 51020
rect 23624 51008 23630 51060
rect 25406 51048 25412 51060
rect 25367 51020 25412 51048
rect 25406 51008 25412 51020
rect 25464 51008 25470 51060
rect 27065 51051 27123 51057
rect 27065 51017 27077 51051
rect 27111 51048 27123 51051
rect 27706 51048 27712 51060
rect 27111 51020 27712 51048
rect 27111 51017 27123 51020
rect 27065 51011 27123 51017
rect 27706 51008 27712 51020
rect 27764 51008 27770 51060
rect 30837 51051 30895 51057
rect 30837 51017 30849 51051
rect 30883 51048 30895 51051
rect 31754 51048 31760 51060
rect 30883 51020 31760 51048
rect 30883 51017 30895 51020
rect 30837 51011 30895 51017
rect 31754 51008 31760 51020
rect 31812 51008 31818 51060
rect 32858 51048 32864 51060
rect 32819 51020 32864 51048
rect 32858 51008 32864 51020
rect 32916 51008 32922 51060
rect 36262 51008 36268 51060
rect 36320 51048 36326 51060
rect 36998 51048 37004 51060
rect 36320 51020 37004 51048
rect 36320 51008 36326 51020
rect 36998 51008 37004 51020
rect 37056 51008 37062 51060
rect 37921 51051 37979 51057
rect 37921 51017 37933 51051
rect 37967 51048 37979 51051
rect 38010 51048 38016 51060
rect 37967 51020 38016 51048
rect 37967 51017 37979 51020
rect 37921 51011 37979 51017
rect 38010 51008 38016 51020
rect 38068 51008 38074 51060
rect 2041 50983 2099 50989
rect 2041 50949 2053 50983
rect 2087 50980 2099 50983
rect 7006 50980 7012 50992
rect 2087 50952 7012 50980
rect 2087 50949 2099 50952
rect 2041 50943 2099 50949
rect 7006 50940 7012 50952
rect 7064 50940 7070 50992
rect 22462 50940 22468 50992
rect 22520 50980 22526 50992
rect 23014 50980 23020 50992
rect 22520 50952 23020 50980
rect 22520 50940 22526 50952
rect 23014 50940 23020 50952
rect 23072 50940 23078 50992
rect 24854 50940 24860 50992
rect 24912 50980 24918 50992
rect 24912 50952 27016 50980
rect 24912 50940 24918 50952
rect 6886 50884 26929 50912
rect 1854 50844 1860 50856
rect 1815 50816 1860 50844
rect 1854 50804 1860 50816
rect 1912 50804 1918 50856
rect 4062 50804 4068 50856
rect 4120 50844 4126 50856
rect 6886 50844 6914 50884
rect 4120 50816 6914 50844
rect 4120 50804 4126 50816
rect 21542 50804 21548 50856
rect 21600 50844 21606 50856
rect 23477 50847 23535 50853
rect 23477 50844 23489 50847
rect 21600 50816 23489 50844
rect 21600 50804 21606 50816
rect 23477 50813 23489 50816
rect 23523 50813 23535 50847
rect 26510 50844 26516 50856
rect 26471 50816 26516 50844
rect 23477 50807 23535 50813
rect 26510 50804 26516 50816
rect 26568 50804 26574 50856
rect 26901 50853 26929 50884
rect 26886 50847 26944 50853
rect 26886 50813 26898 50847
rect 26932 50813 26944 50847
rect 26988 50844 27016 50952
rect 34330 50940 34336 50992
rect 34388 50980 34394 50992
rect 35894 50980 35900 50992
rect 34388 50952 35900 50980
rect 34388 50940 34394 50952
rect 35894 50940 35900 50952
rect 35952 50940 35958 50992
rect 37274 50980 37280 50992
rect 36464 50952 37280 50980
rect 35526 50912 35532 50924
rect 28828 50884 35532 50912
rect 28261 50847 28319 50853
rect 28261 50844 28273 50847
rect 26988 50816 28273 50844
rect 26886 50807 26944 50813
rect 28261 50813 28273 50816
rect 28307 50813 28319 50847
rect 28261 50807 28319 50813
rect 28537 50847 28595 50853
rect 28537 50813 28549 50847
rect 28583 50844 28595 50847
rect 28626 50844 28632 50856
rect 28583 50816 28632 50844
rect 28583 50813 28595 50816
rect 28537 50807 28595 50813
rect 28626 50804 28632 50816
rect 28684 50804 28690 50856
rect 28828 50853 28856 50884
rect 35526 50872 35532 50884
rect 35584 50912 35590 50924
rect 36354 50912 36360 50924
rect 35584 50884 36360 50912
rect 35584 50872 35590 50884
rect 36354 50872 36360 50884
rect 36412 50872 36418 50924
rect 28813 50847 28871 50853
rect 28813 50813 28825 50847
rect 28859 50813 28871 50847
rect 28813 50807 28871 50813
rect 28905 50847 28963 50853
rect 28905 50813 28917 50847
rect 28951 50844 28963 50847
rect 36464 50844 36492 50952
rect 37274 50940 37280 50952
rect 37332 50940 37338 50992
rect 37458 50912 37464 50924
rect 36740 50884 37464 50912
rect 36740 50853 36768 50884
rect 37458 50872 37464 50884
rect 37516 50872 37522 50924
rect 38746 50912 38752 50924
rect 37936 50884 38752 50912
rect 28951 50816 36492 50844
rect 36725 50847 36783 50853
rect 28951 50813 28963 50816
rect 28905 50807 28963 50813
rect 36725 50813 36737 50847
rect 36771 50813 36783 50847
rect 36725 50807 36783 50813
rect 36814 50804 36820 50856
rect 36872 50844 36878 50856
rect 37001 50847 37059 50853
rect 36872 50816 36917 50844
rect 36872 50804 36878 50816
rect 37001 50813 37013 50847
rect 37047 50813 37059 50847
rect 37001 50807 37059 50813
rect 37229 50847 37287 50853
rect 37229 50813 37241 50847
rect 37275 50844 37287 50847
rect 37936 50844 37964 50884
rect 38746 50872 38752 50884
rect 38804 50872 38810 50924
rect 38102 50844 38108 50856
rect 37275 50816 37964 50844
rect 38063 50816 38108 50844
rect 37275 50813 37287 50816
rect 37229 50807 37287 50813
rect 4614 50736 4620 50788
rect 4672 50776 4678 50788
rect 20441 50779 20499 50785
rect 20441 50776 20453 50779
rect 4672 50748 20453 50776
rect 4672 50736 4678 50748
rect 20441 50745 20453 50748
rect 20487 50745 20499 50779
rect 22465 50779 22523 50785
rect 22465 50776 22477 50779
rect 20441 50739 20499 50745
rect 22066 50748 22477 50776
rect 18414 50668 18420 50720
rect 18472 50708 18478 50720
rect 22066 50708 22094 50748
rect 22465 50745 22477 50748
rect 22511 50745 22523 50779
rect 22465 50739 22523 50745
rect 23014 50736 23020 50788
rect 23072 50776 23078 50788
rect 25317 50779 25375 50785
rect 25317 50776 25329 50779
rect 23072 50748 25329 50776
rect 23072 50736 23078 50748
rect 25317 50745 25329 50748
rect 25363 50745 25375 50779
rect 25317 50739 25375 50745
rect 26326 50736 26332 50788
rect 26384 50776 26390 50788
rect 26697 50779 26755 50785
rect 26697 50776 26709 50779
rect 26384 50748 26709 50776
rect 26384 50736 26390 50748
rect 26697 50745 26709 50748
rect 26743 50745 26755 50779
rect 26697 50739 26755 50745
rect 18472 50680 22094 50708
rect 26712 50708 26740 50739
rect 26786 50736 26792 50788
rect 26844 50776 26850 50788
rect 26844 50748 26889 50776
rect 26844 50736 26850 50748
rect 27982 50736 27988 50788
rect 28040 50776 28046 50788
rect 30561 50779 30619 50785
rect 30561 50776 30573 50779
rect 28040 50748 30573 50776
rect 28040 50736 28046 50748
rect 30561 50745 30573 50748
rect 30607 50745 30619 50779
rect 32766 50776 32772 50788
rect 32727 50748 32772 50776
rect 30561 50739 30619 50745
rect 32766 50736 32772 50748
rect 32824 50736 32830 50788
rect 36906 50736 36912 50788
rect 36964 50776 36970 50788
rect 37016 50776 37044 50807
rect 38102 50804 38108 50816
rect 38160 50804 38166 50856
rect 36964 50748 37044 50776
rect 37093 50779 37151 50785
rect 36964 50736 36970 50748
rect 37093 50745 37105 50779
rect 37139 50745 37151 50779
rect 37093 50739 37151 50745
rect 27522 50708 27528 50720
rect 26712 50680 27528 50708
rect 18472 50668 18478 50680
rect 27522 50668 27528 50680
rect 27580 50668 27586 50720
rect 27706 50668 27712 50720
rect 27764 50708 27770 50720
rect 28353 50711 28411 50717
rect 28353 50708 28365 50711
rect 27764 50680 28365 50708
rect 27764 50668 27770 50680
rect 28353 50677 28365 50680
rect 28399 50677 28411 50711
rect 28353 50671 28411 50677
rect 36998 50668 37004 50720
rect 37056 50708 37062 50720
rect 37108 50708 37136 50739
rect 37366 50708 37372 50720
rect 37056 50680 37136 50708
rect 37327 50680 37372 50708
rect 37056 50668 37062 50680
rect 37366 50668 37372 50680
rect 37424 50668 37430 50720
rect 1104 50618 38824 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 38824 50618
rect 1104 50544 38824 50566
rect 25314 50504 25320 50516
rect 25275 50476 25320 50504
rect 25314 50464 25320 50476
rect 25372 50464 25378 50516
rect 36906 50464 36912 50516
rect 36964 50464 36970 50516
rect 36998 50464 37004 50516
rect 37056 50504 37062 50516
rect 37056 50476 37136 50504
rect 37056 50464 37062 50476
rect 36924 50436 36952 50464
rect 36924 50408 37044 50436
rect 7282 50368 7288 50380
rect 7243 50340 7288 50368
rect 7282 50328 7288 50340
rect 7340 50328 7346 50380
rect 12250 50328 12256 50380
rect 12308 50368 12314 50380
rect 25225 50371 25283 50377
rect 25225 50368 25237 50371
rect 12308 50340 25237 50368
rect 12308 50328 12314 50340
rect 25225 50337 25237 50340
rect 25271 50337 25283 50371
rect 25225 50331 25283 50337
rect 35802 50328 35808 50380
rect 35860 50368 35866 50380
rect 36906 50377 36912 50380
rect 36081 50371 36139 50377
rect 36081 50368 36093 50371
rect 35860 50340 36093 50368
rect 35860 50328 35866 50340
rect 36081 50337 36093 50340
rect 36127 50337 36139 50371
rect 36081 50331 36139 50337
rect 36725 50371 36783 50377
rect 36725 50337 36737 50371
rect 36771 50337 36783 50371
rect 36725 50331 36783 50337
rect 36873 50371 36912 50377
rect 36873 50337 36885 50371
rect 36873 50331 36912 50337
rect 20990 50260 20996 50312
rect 21048 50300 21054 50312
rect 27982 50300 27988 50312
rect 21048 50272 27988 50300
rect 21048 50260 21054 50272
rect 27982 50260 27988 50272
rect 28040 50260 28046 50312
rect 29914 50260 29920 50312
rect 29972 50300 29978 50312
rect 29972 50272 36308 50300
rect 29972 50260 29978 50272
rect 21082 50192 21088 50244
rect 21140 50232 21146 50244
rect 21140 50204 22094 50232
rect 21140 50192 21146 50204
rect 7466 50164 7472 50176
rect 7427 50136 7472 50164
rect 7466 50124 7472 50136
rect 7524 50124 7530 50176
rect 22066 50164 22094 50204
rect 26510 50192 26516 50244
rect 26568 50232 26574 50244
rect 34514 50232 34520 50244
rect 26568 50204 34520 50232
rect 26568 50192 26574 50204
rect 34514 50192 34520 50204
rect 34572 50192 34578 50244
rect 36280 50241 36308 50272
rect 36265 50235 36323 50241
rect 36265 50201 36277 50235
rect 36311 50201 36323 50235
rect 36740 50232 36768 50331
rect 36906 50328 36912 50331
rect 36964 50328 36970 50380
rect 37016 50377 37044 50408
rect 37108 50377 37136 50476
rect 37001 50371 37059 50377
rect 37001 50337 37013 50371
rect 37047 50337 37059 50371
rect 37001 50331 37059 50337
rect 37093 50371 37151 50377
rect 37093 50337 37105 50371
rect 37139 50337 37151 50371
rect 37093 50331 37151 50337
rect 37231 50371 37289 50377
rect 37231 50337 37243 50371
rect 37277 50368 37289 50371
rect 38654 50368 38660 50380
rect 37277 50340 38660 50368
rect 37277 50337 37289 50340
rect 37231 50331 37289 50337
rect 37016 50300 37044 50331
rect 38654 50328 38660 50340
rect 38712 50328 38718 50380
rect 37550 50300 37556 50312
rect 37016 50272 37556 50300
rect 37550 50260 37556 50272
rect 37608 50260 37614 50312
rect 37458 50232 37464 50244
rect 36740 50204 37464 50232
rect 36265 50195 36323 50201
rect 37458 50192 37464 50204
rect 37516 50192 37522 50244
rect 29362 50164 29368 50176
rect 22066 50136 29368 50164
rect 29362 50124 29368 50136
rect 29420 50124 29426 50176
rect 32582 50124 32588 50176
rect 32640 50164 32646 50176
rect 37369 50167 37427 50173
rect 37369 50164 37381 50167
rect 32640 50136 37381 50164
rect 32640 50124 32646 50136
rect 37369 50133 37381 50136
rect 37415 50133 37427 50167
rect 37369 50127 37427 50133
rect 1104 50074 38824 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 38824 50074
rect 1104 50000 38824 50022
rect 27065 49963 27123 49969
rect 27065 49929 27077 49963
rect 27111 49960 27123 49963
rect 27890 49960 27896 49972
rect 27111 49932 27896 49960
rect 27111 49929 27123 49932
rect 27065 49923 27123 49929
rect 27890 49920 27896 49932
rect 27948 49920 27954 49972
rect 36081 49963 36139 49969
rect 36081 49929 36093 49963
rect 36127 49960 36139 49963
rect 36814 49960 36820 49972
rect 36127 49932 36820 49960
rect 36127 49929 36139 49932
rect 36081 49923 36139 49929
rect 36814 49920 36820 49932
rect 36872 49920 36878 49972
rect 37366 49960 37372 49972
rect 36924 49932 37372 49960
rect 2041 49895 2099 49901
rect 2041 49861 2053 49895
rect 2087 49892 2099 49895
rect 8386 49892 8392 49904
rect 2087 49864 8392 49892
rect 2087 49861 2099 49864
rect 2041 49855 2099 49861
rect 8386 49852 8392 49864
rect 8444 49852 8450 49904
rect 21358 49852 21364 49904
rect 21416 49892 21422 49904
rect 28534 49892 28540 49904
rect 21416 49864 28540 49892
rect 21416 49852 21422 49864
rect 28534 49852 28540 49864
rect 28592 49852 28598 49904
rect 34330 49892 34336 49904
rect 31726 49864 34336 49892
rect 31726 49824 31754 49864
rect 34330 49852 34336 49864
rect 34388 49852 34394 49904
rect 36924 49892 36952 49932
rect 37366 49920 37372 49932
rect 37424 49920 37430 49972
rect 37918 49960 37924 49972
rect 37879 49932 37924 49960
rect 37918 49920 37924 49932
rect 37976 49920 37982 49972
rect 37090 49892 37096 49904
rect 34440 49864 36952 49892
rect 37016 49864 37096 49892
rect 26528 49796 31754 49824
rect 1854 49756 1860 49768
rect 1815 49728 1860 49756
rect 1854 49716 1860 49728
rect 1912 49716 1918 49768
rect 23198 49716 23204 49768
rect 23256 49756 23262 49768
rect 26528 49765 26556 49796
rect 34054 49784 34060 49836
rect 34112 49824 34118 49836
rect 34440 49824 34468 49864
rect 37016 49824 37044 49864
rect 37090 49852 37096 49864
rect 37148 49852 37154 49904
rect 37366 49824 37372 49836
rect 34112 49796 34468 49824
rect 36740 49796 37044 49824
rect 37154 49796 37372 49824
rect 34112 49784 34118 49796
rect 26513 49759 26571 49765
rect 23256 49728 26464 49756
rect 23256 49716 23262 49728
rect 1670 49648 1676 49700
rect 1728 49688 1734 49700
rect 7650 49688 7656 49700
rect 1728 49660 7656 49688
rect 1728 49648 1734 49660
rect 7650 49648 7656 49660
rect 7708 49648 7714 49700
rect 7742 49648 7748 49700
rect 7800 49688 7806 49700
rect 8386 49688 8392 49700
rect 7800 49660 8392 49688
rect 7800 49648 7806 49660
rect 8386 49648 8392 49660
rect 8444 49648 8450 49700
rect 8938 49648 8944 49700
rect 8996 49688 9002 49700
rect 10134 49688 10140 49700
rect 8996 49660 10140 49688
rect 8996 49648 9002 49660
rect 10134 49648 10140 49660
rect 10192 49648 10198 49700
rect 26436 49688 26464 49728
rect 26513 49725 26525 49759
rect 26559 49725 26571 49759
rect 26886 49759 26944 49765
rect 26886 49756 26898 49759
rect 26513 49719 26571 49725
rect 26620 49728 26898 49756
rect 26620 49688 26648 49728
rect 26886 49725 26898 49728
rect 26932 49725 26944 49759
rect 27522 49756 27528 49768
rect 26886 49719 26944 49725
rect 26988 49728 27528 49756
rect 26436 49660 26648 49688
rect 26697 49691 26755 49697
rect 26697 49657 26709 49691
rect 26743 49657 26755 49691
rect 26697 49651 26755 49657
rect 26712 49620 26740 49651
rect 26786 49648 26792 49700
rect 26844 49688 26850 49700
rect 26844 49660 26889 49688
rect 26844 49648 26850 49660
rect 26988 49620 27016 49728
rect 27522 49716 27528 49728
rect 27580 49716 27586 49768
rect 36262 49756 36268 49768
rect 36223 49728 36268 49756
rect 36262 49716 36268 49728
rect 36320 49716 36326 49768
rect 36740 49765 36768 49796
rect 36725 49759 36783 49765
rect 36725 49725 36737 49759
rect 36771 49725 36783 49759
rect 36725 49719 36783 49725
rect 36814 49716 36820 49768
rect 36872 49756 36878 49768
rect 37001 49759 37059 49765
rect 36872 49728 36917 49756
rect 36872 49716 36878 49728
rect 37001 49725 37013 49759
rect 37047 49756 37059 49759
rect 37154 49756 37182 49796
rect 37366 49784 37372 49796
rect 37424 49784 37430 49836
rect 38562 49824 38568 49836
rect 37936 49796 38568 49824
rect 37047 49728 37182 49756
rect 37231 49759 37289 49765
rect 37047 49725 37059 49728
rect 37001 49719 37059 49725
rect 37231 49725 37243 49759
rect 37277 49756 37289 49759
rect 37936 49756 37964 49796
rect 38562 49784 38568 49796
rect 38620 49784 38626 49836
rect 38102 49756 38108 49768
rect 37277 49728 37964 49756
rect 38063 49728 38108 49756
rect 37277 49725 37289 49728
rect 37231 49719 37289 49725
rect 38102 49716 38108 49728
rect 38160 49716 38166 49768
rect 29362 49648 29368 49700
rect 29420 49688 29426 49700
rect 37090 49688 37096 49700
rect 29420 49660 36216 49688
rect 37051 49660 37096 49688
rect 29420 49648 29426 49660
rect 26712 49592 27016 49620
rect 34146 49580 34152 49632
rect 34204 49620 34210 49632
rect 35710 49620 35716 49632
rect 34204 49592 35716 49620
rect 34204 49580 34210 49592
rect 35710 49580 35716 49592
rect 35768 49580 35774 49632
rect 36188 49620 36216 49660
rect 37090 49648 37096 49660
rect 37148 49648 37154 49700
rect 37369 49623 37427 49629
rect 37369 49620 37381 49623
rect 36188 49592 37381 49620
rect 37369 49589 37381 49592
rect 37415 49589 37427 49623
rect 37369 49583 37427 49589
rect 1104 49530 38824 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 38824 49530
rect 1104 49456 38824 49478
rect 24486 49416 24492 49428
rect 23124 49388 24492 49416
rect 2041 49351 2099 49357
rect 2041 49317 2053 49351
rect 2087 49348 2099 49351
rect 8018 49348 8024 49360
rect 2087 49320 8024 49348
rect 2087 49317 2099 49320
rect 2041 49311 2099 49317
rect 8018 49308 8024 49320
rect 8076 49308 8082 49360
rect 1854 49280 1860 49292
rect 1815 49252 1860 49280
rect 1854 49240 1860 49252
rect 1912 49240 1918 49292
rect 23124 49289 23152 49388
rect 24486 49376 24492 49388
rect 24544 49376 24550 49428
rect 35526 49376 35532 49428
rect 35584 49416 35590 49428
rect 37550 49416 37556 49428
rect 35584 49388 37556 49416
rect 35584 49376 35590 49388
rect 37550 49376 37556 49388
rect 37608 49376 37614 49428
rect 27706 49348 27712 49360
rect 23400 49320 27712 49348
rect 23400 49289 23428 49320
rect 27706 49308 27712 49320
rect 27764 49308 27770 49360
rect 35710 49308 35716 49360
rect 35768 49348 35774 49360
rect 36909 49351 36967 49357
rect 35768 49320 36768 49348
rect 35768 49308 35774 49320
rect 23109 49283 23167 49289
rect 23109 49249 23121 49283
rect 23155 49249 23167 49283
rect 23109 49243 23167 49249
rect 23385 49283 23443 49289
rect 23385 49249 23397 49283
rect 23431 49249 23443 49283
rect 23385 49243 23443 49249
rect 23845 49283 23903 49289
rect 23845 49249 23857 49283
rect 23891 49280 23903 49283
rect 25866 49280 25872 49292
rect 23891 49252 25872 49280
rect 23891 49249 23903 49252
rect 23845 49243 23903 49249
rect 25866 49240 25872 49252
rect 25924 49240 25930 49292
rect 35618 49280 35624 49292
rect 35579 49252 35624 49280
rect 35618 49240 35624 49252
rect 35676 49240 35682 49292
rect 35802 49280 35808 49292
rect 35763 49252 35808 49280
rect 35802 49240 35808 49252
rect 35860 49240 35866 49292
rect 35897 49283 35955 49289
rect 35897 49249 35909 49283
rect 35943 49249 35955 49283
rect 35897 49243 35955 49249
rect 35989 49283 36047 49289
rect 35989 49249 36001 49283
rect 36035 49280 36047 49283
rect 36630 49280 36636 49292
rect 36035 49252 36492 49280
rect 36591 49252 36636 49280
rect 36035 49249 36047 49252
rect 35989 49243 36047 49249
rect 2038 49172 2044 49224
rect 2096 49212 2102 49224
rect 22186 49212 22192 49224
rect 2096 49184 22192 49212
rect 2096 49172 2102 49184
rect 22186 49172 22192 49184
rect 22244 49172 22250 49224
rect 23474 49172 23480 49224
rect 23532 49212 23538 49224
rect 23937 49215 23995 49221
rect 23937 49212 23949 49215
rect 23532 49184 23949 49212
rect 23532 49172 23538 49184
rect 23937 49181 23949 49184
rect 23983 49181 23995 49215
rect 35912 49212 35940 49243
rect 36354 49212 36360 49224
rect 35912 49184 36360 49212
rect 23937 49175 23995 49181
rect 36354 49172 36360 49184
rect 36412 49172 36418 49224
rect 8202 49104 8208 49156
rect 8260 49144 8266 49156
rect 24213 49147 24271 49153
rect 24213 49144 24225 49147
rect 8260 49116 24225 49144
rect 8260 49104 8266 49116
rect 24213 49113 24225 49116
rect 24259 49113 24271 49147
rect 24213 49107 24271 49113
rect 35618 49104 35624 49156
rect 35676 49144 35682 49156
rect 36464 49144 36492 49252
rect 36630 49240 36636 49252
rect 36688 49240 36694 49292
rect 36740 49289 36768 49320
rect 36909 49317 36921 49351
rect 36955 49348 36967 49351
rect 37366 49348 37372 49360
rect 36955 49320 37372 49348
rect 36955 49317 36967 49320
rect 36909 49311 36967 49317
rect 37366 49308 37372 49320
rect 37424 49308 37430 49360
rect 36726 49283 36784 49289
rect 36726 49249 36738 49283
rect 36772 49249 36784 49283
rect 36998 49280 37004 49292
rect 36959 49252 37004 49280
rect 36726 49243 36784 49249
rect 36998 49240 37004 49252
rect 37056 49240 37062 49292
rect 37139 49283 37197 49289
rect 37139 49249 37151 49283
rect 37185 49280 37197 49283
rect 39574 49280 39580 49292
rect 37185 49252 39580 49280
rect 37185 49249 37197 49252
rect 37139 49243 37197 49249
rect 39574 49240 39580 49252
rect 39632 49240 39638 49292
rect 35676 49116 36492 49144
rect 35676 49104 35682 49116
rect 36173 49079 36231 49085
rect 36173 49045 36185 49079
rect 36219 49076 36231 49079
rect 36538 49076 36544 49088
rect 36219 49048 36544 49076
rect 36219 49045 36231 49048
rect 36173 49039 36231 49045
rect 36538 49036 36544 49048
rect 36596 49036 36602 49088
rect 37274 49076 37280 49088
rect 37235 49048 37280 49076
rect 37274 49036 37280 49048
rect 37332 49036 37338 49088
rect 1104 48986 38824 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 38824 48986
rect 1104 48912 38824 48934
rect 28902 48832 28908 48884
rect 28960 48872 28966 48884
rect 29454 48872 29460 48884
rect 28960 48844 29460 48872
rect 28960 48832 28966 48844
rect 29454 48832 29460 48844
rect 29512 48832 29518 48884
rect 35989 48875 36047 48881
rect 35989 48841 36001 48875
rect 36035 48872 36047 48875
rect 36906 48872 36912 48884
rect 36035 48844 36912 48872
rect 36035 48841 36047 48844
rect 35989 48835 36047 48841
rect 36906 48832 36912 48844
rect 36964 48832 36970 48884
rect 37734 48832 37740 48884
rect 37792 48872 37798 48884
rect 38013 48875 38071 48881
rect 38013 48872 38025 48875
rect 37792 48844 38025 48872
rect 37792 48832 37798 48844
rect 38013 48841 38025 48844
rect 38059 48841 38071 48875
rect 38013 48835 38071 48841
rect 27706 48764 27712 48816
rect 27764 48804 27770 48816
rect 37274 48804 37280 48816
rect 27764 48776 37280 48804
rect 27764 48764 27770 48776
rect 37274 48764 37280 48776
rect 37332 48764 37338 48816
rect 20070 48696 20076 48748
rect 20128 48736 20134 48748
rect 21266 48736 21272 48748
rect 20128 48708 21272 48736
rect 20128 48696 20134 48708
rect 21266 48696 21272 48708
rect 21324 48696 21330 48748
rect 34606 48696 34612 48748
rect 34664 48736 34670 48748
rect 35158 48736 35164 48748
rect 34664 48708 35164 48736
rect 34664 48696 34670 48708
rect 35158 48696 35164 48708
rect 35216 48696 35222 48748
rect 37366 48736 37372 48748
rect 36924 48708 37372 48736
rect 7193 48671 7251 48677
rect 7193 48637 7205 48671
rect 7239 48668 7251 48671
rect 7282 48668 7288 48680
rect 7239 48640 7288 48668
rect 7239 48637 7251 48640
rect 7193 48631 7251 48637
rect 7282 48628 7288 48640
rect 7340 48628 7346 48680
rect 36173 48671 36231 48677
rect 36173 48637 36185 48671
rect 36219 48668 36231 48671
rect 36262 48668 36268 48680
rect 36219 48640 36268 48668
rect 36219 48637 36231 48640
rect 36173 48631 36231 48637
rect 36262 48628 36268 48640
rect 36320 48628 36326 48680
rect 36446 48628 36452 48680
rect 36504 48668 36510 48680
rect 36633 48671 36691 48677
rect 36633 48668 36645 48671
rect 36504 48640 36645 48668
rect 36504 48628 36510 48640
rect 36633 48637 36645 48640
rect 36679 48637 36691 48671
rect 36633 48631 36691 48637
rect 36726 48671 36784 48677
rect 36726 48637 36738 48671
rect 36772 48637 36784 48671
rect 36726 48631 36784 48637
rect 34606 48560 34612 48612
rect 34664 48600 34670 48612
rect 36740 48600 36768 48631
rect 36924 48612 36952 48708
rect 37366 48696 37372 48708
rect 37424 48696 37430 48748
rect 37139 48671 37197 48677
rect 37139 48637 37151 48671
rect 37185 48668 37197 48671
rect 38838 48668 38844 48680
rect 37185 48640 38844 48668
rect 37185 48637 37197 48640
rect 37139 48631 37197 48637
rect 38838 48628 38844 48640
rect 38896 48628 38902 48680
rect 36906 48600 36912 48612
rect 34664 48572 36768 48600
rect 36867 48572 36912 48600
rect 34664 48560 34670 48572
rect 36906 48560 36912 48572
rect 36964 48560 36970 48612
rect 36998 48560 37004 48612
rect 37056 48600 37062 48612
rect 37056 48572 37101 48600
rect 37056 48560 37062 48572
rect 37734 48560 37740 48612
rect 37792 48600 37798 48612
rect 37921 48603 37979 48609
rect 37921 48600 37933 48603
rect 37792 48572 37933 48600
rect 37792 48560 37798 48572
rect 37921 48569 37933 48572
rect 37967 48569 37979 48603
rect 37921 48563 37979 48569
rect 7374 48532 7380 48544
rect 7335 48504 7380 48532
rect 7374 48492 7380 48504
rect 7432 48492 7438 48544
rect 37090 48492 37096 48544
rect 37148 48532 37154 48544
rect 37277 48535 37335 48541
rect 37277 48532 37289 48535
rect 37148 48504 37289 48532
rect 37148 48492 37154 48504
rect 37277 48501 37289 48504
rect 37323 48501 37335 48535
rect 37277 48495 37335 48501
rect 1104 48442 38824 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 38824 48442
rect 1104 48368 38824 48390
rect 1854 48260 1860 48272
rect 1815 48232 1860 48260
rect 1854 48220 1860 48232
rect 1912 48220 1918 48272
rect 2038 48260 2044 48272
rect 1999 48232 2044 48260
rect 2038 48220 2044 48232
rect 2096 48220 2102 48272
rect 2314 48220 2320 48272
rect 2372 48260 2378 48272
rect 2372 48232 6914 48260
rect 2372 48220 2378 48232
rect 6886 48192 6914 48232
rect 19978 48220 19984 48272
rect 20036 48260 20042 48272
rect 25222 48260 25228 48272
rect 20036 48232 25228 48260
rect 20036 48220 20042 48232
rect 25222 48220 25228 48232
rect 25280 48220 25286 48272
rect 35802 48220 35808 48272
rect 35860 48260 35866 48272
rect 36262 48260 36268 48272
rect 35860 48232 36268 48260
rect 35860 48220 35866 48232
rect 36262 48220 36268 48232
rect 36320 48260 36326 48272
rect 37001 48263 37059 48269
rect 37001 48260 37013 48263
rect 36320 48232 37013 48260
rect 36320 48220 36326 48232
rect 37001 48229 37013 48232
rect 37047 48229 37059 48263
rect 37001 48223 37059 48229
rect 37093 48263 37151 48269
rect 37093 48229 37105 48263
rect 37139 48260 37151 48263
rect 37274 48260 37280 48272
rect 37139 48232 37280 48260
rect 37139 48229 37151 48232
rect 37093 48223 37151 48229
rect 37274 48220 37280 48232
rect 37332 48220 37338 48272
rect 8757 48195 8815 48201
rect 8757 48192 8769 48195
rect 6886 48164 8769 48192
rect 8757 48161 8769 48164
rect 8803 48161 8815 48195
rect 35526 48192 35532 48204
rect 35487 48164 35532 48192
rect 8757 48155 8815 48161
rect 35526 48152 35532 48164
rect 35584 48152 35590 48204
rect 36354 48192 36360 48204
rect 36315 48164 36360 48192
rect 36354 48152 36360 48164
rect 36412 48152 36418 48204
rect 36630 48152 36636 48204
rect 36688 48192 36694 48204
rect 36817 48195 36875 48201
rect 36817 48192 36829 48195
rect 36688 48164 36829 48192
rect 36688 48152 36694 48164
rect 36817 48161 36829 48164
rect 36863 48161 36875 48195
rect 36817 48155 36875 48161
rect 37185 48195 37243 48201
rect 37185 48161 37197 48195
rect 37231 48192 37243 48195
rect 38562 48192 38568 48204
rect 37231 48164 38568 48192
rect 37231 48161 37243 48164
rect 37185 48155 37243 48161
rect 38562 48152 38568 48164
rect 38620 48152 38626 48204
rect 7466 48084 7472 48136
rect 7524 48124 7530 48136
rect 8573 48127 8631 48133
rect 8573 48124 8585 48127
rect 7524 48096 8585 48124
rect 7524 48084 7530 48096
rect 8573 48093 8585 48096
rect 8619 48093 8631 48127
rect 8573 48087 8631 48093
rect 35158 48084 35164 48136
rect 35216 48124 35222 48136
rect 37918 48124 37924 48136
rect 35216 48096 37924 48124
rect 35216 48084 35222 48096
rect 37918 48084 37924 48096
rect 37976 48084 37982 48136
rect 22094 48016 22100 48068
rect 22152 48056 22158 48068
rect 28534 48056 28540 48068
rect 22152 48028 28540 48056
rect 22152 48016 22158 48028
rect 28534 48016 28540 48028
rect 28592 48016 28598 48068
rect 35434 48016 35440 48068
rect 35492 48056 35498 48068
rect 35713 48059 35771 48065
rect 35713 48056 35725 48059
rect 35492 48028 35725 48056
rect 35492 48016 35498 48028
rect 35713 48025 35725 48028
rect 35759 48025 35771 48059
rect 35713 48019 35771 48025
rect 36173 48059 36231 48065
rect 36173 48025 36185 48059
rect 36219 48056 36231 48059
rect 38194 48056 38200 48068
rect 36219 48028 38200 48056
rect 36219 48025 36231 48028
rect 36173 48019 36231 48025
rect 38194 48016 38200 48028
rect 38252 48016 38258 48068
rect 8941 47991 8999 47997
rect 8941 47957 8953 47991
rect 8987 47988 8999 47991
rect 14642 47988 14648 48000
rect 8987 47960 14648 47988
rect 8987 47957 8999 47960
rect 8941 47951 8999 47957
rect 14642 47948 14648 47960
rect 14700 47948 14706 48000
rect 22278 47948 22284 48000
rect 22336 47988 22342 48000
rect 27890 47988 27896 48000
rect 22336 47960 27896 47988
rect 22336 47948 22342 47960
rect 27890 47948 27896 47960
rect 27948 47948 27954 48000
rect 37366 47988 37372 48000
rect 37327 47960 37372 47988
rect 37366 47948 37372 47960
rect 37424 47948 37430 48000
rect 1104 47898 38824 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 38824 47898
rect 1104 47824 38824 47846
rect 26881 47787 26939 47793
rect 26881 47753 26893 47787
rect 26927 47784 26939 47787
rect 27338 47784 27344 47796
rect 26927 47756 27344 47784
rect 26927 47753 26939 47756
rect 26881 47747 26939 47753
rect 27338 47744 27344 47756
rect 27396 47744 27402 47796
rect 35894 47744 35900 47796
rect 35952 47784 35958 47796
rect 36081 47787 36139 47793
rect 36081 47784 36093 47787
rect 35952 47756 36093 47784
rect 35952 47744 35958 47756
rect 36081 47753 36093 47756
rect 36127 47753 36139 47787
rect 36081 47747 36139 47753
rect 2038 47676 2044 47728
rect 2096 47716 2102 47728
rect 23198 47716 23204 47728
rect 2096 47688 23204 47716
rect 2096 47676 2102 47688
rect 23198 47676 23204 47688
rect 23256 47676 23262 47728
rect 26234 47676 26240 47728
rect 26292 47716 26298 47728
rect 26292 47688 27384 47716
rect 26292 47676 26298 47688
rect 27356 47660 27384 47688
rect 36354 47676 36360 47728
rect 36412 47716 36418 47728
rect 36630 47716 36636 47728
rect 36412 47688 36636 47716
rect 36412 47676 36418 47688
rect 36630 47676 36636 47688
rect 36688 47716 36694 47728
rect 37182 47716 37188 47728
rect 36688 47688 37188 47716
rect 36688 47676 36694 47688
rect 37182 47676 37188 47688
rect 37240 47716 37246 47728
rect 37240 47688 37872 47716
rect 37240 47676 37246 47688
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 7466 47608 7472 47660
rect 7524 47648 7530 47660
rect 8205 47651 8263 47657
rect 8205 47648 8217 47651
rect 7524 47620 8217 47648
rect 7524 47608 7530 47620
rect 8205 47617 8217 47620
rect 8251 47648 8263 47651
rect 9493 47651 9551 47657
rect 9493 47648 9505 47651
rect 8251 47620 9505 47648
rect 8251 47617 8263 47620
rect 8205 47611 8263 47617
rect 9493 47617 9505 47620
rect 9539 47617 9551 47651
rect 9493 47611 9551 47617
rect 26602 47608 26608 47660
rect 26660 47648 26666 47660
rect 27062 47648 27068 47660
rect 26660 47620 27068 47648
rect 26660 47608 26666 47620
rect 27062 47608 27068 47620
rect 27120 47608 27126 47660
rect 27338 47608 27344 47660
rect 27396 47608 27402 47660
rect 27890 47608 27896 47660
rect 27948 47648 27954 47660
rect 27948 47620 37596 47648
rect 27948 47608 27954 47620
rect 1394 47580 1400 47592
rect 1355 47552 1400 47580
rect 1394 47540 1400 47552
rect 1452 47540 1458 47592
rect 7006 47540 7012 47592
rect 7064 47580 7070 47592
rect 7101 47583 7159 47589
rect 7101 47580 7113 47583
rect 7064 47552 7113 47580
rect 7064 47540 7070 47552
rect 7101 47549 7113 47552
rect 7147 47580 7159 47583
rect 7282 47580 7288 47592
rect 7147 47552 7288 47580
rect 7147 47549 7159 47552
rect 7101 47543 7159 47549
rect 7282 47540 7288 47552
rect 7340 47540 7346 47592
rect 8386 47580 8392 47592
rect 8347 47552 8392 47580
rect 8386 47540 8392 47552
rect 8444 47540 8450 47592
rect 9677 47583 9735 47589
rect 9677 47549 9689 47583
rect 9723 47580 9735 47583
rect 9766 47580 9772 47592
rect 9723 47552 9772 47580
rect 9723 47549 9735 47552
rect 9677 47543 9735 47549
rect 9766 47540 9772 47552
rect 9824 47540 9830 47592
rect 26329 47583 26387 47589
rect 26329 47580 26341 47583
rect 26160 47552 26341 47580
rect 2590 47472 2596 47524
rect 2648 47512 2654 47524
rect 8202 47512 8208 47524
rect 2648 47484 8208 47512
rect 2648 47472 2654 47484
rect 8202 47472 8208 47484
rect 8260 47472 8266 47524
rect 8573 47515 8631 47521
rect 8573 47481 8585 47515
rect 8619 47512 8631 47515
rect 13262 47512 13268 47524
rect 8619 47484 13268 47512
rect 8619 47481 8631 47484
rect 8573 47475 8631 47481
rect 13262 47472 13268 47484
rect 13320 47472 13326 47524
rect 7282 47444 7288 47456
rect 7243 47416 7288 47444
rect 7282 47404 7288 47416
rect 7340 47404 7346 47456
rect 9861 47447 9919 47453
rect 9861 47413 9873 47447
rect 9907 47444 9919 47447
rect 10226 47444 10232 47456
rect 9907 47416 10232 47444
rect 9907 47413 9919 47416
rect 9861 47407 9919 47413
rect 10226 47404 10232 47416
rect 10284 47404 10290 47456
rect 26160 47444 26188 47552
rect 26329 47549 26341 47552
rect 26375 47549 26387 47583
rect 26329 47543 26387 47549
rect 26418 47540 26424 47592
rect 26476 47580 26482 47592
rect 26702 47583 26760 47589
rect 26702 47580 26714 47583
rect 26476 47552 26714 47580
rect 26476 47540 26482 47552
rect 26702 47549 26714 47552
rect 26748 47549 26760 47583
rect 26702 47543 26760 47549
rect 35802 47540 35808 47592
rect 35860 47580 35866 47592
rect 35897 47583 35955 47589
rect 35897 47580 35909 47583
rect 35860 47552 35909 47580
rect 35860 47540 35866 47552
rect 35897 47549 35909 47552
rect 35943 47549 35955 47583
rect 35897 47543 35955 47549
rect 35986 47540 35992 47592
rect 36044 47580 36050 47592
rect 36541 47583 36599 47589
rect 36541 47580 36553 47583
rect 36044 47552 36553 47580
rect 36044 47540 36050 47552
rect 36541 47549 36553 47552
rect 36587 47549 36599 47583
rect 36541 47543 36599 47549
rect 36630 47540 36636 47592
rect 36688 47580 36694 47592
rect 36817 47583 36875 47589
rect 36817 47580 36829 47583
rect 36688 47552 36829 47580
rect 36688 47540 36694 47552
rect 36817 47549 36829 47552
rect 36863 47549 36875 47583
rect 36817 47543 36875 47549
rect 36909 47583 36967 47589
rect 36909 47549 36921 47583
rect 36955 47580 36967 47583
rect 37274 47580 37280 47592
rect 36955 47552 37280 47580
rect 36955 47549 36967 47552
rect 36909 47543 36967 47549
rect 37274 47540 37280 47552
rect 37332 47540 37338 47592
rect 37568 47589 37596 47620
rect 37844 47589 37872 47688
rect 37553 47583 37611 47589
rect 37553 47549 37565 47583
rect 37599 47549 37611 47583
rect 37553 47543 37611 47549
rect 37829 47583 37887 47589
rect 37829 47549 37841 47583
rect 37875 47549 37887 47583
rect 37829 47543 37887 47549
rect 37921 47583 37979 47589
rect 37921 47549 37933 47583
rect 37967 47549 37979 47583
rect 37921 47543 37979 47549
rect 26510 47512 26516 47524
rect 26471 47484 26516 47512
rect 26510 47472 26516 47484
rect 26568 47472 26574 47524
rect 26602 47472 26608 47524
rect 26660 47512 26666 47524
rect 26660 47484 26705 47512
rect 26660 47472 26666 47484
rect 36262 47472 36268 47524
rect 36320 47512 36326 47524
rect 36725 47515 36783 47521
rect 36725 47512 36737 47515
rect 36320 47484 36737 47512
rect 36320 47472 36326 47484
rect 36725 47481 36737 47484
rect 36771 47512 36783 47515
rect 37182 47512 37188 47524
rect 36771 47484 37188 47512
rect 36771 47481 36783 47484
rect 36725 47475 36783 47481
rect 37182 47472 37188 47484
rect 37240 47512 37246 47524
rect 37737 47515 37795 47521
rect 37737 47512 37749 47515
rect 37240 47484 37749 47512
rect 37240 47472 37246 47484
rect 37737 47481 37749 47484
rect 37783 47481 37795 47515
rect 37737 47475 37795 47481
rect 27890 47444 27896 47456
rect 26160 47416 27896 47444
rect 27890 47404 27896 47416
rect 27948 47404 27954 47456
rect 35986 47404 35992 47456
rect 36044 47444 36050 47456
rect 36354 47444 36360 47456
rect 36044 47416 36360 47444
rect 36044 47404 36050 47416
rect 36354 47404 36360 47416
rect 36412 47404 36418 47456
rect 36446 47404 36452 47456
rect 36504 47444 36510 47456
rect 37093 47447 37151 47453
rect 37093 47444 37105 47447
rect 36504 47416 37105 47444
rect 36504 47404 36510 47416
rect 37093 47413 37105 47416
rect 37139 47413 37151 47447
rect 37093 47407 37151 47413
rect 37458 47404 37464 47456
rect 37516 47444 37522 47456
rect 37936 47444 37964 47543
rect 38102 47444 38108 47456
rect 37516 47416 37964 47444
rect 38063 47416 38108 47444
rect 37516 47404 37522 47416
rect 38102 47404 38108 47416
rect 38160 47404 38166 47456
rect 1104 47354 38824 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 38824 47354
rect 1104 47280 38824 47302
rect 4798 47200 4804 47252
rect 4856 47240 4862 47252
rect 8386 47240 8392 47252
rect 4856 47212 8392 47240
rect 4856 47200 4862 47212
rect 8386 47200 8392 47212
rect 8444 47200 8450 47252
rect 26418 47240 26424 47252
rect 12406 47212 26424 47240
rect 12406 47172 12434 47212
rect 26418 47200 26424 47212
rect 26476 47200 26482 47252
rect 26602 47200 26608 47252
rect 26660 47200 26666 47252
rect 33318 47200 33324 47252
rect 33376 47240 33382 47252
rect 35437 47243 35495 47249
rect 35437 47240 35449 47243
rect 33376 47212 35449 47240
rect 33376 47200 33382 47212
rect 35437 47209 35449 47212
rect 35483 47209 35495 47243
rect 35437 47203 35495 47209
rect 35897 47243 35955 47249
rect 35897 47209 35909 47243
rect 35943 47240 35955 47243
rect 36814 47240 36820 47252
rect 35943 47212 36820 47240
rect 35943 47209 35955 47212
rect 35897 47203 35955 47209
rect 36814 47200 36820 47212
rect 36872 47200 36878 47252
rect 6886 47144 12434 47172
rect 26513 47175 26571 47181
rect 2314 46860 2320 46912
rect 2372 46900 2378 46912
rect 6886 46900 6914 47144
rect 26513 47141 26525 47175
rect 26559 47172 26571 47175
rect 26620 47172 26648 47200
rect 34054 47172 34060 47184
rect 26559 47144 26648 47172
rect 33336 47144 34060 47172
rect 26559 47141 26571 47144
rect 26513 47135 26571 47141
rect 33336 47116 33364 47144
rect 34054 47132 34060 47144
rect 34112 47132 34118 47184
rect 7558 47104 7564 47116
rect 7519 47076 7564 47104
rect 7558 47064 7564 47076
rect 7616 47064 7622 47116
rect 8294 47064 8300 47116
rect 8352 47104 8358 47116
rect 8389 47107 8447 47113
rect 8389 47104 8401 47107
rect 8352 47076 8401 47104
rect 8352 47064 8358 47076
rect 8389 47073 8401 47076
rect 8435 47073 8447 47107
rect 9214 47104 9220 47116
rect 9175 47076 9220 47104
rect 8389 47067 8447 47073
rect 9214 47064 9220 47076
rect 9272 47064 9278 47116
rect 10042 47104 10048 47116
rect 10003 47076 10048 47104
rect 10042 47064 10048 47076
rect 10100 47064 10106 47116
rect 26234 47104 26240 47116
rect 26195 47076 26240 47104
rect 26234 47064 26240 47076
rect 26292 47064 26298 47116
rect 26418 47104 26424 47116
rect 26379 47076 26424 47104
rect 26418 47064 26424 47076
rect 26476 47064 26482 47116
rect 26610 47107 26668 47113
rect 26610 47073 26622 47107
rect 26656 47073 26668 47107
rect 26610 47067 26668 47073
rect 7377 47039 7435 47045
rect 7377 47005 7389 47039
rect 7423 47036 7435 47039
rect 7466 47036 7472 47048
rect 7423 47008 7472 47036
rect 7423 47005 7435 47008
rect 7377 46999 7435 47005
rect 7466 46996 7472 47008
rect 7524 47036 7530 47048
rect 8205 47039 8263 47045
rect 8205 47036 8217 47039
rect 7524 47008 8217 47036
rect 7524 46996 7530 47008
rect 8205 47005 8217 47008
rect 8251 47005 8263 47039
rect 9030 47036 9036 47048
rect 8991 47008 9036 47036
rect 8205 46999 8263 47005
rect 9030 46996 9036 47008
rect 9088 47036 9094 47048
rect 9861 47039 9919 47045
rect 9861 47036 9873 47039
rect 9088 47008 9873 47036
rect 9088 46996 9094 47008
rect 9861 47005 9873 47008
rect 9907 47005 9919 47039
rect 9861 46999 9919 47005
rect 15102 46996 15108 47048
rect 15160 47036 15166 47048
rect 26625 47036 26653 47067
rect 33318 47064 33324 47116
rect 33376 47064 33382 47116
rect 35250 47104 35256 47116
rect 35211 47076 35256 47104
rect 35250 47064 35256 47076
rect 35308 47064 35314 47116
rect 35802 47064 35808 47116
rect 35860 47104 35866 47116
rect 36081 47107 36139 47113
rect 36081 47104 36093 47107
rect 35860 47076 36093 47104
rect 35860 47064 35866 47076
rect 36081 47073 36093 47076
rect 36127 47073 36139 47107
rect 36081 47067 36139 47073
rect 36541 47107 36599 47113
rect 36541 47073 36553 47107
rect 36587 47104 36599 47107
rect 36630 47104 36636 47116
rect 36587 47076 36636 47104
rect 36587 47073 36599 47076
rect 36541 47067 36599 47073
rect 36630 47064 36636 47076
rect 36688 47064 36694 47116
rect 34054 47036 34060 47048
rect 15160 47008 26653 47036
rect 26712 47008 34060 47036
rect 15160 46996 15166 47008
rect 7745 46971 7803 46977
rect 7745 46937 7757 46971
rect 7791 46968 7803 46971
rect 7834 46968 7840 46980
rect 7791 46940 7840 46968
rect 7791 46937 7803 46940
rect 7745 46931 7803 46937
rect 7834 46928 7840 46940
rect 7892 46928 7898 46980
rect 8573 46971 8631 46977
rect 8573 46937 8585 46971
rect 8619 46968 8631 46971
rect 9214 46968 9220 46980
rect 8619 46940 9220 46968
rect 8619 46937 8631 46940
rect 8573 46931 8631 46937
rect 9214 46928 9220 46940
rect 9272 46928 9278 46980
rect 10229 46971 10287 46977
rect 10229 46937 10241 46971
rect 10275 46968 10287 46971
rect 17218 46968 17224 46980
rect 10275 46940 17224 46968
rect 10275 46937 10287 46940
rect 10229 46931 10287 46937
rect 17218 46928 17224 46940
rect 17276 46928 17282 46980
rect 26234 46928 26240 46980
rect 26292 46968 26298 46980
rect 26712 46968 26740 47008
rect 34054 46996 34060 47008
rect 34112 46996 34118 47048
rect 35434 46996 35440 47048
rect 35492 47036 35498 47048
rect 37274 47036 37280 47048
rect 35492 47008 37280 47036
rect 35492 46996 35498 47008
rect 37274 46996 37280 47008
rect 37332 46996 37338 47048
rect 26292 46940 26740 46968
rect 26789 46971 26847 46977
rect 26292 46928 26298 46940
rect 26789 46937 26801 46971
rect 26835 46968 26847 46971
rect 28074 46968 28080 46980
rect 26835 46940 28080 46968
rect 26835 46937 26847 46940
rect 26789 46931 26847 46937
rect 28074 46928 28080 46940
rect 28132 46928 28138 46980
rect 36725 46971 36783 46977
rect 36725 46937 36737 46971
rect 36771 46968 36783 46971
rect 39206 46968 39212 46980
rect 36771 46940 39212 46968
rect 36771 46937 36783 46940
rect 36725 46931 36783 46937
rect 39206 46928 39212 46940
rect 39264 46928 39270 46980
rect 9398 46900 9404 46912
rect 2372 46872 6914 46900
rect 9359 46872 9404 46900
rect 2372 46860 2378 46872
rect 9398 46860 9404 46872
rect 9456 46860 9462 46912
rect 22462 46860 22468 46912
rect 22520 46900 22526 46912
rect 27982 46900 27988 46912
rect 22520 46872 27988 46900
rect 22520 46860 22526 46872
rect 27982 46860 27988 46872
rect 28040 46860 28046 46912
rect 28626 46860 28632 46912
rect 28684 46900 28690 46912
rect 30282 46900 30288 46912
rect 28684 46872 30288 46900
rect 28684 46860 28690 46872
rect 30282 46860 30288 46872
rect 30340 46860 30346 46912
rect 36906 46860 36912 46912
rect 36964 46900 36970 46912
rect 38010 46900 38016 46912
rect 36964 46872 38016 46900
rect 36964 46860 36970 46872
rect 38010 46860 38016 46872
rect 38068 46860 38074 46912
rect 1104 46810 38824 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 38824 46810
rect 1104 46736 38824 46758
rect 26881 46699 26939 46705
rect 26881 46665 26893 46699
rect 26927 46696 26939 46699
rect 28902 46696 28908 46708
rect 26927 46668 28908 46696
rect 26927 46665 26939 46668
rect 26881 46659 26939 46665
rect 28902 46656 28908 46668
rect 28960 46656 28966 46708
rect 35986 46656 35992 46708
rect 36044 46696 36050 46708
rect 36044 46668 38056 46696
rect 36044 46656 36050 46668
rect 15102 46628 15108 46640
rect 6886 46600 15108 46628
rect 1394 46560 1400 46572
rect 1355 46532 1400 46560
rect 1394 46520 1400 46532
rect 1452 46520 1458 46572
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46560 1731 46563
rect 4062 46560 4068 46572
rect 1719 46532 4068 46560
rect 1719 46529 1731 46532
rect 1673 46523 1731 46529
rect 4062 46520 4068 46532
rect 4120 46520 4126 46572
rect 2130 46452 2136 46504
rect 2188 46492 2194 46504
rect 6886 46492 6914 46600
rect 15102 46588 15108 46600
rect 15160 46588 15166 46640
rect 30374 46628 30380 46640
rect 26436 46600 30380 46628
rect 9398 46520 9404 46572
rect 9456 46560 9462 46572
rect 17402 46560 17408 46572
rect 9456 46532 17408 46560
rect 9456 46520 9462 46532
rect 17402 46520 17408 46532
rect 17460 46520 17466 46572
rect 26436 46560 26464 46600
rect 30374 46588 30380 46600
rect 30432 46588 30438 46640
rect 36173 46631 36231 46637
rect 36173 46597 36185 46631
rect 36219 46628 36231 46631
rect 36906 46628 36912 46640
rect 36219 46600 36912 46628
rect 36219 46597 36231 46600
rect 36173 46591 36231 46597
rect 36906 46588 36912 46600
rect 36964 46588 36970 46640
rect 37093 46631 37151 46637
rect 37093 46597 37105 46631
rect 37139 46628 37151 46631
rect 37826 46628 37832 46640
rect 37139 46600 37832 46628
rect 37139 46597 37151 46600
rect 37093 46591 37151 46597
rect 37826 46588 37832 46600
rect 37884 46588 37890 46640
rect 26344 46532 26464 46560
rect 7006 46492 7012 46504
rect 2188 46464 6914 46492
rect 6967 46464 7012 46492
rect 2188 46452 2194 46464
rect 7006 46452 7012 46464
rect 7064 46452 7070 46504
rect 7742 46452 7748 46504
rect 7800 46492 7806 46504
rect 8205 46495 8263 46501
rect 8205 46492 8217 46495
rect 7800 46464 8217 46492
rect 7800 46452 7806 46464
rect 8205 46461 8217 46464
rect 8251 46461 8263 46495
rect 8386 46492 8392 46504
rect 8347 46464 8392 46492
rect 8205 46455 8263 46461
rect 8220 46424 8248 46455
rect 8386 46452 8392 46464
rect 8444 46452 8450 46504
rect 9493 46495 9551 46501
rect 9493 46461 9505 46495
rect 9539 46461 9551 46495
rect 9674 46492 9680 46504
rect 9635 46464 9680 46492
rect 9493 46455 9551 46461
rect 9030 46424 9036 46436
rect 8220 46396 9036 46424
rect 9030 46384 9036 46396
rect 9088 46424 9094 46436
rect 9508 46424 9536 46455
rect 9674 46452 9680 46464
rect 9732 46452 9738 46504
rect 26344 46501 26372 46532
rect 28902 46520 28908 46572
rect 28960 46560 28966 46572
rect 29362 46560 29368 46572
rect 28960 46532 29368 46560
rect 28960 46520 28966 46532
rect 29362 46520 29368 46532
rect 29420 46520 29426 46572
rect 31726 46532 37596 46560
rect 26329 46495 26387 46501
rect 26329 46461 26341 46495
rect 26375 46461 26387 46495
rect 26329 46455 26387 46461
rect 26418 46452 26424 46504
rect 26476 46492 26482 46504
rect 26702 46495 26760 46501
rect 26702 46492 26714 46495
rect 26476 46464 26714 46492
rect 26476 46452 26482 46464
rect 26702 46461 26714 46464
rect 26748 46461 26760 46495
rect 26702 46455 26760 46461
rect 27982 46452 27988 46504
rect 28040 46492 28046 46504
rect 31726 46492 31754 46532
rect 36354 46492 36360 46504
rect 28040 46464 31754 46492
rect 36315 46464 36360 46492
rect 28040 46452 28046 46464
rect 36354 46452 36360 46464
rect 36412 46452 36418 46504
rect 37568 46501 37596 46532
rect 37553 46495 37611 46501
rect 37553 46461 37565 46495
rect 37599 46461 37611 46495
rect 37918 46492 37924 46504
rect 37879 46464 37924 46492
rect 37553 46455 37611 46461
rect 37918 46452 37924 46464
rect 37976 46452 37982 46504
rect 26510 46424 26516 46436
rect 9088 46396 9536 46424
rect 26471 46396 26516 46424
rect 9088 46384 9094 46396
rect 26510 46384 26516 46396
rect 26568 46384 26574 46436
rect 26602 46384 26608 46436
rect 26660 46424 26666 46436
rect 26660 46396 26753 46424
rect 26660 46384 26666 46396
rect 35158 46384 35164 46436
rect 35216 46424 35222 46436
rect 36909 46427 36967 46433
rect 36909 46424 36921 46427
rect 35216 46396 36921 46424
rect 35216 46384 35222 46396
rect 36909 46393 36921 46396
rect 36955 46393 36967 46427
rect 36909 46387 36967 46393
rect 37182 46384 37188 46436
rect 37240 46424 37246 46436
rect 37737 46427 37795 46433
rect 37737 46424 37749 46427
rect 37240 46396 37749 46424
rect 37240 46384 37246 46396
rect 37737 46393 37749 46396
rect 37783 46393 37795 46427
rect 37737 46387 37795 46393
rect 37829 46427 37887 46433
rect 37829 46393 37841 46427
rect 37875 46424 37887 46427
rect 38028 46424 38056 46668
rect 37875 46396 38056 46424
rect 37875 46393 37887 46396
rect 37829 46387 37887 46393
rect 7190 46356 7196 46368
rect 7151 46328 7196 46356
rect 7190 46316 7196 46328
rect 7248 46316 7254 46368
rect 8570 46356 8576 46368
rect 8531 46328 8576 46356
rect 8570 46316 8576 46328
rect 8628 46316 8634 46368
rect 9858 46356 9864 46368
rect 9819 46328 9864 46356
rect 9858 46316 9864 46328
rect 9916 46316 9922 46368
rect 26234 46316 26240 46368
rect 26292 46356 26298 46368
rect 26620 46356 26648 46384
rect 26292 46328 26648 46356
rect 26292 46316 26298 46328
rect 30742 46316 30748 46368
rect 30800 46356 30806 46368
rect 31202 46356 31208 46368
rect 30800 46328 31208 46356
rect 30800 46316 30806 46328
rect 31202 46316 31208 46328
rect 31260 46316 31266 46368
rect 37274 46316 37280 46368
rect 37332 46356 37338 46368
rect 38105 46359 38163 46365
rect 38105 46356 38117 46359
rect 37332 46328 38117 46356
rect 37332 46316 37338 46328
rect 38105 46325 38117 46328
rect 38151 46325 38163 46359
rect 38105 46319 38163 46325
rect 1104 46266 38824 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 38824 46266
rect 1104 46192 38824 46214
rect 2774 46112 2780 46164
rect 2832 46152 2838 46164
rect 26418 46152 26424 46164
rect 2832 46124 26424 46152
rect 2832 46112 2838 46124
rect 26418 46112 26424 46124
rect 26476 46112 26482 46164
rect 32858 46152 32864 46164
rect 26528 46124 32864 46152
rect 2038 46084 2044 46096
rect 1999 46056 2044 46084
rect 2038 46044 2044 46056
rect 2096 46044 2102 46096
rect 6270 46044 6276 46096
rect 6328 46084 6334 46096
rect 26528 46084 26556 46124
rect 32858 46112 32864 46124
rect 32916 46112 32922 46164
rect 35253 46155 35311 46161
rect 35253 46121 35265 46155
rect 35299 46152 35311 46155
rect 35710 46152 35716 46164
rect 35299 46124 35716 46152
rect 35299 46121 35311 46124
rect 35253 46115 35311 46121
rect 35710 46112 35716 46124
rect 35768 46112 35774 46164
rect 35897 46155 35955 46161
rect 35897 46121 35909 46155
rect 35943 46152 35955 46155
rect 36722 46152 36728 46164
rect 35943 46124 36728 46152
rect 35943 46121 35955 46124
rect 35897 46115 35955 46121
rect 36722 46112 36728 46124
rect 36780 46112 36786 46164
rect 37185 46155 37243 46161
rect 37185 46121 37197 46155
rect 37231 46121 37243 46155
rect 37185 46115 37243 46121
rect 6328 46056 6914 46084
rect 6328 46044 6334 46056
rect 1854 46016 1860 46028
rect 1815 45988 1860 46016
rect 1854 45976 1860 45988
rect 1912 45976 1918 46028
rect 6886 46016 6914 46056
rect 26252 46056 26556 46084
rect 9125 46019 9183 46025
rect 9125 46016 9137 46019
rect 6886 45988 9137 46016
rect 9125 45985 9137 45988
rect 9171 45985 9183 46019
rect 9125 45979 9183 45985
rect 16298 45976 16304 46028
rect 16356 46016 16362 46028
rect 21358 46016 21364 46028
rect 16356 45988 21364 46016
rect 16356 45976 16362 45988
rect 21358 45976 21364 45988
rect 21416 45976 21422 46028
rect 26252 46025 26280 46056
rect 29914 46044 29920 46096
rect 29972 46084 29978 46096
rect 37200 46084 37228 46115
rect 38286 46112 38292 46164
rect 38344 46152 38350 46164
rect 38654 46152 38660 46164
rect 38344 46124 38660 46152
rect 38344 46112 38350 46124
rect 38654 46112 38660 46124
rect 38712 46112 38718 46164
rect 29972 46056 37228 46084
rect 29972 46044 29978 46056
rect 26237 46019 26295 46025
rect 26237 45985 26249 46019
rect 26283 45985 26295 46019
rect 26418 46016 26424 46028
rect 26379 45988 26424 46016
rect 26237 45979 26295 45985
rect 26418 45976 26424 45988
rect 26476 45976 26482 46028
rect 26513 46019 26571 46025
rect 26513 45985 26525 46019
rect 26559 45985 26571 46019
rect 26513 45979 26571 45985
rect 26610 46019 26668 46025
rect 26610 45985 26622 46019
rect 26656 45985 26668 46019
rect 26610 45979 26668 45985
rect 35437 46019 35495 46025
rect 35437 45985 35449 46019
rect 35483 46016 35495 46019
rect 35710 46016 35716 46028
rect 35483 45988 35716 46016
rect 35483 45985 35495 45988
rect 35437 45979 35495 45985
rect 7742 45908 7748 45960
rect 7800 45948 7806 45960
rect 8941 45951 8999 45957
rect 8941 45948 8953 45951
rect 7800 45920 8953 45948
rect 7800 45908 7806 45920
rect 8941 45917 8953 45920
rect 8987 45917 8999 45951
rect 26528 45948 26556 45979
rect 8941 45911 8999 45917
rect 26252 45920 26556 45948
rect 26252 45892 26280 45920
rect 26234 45840 26240 45892
rect 26292 45840 26298 45892
rect 9306 45812 9312 45824
rect 9267 45784 9312 45812
rect 9306 45772 9312 45784
rect 9364 45772 9370 45824
rect 20714 45772 20720 45824
rect 20772 45812 20778 45824
rect 26625 45812 26653 45979
rect 35710 45976 35716 45988
rect 35768 45976 35774 46028
rect 35802 45976 35808 46028
rect 35860 46016 35866 46028
rect 36081 46019 36139 46025
rect 36081 46016 36093 46019
rect 35860 45988 36093 46016
rect 35860 45976 35866 45988
rect 36081 45985 36093 45988
rect 36127 45985 36139 46019
rect 36538 46016 36544 46028
rect 36499 45988 36544 46016
rect 36081 45979 36139 45985
rect 36538 45976 36544 45988
rect 36596 45976 36602 46028
rect 36722 46025 36728 46028
rect 36689 46019 36728 46025
rect 36689 45985 36701 46019
rect 36689 45979 36728 45985
rect 36722 45976 36728 45979
rect 36780 45976 36786 46028
rect 36817 46019 36875 46025
rect 36817 45985 36829 46019
rect 36863 45985 36875 46019
rect 36817 45979 36875 45985
rect 36832 45948 36860 45979
rect 36906 45976 36912 46028
rect 36964 46016 36970 46028
rect 37045 46019 37103 46025
rect 36964 45988 37009 46016
rect 36964 45976 36970 45988
rect 37045 45985 37057 46019
rect 37091 45985 37103 46019
rect 37045 45979 37103 45985
rect 36556 45920 36860 45948
rect 36556 45892 36584 45920
rect 26789 45883 26847 45889
rect 26789 45849 26801 45883
rect 26835 45880 26847 45883
rect 27338 45880 27344 45892
rect 26835 45852 27344 45880
rect 26835 45849 26847 45852
rect 26789 45843 26847 45849
rect 27338 45840 27344 45852
rect 27396 45840 27402 45892
rect 31110 45840 31116 45892
rect 31168 45880 31174 45892
rect 32674 45880 32680 45892
rect 31168 45852 32680 45880
rect 31168 45840 31174 45852
rect 32674 45840 32680 45852
rect 32732 45840 32738 45892
rect 36078 45840 36084 45892
rect 36136 45880 36142 45892
rect 36354 45880 36360 45892
rect 36136 45852 36360 45880
rect 36136 45840 36142 45852
rect 36354 45840 36360 45852
rect 36412 45840 36418 45892
rect 36538 45840 36544 45892
rect 36596 45840 36602 45892
rect 20772 45784 26653 45812
rect 20772 45772 20778 45784
rect 33962 45772 33968 45824
rect 34020 45812 34026 45824
rect 37062 45812 37090 45979
rect 34020 45784 37090 45812
rect 34020 45772 34026 45784
rect 1104 45722 38824 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 38824 45722
rect 1104 45648 38824 45670
rect 7742 45608 7748 45620
rect 7703 45580 7748 45608
rect 7742 45568 7748 45580
rect 7800 45568 7806 45620
rect 33318 45568 33324 45620
rect 33376 45608 33382 45620
rect 33962 45608 33968 45620
rect 33376 45580 33968 45608
rect 33376 45568 33382 45580
rect 33962 45568 33968 45580
rect 34020 45568 34026 45620
rect 36078 45568 36084 45620
rect 36136 45608 36142 45620
rect 36136 45580 36407 45608
rect 36136 45568 36142 45580
rect 12434 45500 12440 45552
rect 12492 45540 12498 45552
rect 17678 45540 17684 45552
rect 12492 45512 17684 45540
rect 12492 45500 12498 45512
rect 17678 45500 17684 45512
rect 17736 45500 17742 45552
rect 26344 45512 26832 45540
rect 7374 45432 7380 45484
rect 7432 45472 7438 45484
rect 8205 45475 8263 45481
rect 8205 45472 8217 45475
rect 7432 45444 8217 45472
rect 7432 45432 7438 45444
rect 8205 45441 8217 45444
rect 8251 45441 8263 45475
rect 8205 45435 8263 45441
rect 18690 45432 18696 45484
rect 18748 45472 18754 45484
rect 21726 45472 21732 45484
rect 18748 45444 21732 45472
rect 18748 45432 18754 45444
rect 21726 45432 21732 45444
rect 21784 45432 21790 45484
rect 7282 45364 7288 45416
rect 7340 45404 7346 45416
rect 7561 45407 7619 45413
rect 7561 45404 7573 45407
rect 7340 45376 7573 45404
rect 7340 45364 7346 45376
rect 7561 45373 7573 45376
rect 7607 45373 7619 45407
rect 7561 45367 7619 45373
rect 8389 45407 8447 45413
rect 8389 45373 8401 45407
rect 8435 45404 8447 45407
rect 9398 45404 9404 45416
rect 8435 45376 9404 45404
rect 8435 45373 8447 45376
rect 8389 45367 8447 45373
rect 9398 45364 9404 45376
rect 9456 45364 9462 45416
rect 9490 45364 9496 45416
rect 9548 45404 9554 45416
rect 9677 45407 9735 45413
rect 9548 45376 9593 45404
rect 9548 45364 9554 45376
rect 9677 45373 9689 45407
rect 9723 45404 9735 45407
rect 9950 45404 9956 45416
rect 9723 45376 9956 45404
rect 9723 45373 9735 45376
rect 9677 45367 9735 45373
rect 9950 45364 9956 45376
rect 10008 45364 10014 45416
rect 26344 45413 26372 45512
rect 26329 45407 26387 45413
rect 26329 45373 26341 45407
rect 26375 45373 26387 45407
rect 26329 45367 26387 45373
rect 26418 45364 26424 45416
rect 26476 45404 26482 45416
rect 26702 45407 26760 45413
rect 26702 45404 26714 45407
rect 26476 45376 26714 45404
rect 26476 45364 26482 45376
rect 26702 45373 26714 45376
rect 26748 45373 26760 45407
rect 26804 45404 26832 45512
rect 28534 45500 28540 45552
rect 28592 45540 28598 45552
rect 35710 45540 35716 45552
rect 28592 45512 35716 45540
rect 28592 45500 28598 45512
rect 35710 45500 35716 45512
rect 35768 45500 35774 45552
rect 35989 45543 36047 45549
rect 35989 45509 36001 45543
rect 36035 45540 36047 45543
rect 36262 45540 36268 45552
rect 36035 45512 36268 45540
rect 36035 45509 36047 45512
rect 35989 45503 36047 45509
rect 36262 45500 36268 45512
rect 36320 45500 36326 45552
rect 28534 45404 28540 45416
rect 26804 45376 28540 45404
rect 26702 45367 26760 45373
rect 28534 45364 28540 45376
rect 28592 45364 28598 45416
rect 35802 45404 35808 45416
rect 35763 45376 35808 45404
rect 35802 45364 35808 45376
rect 35860 45364 35866 45416
rect 36379 45404 36407 45580
rect 37182 45568 37188 45620
rect 37240 45608 37246 45620
rect 37240 45580 37320 45608
rect 37240 45568 37246 45580
rect 36538 45500 36544 45552
rect 36596 45500 36602 45552
rect 36556 45472 36584 45500
rect 36556 45444 36768 45472
rect 36740 45413 36768 45444
rect 36814 45432 36820 45484
rect 36872 45472 36878 45484
rect 37182 45472 37188 45484
rect 36872 45444 37188 45472
rect 36872 45432 36878 45444
rect 37182 45432 37188 45444
rect 37240 45432 37246 45484
rect 36449 45407 36507 45413
rect 36449 45404 36461 45407
rect 36379 45376 36461 45404
rect 36449 45373 36461 45376
rect 36495 45373 36507 45407
rect 36449 45367 36507 45373
rect 36542 45407 36600 45413
rect 36542 45373 36554 45407
rect 36588 45373 36600 45407
rect 36542 45367 36600 45373
rect 36725 45407 36783 45413
rect 36725 45373 36737 45407
rect 36771 45373 36783 45407
rect 36725 45367 36783 45373
rect 36955 45407 37013 45413
rect 36955 45373 36967 45407
rect 37001 45404 37013 45407
rect 37292 45404 37320 45580
rect 37734 45568 37740 45620
rect 37792 45608 37798 45620
rect 37829 45611 37887 45617
rect 37829 45608 37841 45611
rect 37792 45580 37841 45608
rect 37792 45568 37798 45580
rect 37829 45577 37841 45580
rect 37875 45608 37887 45611
rect 38286 45608 38292 45620
rect 37875 45580 38292 45608
rect 37875 45577 37887 45580
rect 37829 45571 37887 45577
rect 38286 45568 38292 45580
rect 38344 45568 38350 45620
rect 37001 45376 37320 45404
rect 37737 45407 37795 45413
rect 37001 45373 37013 45376
rect 36955 45367 37013 45373
rect 37737 45373 37749 45407
rect 37783 45404 37795 45407
rect 38194 45404 38200 45416
rect 37783 45376 38200 45404
rect 37783 45373 37795 45376
rect 37737 45367 37795 45373
rect 17494 45296 17500 45348
rect 17552 45336 17558 45348
rect 21726 45336 21732 45348
rect 17552 45308 21732 45336
rect 17552 45296 17558 45308
rect 21726 45296 21732 45308
rect 21784 45296 21790 45348
rect 26510 45336 26516 45348
rect 26471 45308 26516 45336
rect 26510 45296 26516 45308
rect 26568 45296 26574 45348
rect 26605 45339 26663 45345
rect 26605 45305 26617 45339
rect 26651 45305 26663 45339
rect 26605 45299 26663 45305
rect 26898 45339 26956 45345
rect 26898 45305 26910 45339
rect 26944 45336 26956 45339
rect 27430 45336 27436 45348
rect 26944 45308 27436 45336
rect 26944 45305 26956 45308
rect 26898 45299 26956 45305
rect 8573 45271 8631 45277
rect 8573 45237 8585 45271
rect 8619 45268 8631 45271
rect 8662 45268 8668 45280
rect 8619 45240 8668 45268
rect 8619 45237 8631 45240
rect 8573 45231 8631 45237
rect 8662 45228 8668 45240
rect 8720 45228 8726 45280
rect 9861 45271 9919 45277
rect 9861 45237 9873 45271
rect 9907 45268 9919 45271
rect 15838 45268 15844 45280
rect 9907 45240 15844 45268
rect 9907 45237 9919 45240
rect 9861 45231 9919 45237
rect 15838 45228 15844 45240
rect 15896 45228 15902 45280
rect 26234 45228 26240 45280
rect 26292 45268 26298 45280
rect 26620 45268 26648 45299
rect 27430 45296 27436 45308
rect 27488 45296 27494 45348
rect 31570 45296 31576 45348
rect 31628 45336 31634 45348
rect 31628 45308 36124 45336
rect 31628 45296 31634 45308
rect 26292 45240 26648 45268
rect 36096 45268 36124 45308
rect 36262 45296 36268 45348
rect 36320 45336 36326 45348
rect 36556 45336 36584 45367
rect 36814 45336 36820 45348
rect 36320 45308 36584 45336
rect 36775 45308 36820 45336
rect 36320 45296 36326 45308
rect 36814 45296 36820 45308
rect 36872 45296 36878 45348
rect 37752 45280 37780 45367
rect 38194 45364 38200 45376
rect 38252 45404 38258 45416
rect 39390 45404 39396 45416
rect 38252 45376 39396 45404
rect 38252 45364 38258 45376
rect 39390 45364 39396 45376
rect 39448 45364 39454 45416
rect 37093 45271 37151 45277
rect 37093 45268 37105 45271
rect 36096 45240 37105 45268
rect 26292 45228 26298 45240
rect 37093 45237 37105 45240
rect 37139 45237 37151 45271
rect 37093 45231 37151 45237
rect 37734 45228 37740 45280
rect 37792 45228 37798 45280
rect 1104 45178 38824 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 38824 45178
rect 1104 45104 38824 45126
rect 6362 45024 6368 45076
rect 6420 45064 6426 45076
rect 6420 45036 9720 45064
rect 6420 45024 6426 45036
rect 1854 44996 1860 45008
rect 1815 44968 1860 44996
rect 1854 44956 1860 44968
rect 1912 44956 1918 45008
rect 2041 44999 2099 45005
rect 2041 44965 2053 44999
rect 2087 44996 2099 44999
rect 2314 44996 2320 45008
rect 2087 44968 2320 44996
rect 2087 44965 2099 44968
rect 2041 44959 2099 44965
rect 2314 44956 2320 44968
rect 2372 44956 2378 45008
rect 3510 44956 3516 45008
rect 3568 44996 3574 45008
rect 3568 44968 8892 44996
rect 3568 44956 3574 44968
rect 2222 44888 2228 44940
rect 2280 44928 2286 44940
rect 8864 44937 8892 44968
rect 9692 44937 9720 45036
rect 23474 45024 23480 45076
rect 23532 45064 23538 45076
rect 24213 45067 24271 45073
rect 24213 45064 24225 45067
rect 23532 45036 24225 45064
rect 23532 45024 23538 45036
rect 24213 45033 24225 45036
rect 24259 45064 24271 45067
rect 24394 45064 24400 45076
rect 24259 45036 24400 45064
rect 24259 45033 24271 45036
rect 24213 45027 24271 45033
rect 24394 45024 24400 45036
rect 24452 45024 24458 45076
rect 27430 45024 27436 45076
rect 27488 45064 27494 45076
rect 28810 45064 28816 45076
rect 27488 45036 28816 45064
rect 27488 45024 27494 45036
rect 28810 45024 28816 45036
rect 28868 45024 28874 45076
rect 29086 45024 29092 45076
rect 29144 45064 29150 45076
rect 29730 45064 29736 45076
rect 29144 45036 29736 45064
rect 29144 45024 29150 45036
rect 29730 45024 29736 45036
rect 29788 45024 29794 45076
rect 34514 45024 34520 45076
rect 34572 45064 34578 45076
rect 34701 45067 34759 45073
rect 34701 45064 34713 45067
rect 34572 45036 34713 45064
rect 34572 45024 34578 45036
rect 34701 45033 34713 45036
rect 34747 45033 34759 45067
rect 34701 45027 34759 45033
rect 35345 45067 35403 45073
rect 35345 45033 35357 45067
rect 35391 45064 35403 45067
rect 37734 45064 37740 45076
rect 35391 45036 37740 45064
rect 35391 45033 35403 45036
rect 35345 45027 35403 45033
rect 37734 45024 37740 45036
rect 37792 45024 37798 45076
rect 26881 44999 26939 45005
rect 26881 44965 26893 44999
rect 26927 44996 26939 44999
rect 27522 44996 27528 45008
rect 26927 44968 27528 44996
rect 26927 44965 26939 44968
rect 26881 44959 26939 44965
rect 27522 44956 27528 44968
rect 27580 44956 27586 45008
rect 28905 44999 28963 45005
rect 28905 44965 28917 44999
rect 28951 44996 28963 44999
rect 28994 44996 29000 45008
rect 28951 44968 29000 44996
rect 28951 44965 28963 44968
rect 28905 44959 28963 44965
rect 28994 44956 29000 44968
rect 29052 44956 29058 45008
rect 30006 44996 30012 45008
rect 29932 44968 30012 44996
rect 8021 44931 8079 44937
rect 8021 44928 8033 44931
rect 2280 44900 8033 44928
rect 2280 44888 2286 44900
rect 8021 44897 8033 44900
rect 8067 44897 8079 44931
rect 8021 44891 8079 44897
rect 8849 44931 8907 44937
rect 8849 44897 8861 44931
rect 8895 44897 8907 44931
rect 8849 44891 8907 44897
rect 9677 44931 9735 44937
rect 9677 44897 9689 44931
rect 9723 44897 9735 44931
rect 10502 44928 10508 44940
rect 10463 44900 10508 44928
rect 9677 44891 9735 44897
rect 10502 44888 10508 44900
rect 10560 44888 10566 44940
rect 11146 44888 11152 44940
rect 11204 44928 11210 44940
rect 23014 44928 23020 44940
rect 11204 44900 23020 44928
rect 11204 44888 11210 44900
rect 23014 44888 23020 44900
rect 23072 44888 23078 44940
rect 24026 44928 24032 44940
rect 23987 44900 24032 44928
rect 24026 44888 24032 44900
rect 24084 44888 24090 44940
rect 26602 44888 26608 44940
rect 26660 44928 26666 44940
rect 29932 44937 29960 44968
rect 30006 44956 30012 44968
rect 30064 44956 30070 45008
rect 36078 44956 36084 45008
rect 36136 44956 36142 45008
rect 26697 44931 26755 44937
rect 26697 44928 26709 44931
rect 26660 44900 26709 44928
rect 26660 44888 26666 44900
rect 26697 44897 26709 44900
rect 26743 44897 26755 44931
rect 29733 44931 29791 44937
rect 29733 44928 29745 44931
rect 26697 44891 26755 44897
rect 27586 44900 29745 44928
rect 7837 44863 7895 44869
rect 7837 44829 7849 44863
rect 7883 44860 7895 44863
rect 8665 44863 8723 44869
rect 8665 44860 8677 44863
rect 7883 44832 8677 44860
rect 7883 44829 7895 44832
rect 7837 44823 7895 44829
rect 8665 44829 8677 44832
rect 8711 44860 8723 44863
rect 9490 44860 9496 44872
rect 8711 44832 9496 44860
rect 8711 44829 8723 44832
rect 8665 44823 8723 44829
rect 9490 44820 9496 44832
rect 9548 44860 9554 44872
rect 10321 44863 10379 44869
rect 10321 44860 10333 44863
rect 9548 44832 10333 44860
rect 9548 44820 9554 44832
rect 10321 44829 10333 44832
rect 10367 44829 10379 44863
rect 10321 44823 10379 44829
rect 22186 44820 22192 44872
rect 22244 44860 22250 44872
rect 24044 44860 24072 44888
rect 22244 44832 24072 44860
rect 22244 44820 22250 44832
rect 24486 44820 24492 44872
rect 24544 44860 24550 44872
rect 27586 44860 27614 44900
rect 29733 44897 29745 44900
rect 29779 44897 29791 44931
rect 29733 44891 29791 44897
rect 29917 44931 29975 44937
rect 29917 44897 29929 44931
rect 29963 44897 29975 44931
rect 29917 44891 29975 44897
rect 30193 44931 30251 44937
rect 30193 44897 30205 44931
rect 30239 44928 30251 44931
rect 30282 44928 30288 44940
rect 30239 44900 30288 44928
rect 30239 44897 30251 44900
rect 30193 44891 30251 44897
rect 30282 44888 30288 44900
rect 30340 44888 30346 44940
rect 34514 44928 34520 44940
rect 34475 44900 34520 44928
rect 34514 44888 34520 44900
rect 34572 44888 34578 44940
rect 35161 44931 35219 44937
rect 35161 44897 35173 44931
rect 35207 44897 35219 44931
rect 35161 44891 35219 44897
rect 24544 44832 27614 44860
rect 24544 44820 24550 44832
rect 29178 44820 29184 44872
rect 29236 44860 29242 44872
rect 29825 44863 29883 44869
rect 29825 44860 29837 44863
rect 29236 44832 29837 44860
rect 29236 44820 29242 44832
rect 29825 44829 29837 44832
rect 29871 44829 29883 44863
rect 29825 44823 29883 44829
rect 30009 44863 30067 44869
rect 30009 44829 30021 44863
rect 30055 44860 30067 44863
rect 35176 44860 35204 44891
rect 35250 44888 35256 44940
rect 35308 44928 35314 44940
rect 35802 44928 35808 44940
rect 35308 44900 35808 44928
rect 35308 44888 35314 44900
rect 35802 44888 35808 44900
rect 35860 44888 35866 44940
rect 36096 44928 36124 44956
rect 36449 44931 36507 44937
rect 36449 44928 36461 44931
rect 36096 44900 36461 44928
rect 36449 44897 36461 44900
rect 36495 44897 36507 44931
rect 36449 44891 36507 44897
rect 36542 44931 36600 44937
rect 36542 44897 36554 44931
rect 36588 44897 36600 44931
rect 36542 44891 36600 44897
rect 36725 44931 36783 44937
rect 36725 44897 36737 44931
rect 36771 44897 36783 44931
rect 36725 44891 36783 44897
rect 35710 44860 35716 44872
rect 30055 44832 30236 44860
rect 35176 44832 35716 44860
rect 30055 44829 30067 44832
rect 30009 44823 30067 44829
rect 30208 44804 30236 44832
rect 35710 44820 35716 44832
rect 35768 44820 35774 44872
rect 36078 44820 36084 44872
rect 36136 44860 36142 44872
rect 36557 44860 36585 44891
rect 36136 44832 36585 44860
rect 36136 44820 36142 44832
rect 9861 44795 9919 44801
rect 9861 44761 9873 44795
rect 9907 44792 9919 44795
rect 11882 44792 11888 44804
rect 9907 44764 11888 44792
rect 9907 44761 9919 44764
rect 9861 44755 9919 44761
rect 11882 44752 11888 44764
rect 11940 44752 11946 44804
rect 28810 44752 28816 44804
rect 28868 44792 28874 44804
rect 28868 44764 30144 44792
rect 28868 44752 28874 44764
rect 8110 44684 8116 44736
rect 8168 44724 8174 44736
rect 8205 44727 8263 44733
rect 8205 44724 8217 44727
rect 8168 44696 8217 44724
rect 8168 44684 8174 44696
rect 8205 44693 8217 44696
rect 8251 44693 8263 44727
rect 9030 44724 9036 44736
rect 8991 44696 9036 44724
rect 8205 44687 8263 44693
rect 9030 44684 9036 44696
rect 9088 44684 9094 44736
rect 10686 44724 10692 44736
rect 10647 44696 10692 44724
rect 10686 44684 10692 44696
rect 10744 44684 10750 44736
rect 27522 44684 27528 44736
rect 27580 44724 27586 44736
rect 28997 44727 29055 44733
rect 28997 44724 29009 44727
rect 27580 44696 29009 44724
rect 27580 44684 27586 44696
rect 28997 44693 29009 44696
rect 29043 44693 29055 44727
rect 29546 44724 29552 44736
rect 29507 44696 29552 44724
rect 28997 44687 29055 44693
rect 29546 44684 29552 44696
rect 29604 44684 29610 44736
rect 30116 44724 30144 44764
rect 30190 44752 30196 44804
rect 30248 44752 30254 44804
rect 30383 44764 36124 44792
rect 30383 44724 30411 44764
rect 35986 44724 35992 44736
rect 30116 44696 30411 44724
rect 35947 44696 35992 44724
rect 35986 44684 35992 44696
rect 36044 44684 36050 44736
rect 36096 44724 36124 44764
rect 36538 44752 36544 44804
rect 36596 44792 36602 44804
rect 36740 44792 36768 44891
rect 36814 44888 36820 44940
rect 36872 44928 36878 44940
rect 36955 44931 37013 44937
rect 36872 44900 36917 44928
rect 36872 44888 36878 44900
rect 36955 44897 36967 44931
rect 37001 44928 37013 44931
rect 38010 44928 38016 44940
rect 37001 44900 38016 44928
rect 37001 44897 37013 44900
rect 36955 44891 37013 44897
rect 38010 44888 38016 44900
rect 38068 44888 38074 44940
rect 36596 44764 36768 44792
rect 36596 44752 36602 44764
rect 37093 44727 37151 44733
rect 37093 44724 37105 44727
rect 36096 44696 37105 44724
rect 37093 44693 37105 44696
rect 37139 44693 37151 44727
rect 37093 44687 37151 44693
rect 1104 44634 38824 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 38824 44634
rect 1104 44560 38824 44582
rect 15102 44480 15108 44532
rect 15160 44520 15166 44532
rect 26418 44520 26424 44532
rect 15160 44492 26424 44520
rect 15160 44480 15166 44492
rect 26418 44480 26424 44492
rect 26476 44480 26482 44532
rect 26786 44480 26792 44532
rect 26844 44520 26850 44532
rect 26973 44523 27031 44529
rect 26973 44520 26985 44523
rect 26844 44492 26985 44520
rect 26844 44480 26850 44492
rect 26973 44489 26985 44492
rect 27019 44489 27031 44523
rect 32950 44520 32956 44532
rect 26973 44483 27031 44489
rect 29196 44492 32956 44520
rect 2041 44455 2099 44461
rect 2041 44421 2053 44455
rect 2087 44452 2099 44455
rect 2130 44452 2136 44464
rect 2087 44424 2136 44452
rect 2087 44421 2099 44424
rect 2041 44415 2099 44421
rect 2130 44412 2136 44424
rect 2188 44412 2194 44464
rect 29196 44461 29224 44492
rect 32950 44480 32956 44492
rect 33008 44480 33014 44532
rect 34606 44520 34612 44532
rect 34567 44492 34612 44520
rect 34606 44480 34612 44492
rect 34664 44480 34670 44532
rect 35897 44523 35955 44529
rect 35897 44489 35909 44523
rect 35943 44520 35955 44523
rect 37182 44520 37188 44532
rect 35943 44492 37188 44520
rect 35943 44489 35955 44492
rect 35897 44483 35955 44489
rect 37182 44480 37188 44492
rect 37240 44480 37246 44532
rect 29181 44455 29239 44461
rect 29181 44421 29193 44455
rect 29227 44421 29239 44455
rect 29181 44415 29239 44421
rect 36446 44412 36452 44464
rect 36504 44412 36510 44464
rect 36906 44412 36912 44464
rect 36964 44452 36970 44464
rect 38105 44455 38163 44461
rect 38105 44452 38117 44455
rect 36964 44424 38117 44452
rect 36964 44412 36970 44424
rect 38105 44421 38117 44424
rect 38151 44421 38163 44455
rect 38105 44415 38163 44421
rect 6546 44344 6552 44396
rect 6604 44384 6610 44396
rect 9493 44387 9551 44393
rect 9493 44384 9505 44387
rect 6604 44356 7604 44384
rect 6604 44344 6610 44356
rect 1854 44316 1860 44328
rect 1815 44288 1860 44316
rect 1854 44276 1860 44288
rect 1912 44276 1918 44328
rect 7374 44316 7380 44328
rect 7335 44288 7380 44316
rect 7374 44276 7380 44288
rect 7432 44276 7438 44328
rect 7576 44325 7604 44356
rect 8220 44356 9505 44384
rect 8220 44328 8248 44356
rect 9493 44353 9505 44356
rect 9539 44353 9551 44387
rect 9493 44347 9551 44353
rect 9858 44344 9864 44396
rect 9916 44384 9922 44396
rect 17586 44384 17592 44396
rect 9916 44356 17592 44384
rect 9916 44344 9922 44356
rect 17586 44344 17592 44356
rect 17644 44344 17650 44396
rect 19242 44344 19248 44396
rect 19300 44384 19306 44396
rect 33318 44384 33324 44396
rect 19300 44356 33324 44384
rect 19300 44344 19306 44356
rect 33318 44344 33324 44356
rect 33376 44344 33382 44396
rect 7561 44319 7619 44325
rect 7561 44285 7573 44319
rect 7607 44285 7619 44319
rect 8202 44316 8208 44328
rect 8115 44288 8208 44316
rect 7561 44279 7619 44285
rect 7392 44248 7420 44276
rect 8128 44248 8156 44288
rect 8202 44276 8208 44288
rect 8260 44276 8266 44328
rect 8389 44319 8447 44325
rect 8389 44285 8401 44319
rect 8435 44316 8447 44319
rect 8754 44316 8760 44328
rect 8435 44288 8760 44316
rect 8435 44285 8447 44288
rect 8389 44279 8447 44285
rect 8754 44276 8760 44288
rect 8812 44276 8818 44328
rect 9677 44319 9735 44325
rect 9677 44285 9689 44319
rect 9723 44316 9735 44319
rect 10134 44316 10140 44328
rect 9723 44288 10140 44316
rect 9723 44285 9735 44288
rect 9677 44279 9735 44285
rect 10134 44276 10140 44288
rect 10192 44276 10198 44328
rect 22278 44276 22284 44328
rect 22336 44316 22342 44328
rect 29089 44319 29147 44325
rect 29089 44316 29101 44319
rect 22336 44288 29101 44316
rect 22336 44276 22342 44288
rect 29089 44285 29101 44288
rect 29135 44285 29147 44319
rect 29089 44279 29147 44285
rect 29273 44319 29331 44325
rect 29273 44285 29285 44319
rect 29319 44285 29331 44319
rect 29273 44279 29331 44285
rect 29365 44319 29423 44325
rect 29365 44285 29377 44319
rect 29411 44285 29423 44319
rect 29365 44279 29423 44285
rect 29549 44319 29607 44325
rect 29549 44285 29561 44319
rect 29595 44316 29607 44319
rect 30282 44316 30288 44328
rect 29595 44288 30288 44316
rect 29595 44285 29607 44288
rect 29549 44279 29607 44285
rect 7392 44220 8156 44248
rect 8573 44251 8631 44257
rect 8573 44217 8585 44251
rect 8619 44248 8631 44251
rect 13446 44248 13452 44260
rect 8619 44220 13452 44248
rect 8619 44217 8631 44220
rect 8573 44211 8631 44217
rect 13446 44208 13452 44220
rect 13504 44208 13510 44260
rect 26786 44208 26792 44260
rect 26844 44248 26850 44260
rect 26881 44251 26939 44257
rect 26881 44248 26893 44251
rect 26844 44220 26893 44248
rect 26844 44208 26850 44220
rect 26881 44217 26893 44220
rect 26927 44217 26939 44251
rect 26881 44211 26939 44217
rect 28261 44251 28319 44257
rect 28261 44217 28273 44251
rect 28307 44248 28319 44251
rect 29178 44248 29184 44260
rect 28307 44220 29184 44248
rect 28307 44217 28319 44220
rect 28261 44211 28319 44217
rect 29178 44208 29184 44220
rect 29236 44208 29242 44260
rect 1762 44140 1768 44192
rect 1820 44180 1826 44192
rect 5534 44180 5540 44192
rect 1820 44152 5540 44180
rect 1820 44140 1826 44152
rect 5534 44140 5540 44152
rect 5592 44140 5598 44192
rect 7742 44180 7748 44192
rect 7703 44152 7748 44180
rect 7742 44140 7748 44152
rect 7800 44140 7806 44192
rect 9858 44180 9864 44192
rect 9819 44152 9864 44180
rect 9858 44140 9864 44152
rect 9916 44140 9922 44192
rect 27982 44140 27988 44192
rect 28040 44180 28046 44192
rect 28353 44183 28411 44189
rect 28353 44180 28365 44183
rect 28040 44152 28365 44180
rect 28040 44140 28046 44152
rect 28353 44149 28365 44152
rect 28399 44149 28411 44183
rect 28353 44143 28411 44149
rect 28905 44183 28963 44189
rect 28905 44149 28917 44183
rect 28951 44180 28963 44183
rect 28994 44180 29000 44192
rect 28951 44152 29000 44180
rect 28951 44149 28963 44152
rect 28905 44143 28963 44149
rect 28994 44140 29000 44152
rect 29052 44140 29058 44192
rect 29288 44180 29316 44279
rect 29380 44248 29408 44279
rect 30282 44276 30288 44288
rect 30340 44276 30346 44328
rect 34793 44319 34851 44325
rect 34793 44285 34805 44319
rect 34839 44316 34851 44319
rect 35342 44316 35348 44328
rect 34839 44288 35348 44316
rect 34839 44285 34851 44288
rect 34793 44279 34851 44285
rect 35342 44276 35348 44288
rect 35400 44276 35406 44328
rect 36465 44325 36493 44412
rect 37182 44344 37188 44396
rect 37240 44384 37246 44396
rect 37240 44356 37596 44384
rect 37240 44344 37246 44356
rect 37568 44325 37596 44356
rect 36449 44319 36507 44325
rect 36449 44285 36461 44319
rect 36495 44285 36507 44319
rect 36449 44279 36507 44285
rect 36542 44319 36600 44325
rect 36542 44285 36554 44319
rect 36588 44285 36600 44319
rect 36725 44319 36783 44325
rect 36725 44316 36737 44319
rect 36542 44279 36600 44285
rect 36704 44285 36737 44316
rect 36771 44285 36783 44319
rect 36704 44279 36783 44285
rect 36955 44319 37013 44325
rect 36955 44285 36967 44319
rect 37001 44316 37013 44319
rect 37553 44319 37611 44325
rect 37001 44288 37504 44316
rect 37001 44285 37013 44288
rect 36955 44279 37013 44285
rect 30650 44248 30656 44260
rect 29380 44220 30656 44248
rect 30650 44208 30656 44220
rect 30708 44208 30714 44260
rect 35710 44208 35716 44260
rect 35768 44248 35774 44260
rect 35805 44251 35863 44257
rect 35805 44248 35817 44251
rect 35768 44220 35817 44248
rect 35768 44208 35774 44220
rect 35805 44217 35817 44220
rect 35851 44217 35863 44251
rect 35805 44211 35863 44217
rect 35986 44208 35992 44260
rect 36044 44248 36050 44260
rect 36557 44248 36585 44279
rect 36044 44220 36585 44248
rect 36044 44208 36050 44220
rect 31294 44180 31300 44192
rect 29288 44152 31300 44180
rect 31294 44140 31300 44152
rect 31352 44140 31358 44192
rect 35894 44140 35900 44192
rect 35952 44180 35958 44192
rect 36538 44180 36544 44192
rect 35952 44152 36544 44180
rect 35952 44140 35958 44152
rect 36538 44140 36544 44152
rect 36596 44180 36602 44192
rect 36704 44180 36732 44279
rect 36814 44248 36820 44260
rect 36775 44220 36820 44248
rect 36814 44208 36820 44220
rect 36872 44208 36878 44260
rect 36596 44152 36732 44180
rect 37093 44183 37151 44189
rect 36596 44140 36602 44152
rect 37093 44149 37105 44183
rect 37139 44180 37151 44183
rect 37366 44180 37372 44192
rect 37139 44152 37372 44180
rect 37139 44149 37151 44152
rect 37093 44143 37151 44149
rect 37366 44140 37372 44152
rect 37424 44140 37430 44192
rect 37476 44180 37504 44288
rect 37553 44285 37565 44319
rect 37599 44285 37611 44319
rect 37734 44316 37740 44328
rect 37695 44288 37740 44316
rect 37553 44279 37611 44285
rect 37734 44276 37740 44288
rect 37792 44276 37798 44328
rect 37921 44319 37979 44325
rect 37921 44285 37933 44319
rect 37967 44316 37979 44319
rect 38746 44316 38752 44328
rect 37967 44288 38752 44316
rect 37967 44285 37979 44288
rect 37921 44279 37979 44285
rect 38746 44276 38752 44288
rect 38804 44276 38810 44328
rect 37826 44248 37832 44260
rect 37787 44220 37832 44248
rect 37826 44208 37832 44220
rect 37884 44208 37890 44260
rect 38470 44180 38476 44192
rect 37476 44152 38476 44180
rect 38470 44140 38476 44152
rect 38528 44140 38534 44192
rect 1104 44090 38824 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 38824 44090
rect 1104 44016 38824 44038
rect 1946 43936 1952 43988
rect 2004 43976 2010 43988
rect 9217 43979 9275 43985
rect 2004 43948 6914 43976
rect 2004 43936 2010 43948
rect 6886 43908 6914 43948
rect 9217 43945 9229 43979
rect 9263 43976 9275 43979
rect 9490 43976 9496 43988
rect 9263 43948 9496 43976
rect 9263 43945 9275 43948
rect 9217 43939 9275 43945
rect 9490 43936 9496 43948
rect 9548 43936 9554 43988
rect 29273 43979 29331 43985
rect 29273 43945 29285 43979
rect 29319 43976 29331 43979
rect 34146 43976 34152 43988
rect 29319 43948 34152 43976
rect 29319 43945 29331 43948
rect 29273 43939 29331 43945
rect 34146 43936 34152 43948
rect 34204 43936 34210 43988
rect 34330 43936 34336 43988
rect 34388 43976 34394 43988
rect 35253 43979 35311 43985
rect 35253 43976 35265 43979
rect 34388 43948 35265 43976
rect 34388 43936 34394 43948
rect 35253 43945 35265 43948
rect 35299 43945 35311 43979
rect 35253 43939 35311 43945
rect 35894 43936 35900 43988
rect 35952 43976 35958 43988
rect 35952 43948 36492 43976
rect 35952 43936 35958 43948
rect 9582 43908 9588 43920
rect 6886 43880 9588 43908
rect 9582 43868 9588 43880
rect 9640 43868 9646 43920
rect 22002 43868 22008 43920
rect 22060 43908 22066 43920
rect 35342 43908 35348 43920
rect 22060 43880 35348 43908
rect 22060 43868 22066 43880
rect 35342 43868 35348 43880
rect 35400 43868 35406 43920
rect 36464 43908 36492 43948
rect 36538 43936 36544 43988
rect 36596 43976 36602 43988
rect 37001 43979 37059 43985
rect 36596 43948 36865 43976
rect 36596 43936 36602 43948
rect 36633 43911 36691 43917
rect 36633 43908 36645 43911
rect 36188 43880 36400 43908
rect 36464 43880 36645 43908
rect 8202 43840 8208 43852
rect 8163 43812 8208 43840
rect 8202 43800 8208 43812
rect 8260 43800 8266 43852
rect 8389 43843 8447 43849
rect 8389 43809 8401 43843
rect 8435 43840 8447 43843
rect 8478 43840 8484 43852
rect 8435 43812 8484 43840
rect 8435 43809 8447 43812
rect 8389 43803 8447 43809
rect 8478 43800 8484 43812
rect 8536 43800 8542 43852
rect 9033 43843 9091 43849
rect 9033 43809 9045 43843
rect 9079 43809 9091 43843
rect 9033 43803 9091 43809
rect 7282 43732 7288 43784
rect 7340 43772 7346 43784
rect 9048 43772 9076 43803
rect 29178 43800 29184 43852
rect 29236 43840 29242 43852
rect 29549 43843 29607 43849
rect 29549 43840 29561 43843
rect 29236 43812 29561 43840
rect 29236 43800 29242 43812
rect 29549 43809 29561 43812
rect 29595 43809 29607 43843
rect 29549 43803 29607 43809
rect 29825 43843 29883 43849
rect 29825 43809 29837 43843
rect 29871 43840 29883 43843
rect 30021 43843 30079 43849
rect 29871 43812 29960 43840
rect 29871 43809 29883 43812
rect 29825 43803 29883 43809
rect 7340 43744 9076 43772
rect 29742 43775 29800 43781
rect 7340 43732 7346 43744
rect 8220 43716 8248 43744
rect 29742 43741 29754 43775
rect 29788 43741 29800 43775
rect 29932 43772 29960 43812
rect 30021 43809 30033 43843
rect 30067 43840 30079 43843
rect 30282 43840 30288 43852
rect 30067 43812 30288 43840
rect 30067 43809 30079 43812
rect 30021 43803 30079 43809
rect 30282 43800 30288 43812
rect 30340 43800 30346 43852
rect 30374 43800 30380 43852
rect 30432 43840 30438 43852
rect 31294 43840 31300 43852
rect 30432 43812 31300 43840
rect 30432 43800 30438 43812
rect 31294 43800 31300 43812
rect 31352 43800 31358 43852
rect 35066 43840 35072 43852
rect 35027 43812 35072 43840
rect 35066 43800 35072 43812
rect 35124 43800 35130 43852
rect 35802 43800 35808 43852
rect 35860 43840 35866 43852
rect 35897 43843 35955 43849
rect 35897 43840 35909 43843
rect 35860 43812 35909 43840
rect 35860 43800 35866 43812
rect 35897 43809 35909 43812
rect 35943 43809 35955 43843
rect 35897 43803 35955 43809
rect 31478 43772 31484 43784
rect 29932 43744 31484 43772
rect 29742 43735 29800 43741
rect 8202 43664 8208 43716
rect 8260 43664 8266 43716
rect 29273 43707 29331 43713
rect 29273 43673 29285 43707
rect 29319 43704 29331 43707
rect 29641 43707 29699 43713
rect 29641 43704 29653 43707
rect 29319 43676 29653 43704
rect 29319 43673 29331 43676
rect 29273 43667 29331 43673
rect 29641 43673 29653 43676
rect 29687 43673 29699 43707
rect 29748 43704 29776 43735
rect 31478 43732 31484 43744
rect 31536 43732 31542 43784
rect 31110 43704 31116 43716
rect 29748 43676 31116 43704
rect 29641 43667 29699 43673
rect 31110 43664 31116 43676
rect 31168 43664 31174 43716
rect 36188 43704 36216 43880
rect 36372 43849 36400 43880
rect 36633 43877 36645 43880
rect 36679 43877 36691 43911
rect 36633 43871 36691 43877
rect 36538 43849 36544 43852
rect 36357 43843 36415 43849
rect 36357 43809 36369 43843
rect 36403 43809 36415 43843
rect 36357 43803 36415 43809
rect 36505 43843 36544 43849
rect 36505 43809 36517 43843
rect 36505 43803 36544 43809
rect 36538 43800 36544 43803
rect 36596 43800 36602 43852
rect 36837 43849 36865 43948
rect 37001 43945 37013 43979
rect 37047 43945 37059 43979
rect 37001 43939 37059 43945
rect 37016 43908 37044 43939
rect 37182 43936 37188 43988
rect 37240 43976 37246 43988
rect 37550 43976 37556 43988
rect 37240 43948 37556 43976
rect 37240 43936 37246 43948
rect 37550 43936 37556 43948
rect 37608 43936 37614 43988
rect 38102 43908 38108 43920
rect 37016 43880 38108 43908
rect 38102 43868 38108 43880
rect 38160 43868 38166 43920
rect 36725 43843 36783 43849
rect 36725 43809 36737 43843
rect 36771 43809 36783 43843
rect 36725 43803 36783 43809
rect 36822 43843 36880 43849
rect 36822 43809 36834 43843
rect 36868 43809 36880 43843
rect 36822 43803 36880 43809
rect 36740 43772 36768 43803
rect 37550 43772 37556 43784
rect 36740 43744 37556 43772
rect 37550 43732 37556 43744
rect 37608 43732 37614 43784
rect 37274 43704 37280 43716
rect 36188 43676 37280 43704
rect 37274 43664 37280 43676
rect 37332 43664 37338 43716
rect 8570 43636 8576 43648
rect 8531 43608 8576 43636
rect 8570 43596 8576 43608
rect 8628 43596 8634 43648
rect 29365 43639 29423 43645
rect 29365 43605 29377 43639
rect 29411 43636 29423 43639
rect 30374 43636 30380 43648
rect 29411 43608 30380 43636
rect 29411 43605 29423 43608
rect 29365 43599 29423 43605
rect 30374 43596 30380 43608
rect 30432 43596 30438 43648
rect 35713 43639 35771 43645
rect 35713 43605 35725 43639
rect 35759 43636 35771 43639
rect 39022 43636 39028 43648
rect 35759 43608 39028 43636
rect 35759 43605 35771 43608
rect 35713 43599 35771 43605
rect 39022 43596 39028 43608
rect 39080 43596 39086 43648
rect 1104 43546 38824 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 38824 43546
rect 1104 43472 38824 43494
rect 2038 43392 2044 43444
rect 2096 43432 2102 43444
rect 20714 43432 20720 43444
rect 2096 43404 20720 43432
rect 2096 43392 2102 43404
rect 20714 43392 20720 43404
rect 20772 43392 20778 43444
rect 27065 43435 27123 43441
rect 27065 43401 27077 43435
rect 27111 43432 27123 43435
rect 28626 43432 28632 43444
rect 27111 43404 28632 43432
rect 27111 43401 27123 43404
rect 27065 43395 27123 43401
rect 28626 43392 28632 43404
rect 28684 43392 28690 43444
rect 34609 43435 34667 43441
rect 34609 43401 34621 43435
rect 34655 43432 34667 43435
rect 36722 43432 36728 43444
rect 34655 43404 36728 43432
rect 34655 43401 34667 43404
rect 34609 43395 34667 43401
rect 36722 43392 36728 43404
rect 36780 43392 36786 43444
rect 36817 43435 36875 43441
rect 36817 43401 36829 43435
rect 36863 43432 36875 43435
rect 36998 43432 37004 43444
rect 36863 43404 37004 43432
rect 36863 43401 36875 43404
rect 36817 43395 36875 43401
rect 36998 43392 37004 43404
rect 37056 43392 37062 43444
rect 26510 43324 26516 43376
rect 26568 43364 26574 43376
rect 27338 43364 27344 43376
rect 26568 43336 27344 43364
rect 26568 43324 26574 43336
rect 27338 43324 27344 43336
rect 27396 43324 27402 43376
rect 34514 43324 34520 43376
rect 34572 43364 34578 43376
rect 36538 43364 36544 43376
rect 34572 43336 36544 43364
rect 34572 43324 34578 43336
rect 36538 43324 36544 43336
rect 36596 43324 36602 43376
rect 2041 43299 2099 43305
rect 2041 43265 2053 43299
rect 2087 43296 2099 43299
rect 2682 43296 2688 43308
rect 2087 43268 2688 43296
rect 2087 43265 2099 43268
rect 2041 43259 2099 43265
rect 2682 43256 2688 43268
rect 2740 43256 2746 43308
rect 19150 43256 19156 43308
rect 19208 43296 19214 43308
rect 19208 43268 37596 43296
rect 19208 43256 19214 43268
rect 1854 43228 1860 43240
rect 1815 43200 1860 43228
rect 1854 43188 1860 43200
rect 1912 43188 1918 43240
rect 2130 43188 2136 43240
rect 2188 43228 2194 43240
rect 26510 43228 26516 43240
rect 2188 43200 6914 43228
rect 26471 43200 26516 43228
rect 2188 43188 2194 43200
rect 6886 43160 6914 43200
rect 26510 43188 26516 43200
rect 26568 43188 26574 43240
rect 26886 43231 26944 43237
rect 26886 43228 26898 43231
rect 26620 43200 26898 43228
rect 26620 43160 26648 43200
rect 26886 43197 26898 43200
rect 26932 43197 26944 43231
rect 26886 43191 26944 43197
rect 28074 43188 28080 43240
rect 28132 43228 28138 43240
rect 29089 43231 29147 43237
rect 29089 43228 29101 43231
rect 28132 43200 29101 43228
rect 28132 43188 28138 43200
rect 29089 43197 29101 43200
rect 29135 43197 29147 43231
rect 29089 43191 29147 43197
rect 29181 43231 29239 43237
rect 29181 43197 29193 43231
rect 29227 43197 29239 43231
rect 29181 43191 29239 43197
rect 29273 43231 29331 43237
rect 29273 43197 29285 43231
rect 29319 43197 29331 43231
rect 29273 43191 29331 43197
rect 29365 43231 29423 43237
rect 29365 43197 29377 43231
rect 29411 43228 29423 43231
rect 29454 43228 29460 43240
rect 29411 43200 29460 43228
rect 29411 43197 29423 43200
rect 29365 43191 29423 43197
rect 6886 43132 26648 43160
rect 26697 43163 26755 43169
rect 26697 43129 26709 43163
rect 26743 43129 26755 43163
rect 26697 43123 26755 43129
rect 26789 43163 26847 43169
rect 26789 43129 26801 43163
rect 26835 43160 26847 43163
rect 27522 43160 27528 43172
rect 26835 43132 27528 43160
rect 26835 43129 26847 43132
rect 26789 43123 26847 43129
rect 25866 43052 25872 43104
rect 25924 43092 25930 43104
rect 26712 43092 26740 43123
rect 27522 43120 27528 43132
rect 27580 43120 27586 43172
rect 27982 43092 27988 43104
rect 25924 43064 27988 43092
rect 25924 43052 25930 43064
rect 27982 43052 27988 43064
rect 28040 43052 28046 43104
rect 28902 43092 28908 43104
rect 28863 43064 28908 43092
rect 28902 43052 28908 43064
rect 28960 43052 28966 43104
rect 29196 43092 29224 43191
rect 29288 43160 29316 43191
rect 29454 43188 29460 43200
rect 29512 43188 29518 43240
rect 29549 43231 29607 43237
rect 29549 43197 29561 43231
rect 29595 43228 29607 43231
rect 30006 43228 30012 43240
rect 29595 43200 30012 43228
rect 29595 43197 29607 43200
rect 29549 43191 29607 43197
rect 30006 43188 30012 43200
rect 30064 43228 30070 43240
rect 30282 43228 30288 43240
rect 30064 43200 30288 43228
rect 30064 43188 30070 43200
rect 30282 43188 30288 43200
rect 30340 43188 30346 43240
rect 34793 43231 34851 43237
rect 34793 43197 34805 43231
rect 34839 43228 34851 43231
rect 34974 43228 34980 43240
rect 34839 43200 34980 43228
rect 34839 43197 34851 43200
rect 34793 43191 34851 43197
rect 34974 43188 34980 43200
rect 35032 43188 35038 43240
rect 35434 43188 35440 43240
rect 35492 43228 35498 43240
rect 35713 43231 35771 43237
rect 35713 43228 35725 43231
rect 35492 43200 35725 43228
rect 35492 43188 35498 43200
rect 35713 43197 35725 43200
rect 35759 43197 35771 43231
rect 37458 43228 37464 43240
rect 35713 43191 35771 43197
rect 35820 43200 37464 43228
rect 32490 43160 32496 43172
rect 29288 43132 32496 43160
rect 32490 43120 32496 43132
rect 32548 43120 32554 43172
rect 34606 43120 34612 43172
rect 34664 43160 34670 43172
rect 35820 43160 35848 43200
rect 37458 43188 37464 43200
rect 37516 43188 37522 43240
rect 37568 43237 37596 43268
rect 37553 43231 37611 43237
rect 37553 43197 37565 43231
rect 37599 43197 37611 43231
rect 37734 43228 37740 43240
rect 37695 43200 37740 43228
rect 37553 43191 37611 43197
rect 37734 43188 37740 43200
rect 37792 43188 37798 43240
rect 37967 43231 38025 43237
rect 37967 43197 37979 43231
rect 38013 43228 38025 43231
rect 39022 43228 39028 43240
rect 38013 43200 39028 43228
rect 38013 43197 38025 43200
rect 37967 43191 38025 43197
rect 39022 43188 39028 43200
rect 39080 43188 39086 43240
rect 34664 43132 35848 43160
rect 36725 43163 36783 43169
rect 34664 43120 34670 43132
rect 36725 43129 36737 43163
rect 36771 43160 36783 43163
rect 37090 43160 37096 43172
rect 36771 43132 37096 43160
rect 36771 43129 36783 43132
rect 36725 43123 36783 43129
rect 37090 43120 37096 43132
rect 37148 43120 37154 43172
rect 37826 43160 37832 43172
rect 37787 43132 37832 43160
rect 37826 43120 37832 43132
rect 37884 43120 37890 43172
rect 33042 43092 33048 43104
rect 29196 43064 33048 43092
rect 33042 43052 33048 43064
rect 33100 43052 33106 43104
rect 35897 43095 35955 43101
rect 35897 43061 35909 43095
rect 35943 43092 35955 43095
rect 37182 43092 37188 43104
rect 35943 43064 37188 43092
rect 35943 43061 35955 43064
rect 35897 43055 35955 43061
rect 37182 43052 37188 43064
rect 37240 43052 37246 43104
rect 38102 43092 38108 43104
rect 38063 43064 38108 43092
rect 38102 43052 38108 43064
rect 38160 43052 38166 43104
rect 1104 43002 38824 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 38824 43002
rect 1104 42928 38824 42950
rect 8478 42848 8484 42900
rect 8536 42888 8542 42900
rect 16022 42888 16028 42900
rect 8536 42860 16028 42888
rect 8536 42848 8542 42860
rect 16022 42848 16028 42860
rect 16080 42848 16086 42900
rect 27338 42848 27344 42900
rect 27396 42888 27402 42900
rect 34146 42888 34152 42900
rect 27396 42860 34152 42888
rect 27396 42848 27402 42860
rect 34146 42848 34152 42860
rect 34204 42848 34210 42900
rect 35342 42848 35348 42900
rect 35400 42848 35406 42900
rect 37734 42888 37740 42900
rect 37016 42860 37740 42888
rect 9030 42780 9036 42832
rect 9088 42820 9094 42832
rect 14734 42820 14740 42832
rect 9088 42792 14740 42820
rect 9088 42780 9094 42792
rect 14734 42780 14740 42792
rect 14792 42780 14798 42832
rect 25866 42780 25872 42832
rect 25924 42820 25930 42832
rect 26421 42823 26479 42829
rect 26421 42820 26433 42823
rect 25924 42792 26433 42820
rect 25924 42780 25930 42792
rect 26421 42789 26433 42792
rect 26467 42789 26479 42823
rect 26421 42783 26479 42789
rect 26513 42823 26571 42829
rect 26513 42789 26525 42823
rect 26559 42820 26571 42823
rect 27522 42820 27528 42832
rect 26559 42792 27528 42820
rect 26559 42789 26571 42792
rect 26513 42783 26571 42789
rect 27522 42780 27528 42792
rect 27580 42780 27586 42832
rect 29270 42780 29276 42832
rect 29328 42780 29334 42832
rect 35360 42820 35388 42848
rect 35360 42792 35572 42820
rect 1854 42752 1860 42764
rect 1815 42724 1860 42752
rect 1854 42712 1860 42724
rect 1912 42712 1918 42764
rect 2038 42752 2044 42764
rect 1999 42724 2044 42752
rect 2038 42712 2044 42724
rect 2096 42712 2102 42764
rect 26237 42755 26295 42761
rect 26237 42721 26249 42755
rect 26283 42721 26295 42755
rect 26237 42715 26295 42721
rect 26633 42755 26691 42761
rect 26633 42721 26645 42755
rect 26679 42721 26691 42755
rect 26633 42715 26691 42721
rect 26806 42755 26864 42761
rect 26806 42721 26818 42755
rect 26852 42752 26864 42755
rect 27062 42752 27068 42764
rect 26852 42724 27068 42752
rect 26852 42721 26864 42724
rect 26806 42715 26864 42721
rect 26252 42684 26280 42715
rect 26510 42684 26516 42696
rect 26252 42656 26516 42684
rect 26510 42644 26516 42656
rect 26568 42644 26574 42696
rect 2038 42576 2044 42628
rect 2096 42616 2102 42628
rect 26648 42616 26676 42715
rect 27062 42712 27068 42724
rect 27120 42712 27126 42764
rect 29288 42752 29316 42780
rect 30282 42752 30288 42764
rect 29288 42724 30288 42752
rect 30282 42712 30288 42724
rect 30340 42712 30346 42764
rect 34885 42755 34943 42761
rect 34885 42721 34897 42755
rect 34931 42752 34943 42755
rect 35342 42752 35348 42764
rect 34931 42724 35348 42752
rect 34931 42721 34943 42724
rect 34885 42715 34943 42721
rect 35342 42712 35348 42724
rect 35400 42712 35406 42764
rect 27338 42644 27344 42696
rect 27396 42684 27402 42696
rect 29270 42684 29276 42696
rect 27396 42656 29276 42684
rect 27396 42644 27402 42656
rect 29270 42644 29276 42656
rect 29328 42644 29334 42696
rect 35544 42684 35572 42792
rect 35710 42752 35716 42764
rect 35671 42724 35716 42752
rect 35710 42712 35716 42724
rect 35768 42712 35774 42764
rect 36173 42755 36231 42761
rect 36173 42721 36185 42755
rect 36219 42721 36231 42755
rect 36173 42715 36231 42721
rect 35544 42656 35756 42684
rect 35728 42628 35756 42656
rect 2096 42588 26676 42616
rect 2096 42576 2102 42588
rect 27890 42576 27896 42628
rect 27948 42616 27954 42628
rect 35069 42619 35127 42625
rect 35069 42616 35081 42619
rect 27948 42588 35081 42616
rect 27948 42576 27954 42588
rect 35069 42585 35081 42588
rect 35115 42585 35127 42619
rect 35069 42579 35127 42585
rect 35529 42619 35587 42625
rect 35529 42585 35541 42619
rect 35575 42616 35587 42619
rect 35618 42616 35624 42628
rect 35575 42588 35624 42616
rect 35575 42585 35587 42588
rect 35529 42579 35587 42585
rect 35618 42576 35624 42588
rect 35676 42576 35682 42628
rect 35710 42576 35716 42628
rect 35768 42576 35774 42628
rect 36188 42616 36216 42715
rect 36354 42712 36360 42764
rect 36412 42752 36418 42764
rect 37016 42761 37044 42860
rect 37734 42848 37740 42860
rect 37792 42848 37798 42900
rect 37093 42823 37151 42829
rect 37093 42789 37105 42823
rect 37139 42820 37151 42823
rect 37826 42820 37832 42832
rect 37139 42792 37832 42820
rect 37139 42789 37151 42792
rect 37093 42783 37151 42789
rect 36817 42755 36875 42761
rect 36817 42752 36829 42755
rect 36412 42724 36829 42752
rect 36412 42712 36418 42724
rect 36817 42721 36829 42724
rect 36863 42721 36875 42755
rect 36817 42715 36875 42721
rect 37001 42755 37059 42761
rect 37001 42721 37013 42755
rect 37047 42721 37059 42755
rect 37001 42715 37059 42721
rect 36722 42616 36728 42628
rect 36188 42588 36728 42616
rect 21910 42508 21916 42560
rect 21968 42548 21974 42560
rect 36188 42548 36216 42588
rect 36722 42576 36728 42588
rect 36780 42576 36786 42628
rect 36814 42576 36820 42628
rect 36872 42616 36878 42628
rect 37108 42616 37136 42783
rect 37826 42780 37832 42792
rect 37884 42780 37890 42832
rect 37274 42761 37280 42764
rect 37231 42755 37280 42761
rect 37231 42721 37243 42755
rect 37277 42721 37280 42755
rect 37231 42715 37280 42721
rect 37274 42712 37280 42715
rect 37332 42712 37338 42764
rect 36872 42588 37136 42616
rect 36872 42576 36878 42588
rect 21968 42520 36216 42548
rect 36357 42551 36415 42557
rect 21968 42508 21974 42520
rect 36357 42517 36369 42551
rect 36403 42548 36415 42551
rect 36538 42548 36544 42560
rect 36403 42520 36544 42548
rect 36403 42517 36415 42520
rect 36357 42511 36415 42517
rect 36538 42508 36544 42520
rect 36596 42508 36602 42560
rect 37274 42508 37280 42560
rect 37332 42548 37338 42560
rect 37369 42551 37427 42557
rect 37369 42548 37381 42551
rect 37332 42520 37381 42548
rect 37332 42508 37338 42520
rect 37369 42517 37381 42520
rect 37415 42517 37427 42551
rect 37369 42511 37427 42517
rect 1104 42458 38824 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 38824 42458
rect 1104 42384 38824 42406
rect 25961 42347 26019 42353
rect 25961 42313 25973 42347
rect 26007 42344 26019 42347
rect 26234 42344 26240 42356
rect 26007 42316 26240 42344
rect 26007 42313 26019 42316
rect 25961 42307 26019 42313
rect 26234 42304 26240 42316
rect 26292 42304 26298 42356
rect 27062 42304 27068 42356
rect 27120 42344 27126 42356
rect 28353 42347 28411 42353
rect 27120 42316 28304 42344
rect 27120 42304 27126 42316
rect 26786 42236 26792 42288
rect 26844 42276 26850 42288
rect 26844 42248 26924 42276
rect 26844 42236 26850 42248
rect 6886 42180 8156 42208
rect 3602 42100 3608 42152
rect 3660 42140 3666 42152
rect 6886 42140 6914 42180
rect 3660 42112 6914 42140
rect 3660 42100 3666 42112
rect 7190 42100 7196 42152
rect 7248 42140 7254 42152
rect 7926 42140 7932 42152
rect 7248 42112 7932 42140
rect 7248 42100 7254 42112
rect 7926 42100 7932 42112
rect 7984 42100 7990 42152
rect 8128 42149 8156 42180
rect 26234 42168 26240 42220
rect 26292 42208 26298 42220
rect 26513 42211 26571 42217
rect 26513 42208 26525 42211
rect 26292 42180 26525 42208
rect 26292 42168 26298 42180
rect 26513 42177 26525 42180
rect 26559 42208 26571 42211
rect 26602 42208 26608 42220
rect 26559 42180 26608 42208
rect 26559 42177 26571 42180
rect 26513 42171 26571 42177
rect 26602 42168 26608 42180
rect 26660 42168 26666 42220
rect 8113 42143 8171 42149
rect 8113 42109 8125 42143
rect 8159 42109 8171 42143
rect 8113 42103 8171 42109
rect 26418 42100 26424 42152
rect 26476 42140 26482 42152
rect 26789 42143 26847 42149
rect 26789 42140 26801 42143
rect 26476 42112 26801 42140
rect 26476 42100 26482 42112
rect 26789 42109 26801 42112
rect 26835 42109 26847 42143
rect 26789 42103 26847 42109
rect 8570 42032 8576 42084
rect 8628 42072 8634 42084
rect 10318 42072 10324 42084
rect 8628 42044 10324 42072
rect 8628 42032 8634 42044
rect 10318 42032 10324 42044
rect 10376 42032 10382 42084
rect 25869 42075 25927 42081
rect 25869 42041 25881 42075
rect 25915 42072 25927 42075
rect 26896 42072 26924 42248
rect 27338 42236 27344 42288
rect 27396 42276 27402 42288
rect 28276 42276 28304 42316
rect 28353 42313 28365 42347
rect 28399 42344 28411 42347
rect 28442 42344 28448 42356
rect 28399 42316 28448 42344
rect 28399 42313 28411 42316
rect 28353 42307 28411 42313
rect 28442 42304 28448 42316
rect 28500 42304 28506 42356
rect 34609 42347 34667 42353
rect 34609 42313 34621 42347
rect 34655 42344 34667 42347
rect 36262 42344 36268 42356
rect 34655 42316 36268 42344
rect 34655 42313 34667 42316
rect 34609 42307 34667 42313
rect 36262 42304 36268 42316
rect 36320 42304 36326 42356
rect 37366 42344 37372 42356
rect 36372 42316 37372 42344
rect 31570 42276 31576 42288
rect 27396 42248 28217 42276
rect 28276 42248 31576 42276
rect 27396 42236 27402 42248
rect 27522 42168 27528 42220
rect 27580 42208 27586 42220
rect 27580 42180 28120 42208
rect 27580 42168 27586 42180
rect 27522 42072 27528 42084
rect 25915 42044 27528 42072
rect 25915 42041 25927 42044
rect 25869 42035 25927 42041
rect 27522 42032 27528 42044
rect 27580 42032 27586 42084
rect 8297 42007 8355 42013
rect 8297 41973 8309 42007
rect 8343 42004 8355 42007
rect 14550 42004 14556 42016
rect 8343 41976 14556 42004
rect 8343 41973 8355 41976
rect 8297 41967 8355 41973
rect 14550 41964 14556 41976
rect 14608 41964 14614 42016
rect 26510 41964 26516 42016
rect 26568 42004 26574 42016
rect 26786 42004 26792 42016
rect 26568 41976 26792 42004
rect 26568 41964 26574 41976
rect 26786 41964 26792 41976
rect 26844 42004 26850 42016
rect 27632 42004 27660 42180
rect 27801 42143 27859 42149
rect 27801 42140 27813 42143
rect 26844 41976 27660 42004
rect 27724 42112 27813 42140
rect 27724 42004 27752 42112
rect 27801 42109 27813 42112
rect 27847 42109 27859 42143
rect 27982 42140 27988 42152
rect 27943 42112 27988 42140
rect 27801 42103 27859 42109
rect 27982 42100 27988 42112
rect 28040 42100 28046 42152
rect 28092 42149 28120 42180
rect 28189 42149 28217 42248
rect 31570 42236 31576 42248
rect 31628 42236 31634 42288
rect 33042 42236 33048 42288
rect 33100 42276 33106 42288
rect 36372 42276 36400 42316
rect 37366 42304 37372 42316
rect 37424 42304 37430 42356
rect 37458 42276 37464 42288
rect 33100 42248 36400 42276
rect 36464 42248 37464 42276
rect 33100 42236 33106 42248
rect 33318 42208 33324 42220
rect 28276 42180 33324 42208
rect 28077 42143 28135 42149
rect 28077 42109 28089 42143
rect 28123 42109 28135 42143
rect 28077 42103 28135 42109
rect 28174 42143 28232 42149
rect 28174 42109 28186 42143
rect 28220 42109 28232 42143
rect 28174 42103 28232 42109
rect 28276 42004 28304 42180
rect 33318 42168 33324 42180
rect 33376 42168 33382 42220
rect 28534 42100 28540 42152
rect 28592 42140 28598 42152
rect 28810 42140 28816 42152
rect 28592 42112 28816 42140
rect 28592 42100 28598 42112
rect 28810 42100 28816 42112
rect 28868 42100 28874 42152
rect 28997 42143 29055 42149
rect 28997 42109 29009 42143
rect 29043 42140 29055 42143
rect 29086 42140 29092 42152
rect 29043 42112 29092 42140
rect 29043 42109 29055 42112
rect 28997 42103 29055 42109
rect 29086 42100 29092 42112
rect 29144 42100 29150 42152
rect 34790 42140 34796 42152
rect 34751 42112 34796 42140
rect 34790 42100 34796 42112
rect 34848 42100 34854 42152
rect 36170 42100 36176 42152
rect 36228 42140 36234 42152
rect 36464 42149 36492 42248
rect 37458 42236 37464 42248
rect 37516 42276 37522 42288
rect 37734 42276 37740 42288
rect 37516 42248 37740 42276
rect 37516 42236 37522 42248
rect 37734 42236 37740 42248
rect 37792 42236 37798 42288
rect 36814 42208 36820 42220
rect 36556 42180 36820 42208
rect 36556 42149 36584 42180
rect 36814 42168 36820 42180
rect 36872 42168 36878 42220
rect 37277 42211 37335 42217
rect 37277 42177 37289 42211
rect 37323 42208 37335 42211
rect 38194 42208 38200 42220
rect 37323 42180 38200 42208
rect 37323 42177 37335 42180
rect 37277 42171 37335 42177
rect 38194 42168 38200 42180
rect 38252 42208 38258 42220
rect 38470 42208 38476 42220
rect 38252 42180 38476 42208
rect 38252 42168 38258 42180
rect 38470 42168 38476 42180
rect 38528 42168 38534 42220
rect 36265 42143 36323 42149
rect 36265 42140 36277 42143
rect 36228 42112 36277 42140
rect 36228 42100 36234 42112
rect 36265 42109 36277 42112
rect 36311 42109 36323 42143
rect 36265 42103 36323 42109
rect 36449 42143 36507 42149
rect 36449 42109 36461 42143
rect 36495 42109 36507 42143
rect 36449 42103 36507 42109
rect 36541 42143 36599 42149
rect 36541 42109 36553 42143
rect 36587 42109 36599 42143
rect 36541 42103 36599 42109
rect 36633 42143 36691 42149
rect 36633 42109 36645 42143
rect 36679 42109 36691 42143
rect 36832 42140 36860 42168
rect 37366 42140 37372 42152
rect 36832 42112 37372 42140
rect 36633 42103 36691 42109
rect 36648 42072 36676 42103
rect 37366 42100 37372 42112
rect 37424 42100 37430 42152
rect 37553 42143 37611 42149
rect 37553 42109 37565 42143
rect 37599 42140 37611 42143
rect 37734 42140 37740 42152
rect 37599 42112 37740 42140
rect 37599 42109 37611 42112
rect 37553 42103 37611 42109
rect 37734 42100 37740 42112
rect 37792 42100 37798 42152
rect 38194 42072 38200 42084
rect 36648 42044 38200 42072
rect 38194 42032 38200 42044
rect 38252 42032 38258 42084
rect 27724 41976 28304 42004
rect 26844 41964 26850 41976
rect 28810 41964 28816 42016
rect 28868 42004 28874 42016
rect 29089 42007 29147 42013
rect 29089 42004 29101 42007
rect 28868 41976 29101 42004
rect 28868 41964 28874 41976
rect 29089 41973 29101 41976
rect 29135 41973 29147 42007
rect 29089 41967 29147 41973
rect 36262 41964 36268 42016
rect 36320 42004 36326 42016
rect 36817 42007 36875 42013
rect 36817 42004 36829 42007
rect 36320 41976 36829 42004
rect 36320 41964 36326 41976
rect 36817 41973 36829 41976
rect 36863 41973 36875 42007
rect 36817 41967 36875 41973
rect 1104 41914 38824 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 38824 41914
rect 1104 41840 38824 41862
rect 2774 41760 2780 41812
rect 2832 41800 2838 41812
rect 27338 41800 27344 41812
rect 2832 41772 27344 41800
rect 2832 41760 2838 41772
rect 27338 41760 27344 41772
rect 27396 41760 27402 41812
rect 31110 41800 31116 41812
rect 27632 41772 31116 41800
rect 1854 41732 1860 41744
rect 1815 41704 1860 41732
rect 1854 41692 1860 41704
rect 1912 41692 1918 41744
rect 5534 41692 5540 41744
rect 5592 41732 5598 41744
rect 5592 41704 8984 41732
rect 5592 41692 5598 41704
rect 5074 41624 5080 41676
rect 5132 41664 5138 41676
rect 8956 41673 8984 41704
rect 9490 41692 9496 41744
rect 9548 41732 9554 41744
rect 22094 41732 22100 41744
rect 9548 41704 22100 41732
rect 9548 41692 9554 41704
rect 22094 41692 22100 41704
rect 22152 41692 22158 41744
rect 25866 41692 25872 41744
rect 25924 41732 25930 41744
rect 26418 41732 26424 41744
rect 25924 41704 26424 41732
rect 25924 41692 25930 41704
rect 26418 41692 26424 41704
rect 26476 41692 26482 41744
rect 8113 41667 8171 41673
rect 8113 41664 8125 41667
rect 5132 41636 8125 41664
rect 5132 41624 5138 41636
rect 8113 41633 8125 41636
rect 8159 41633 8171 41667
rect 8113 41627 8171 41633
rect 8941 41667 8999 41673
rect 8941 41633 8953 41667
rect 8987 41633 8999 41667
rect 8941 41627 8999 41633
rect 20070 41624 20076 41676
rect 20128 41664 20134 41676
rect 26237 41667 26295 41673
rect 20128 41636 20208 41664
rect 20128 41624 20134 41636
rect 7926 41596 7932 41608
rect 7887 41568 7932 41596
rect 7926 41556 7932 41568
rect 7984 41596 7990 41608
rect 8757 41599 8815 41605
rect 8757 41596 8769 41599
rect 7984 41568 8769 41596
rect 7984 41556 7990 41568
rect 8757 41565 8769 41568
rect 8803 41565 8815 41599
rect 15102 41596 15108 41608
rect 8757 41559 8815 41565
rect 8864 41568 15108 41596
rect 2041 41531 2099 41537
rect 2041 41497 2053 41531
rect 2087 41528 2099 41531
rect 2087 41500 8524 41528
rect 2087 41497 2099 41500
rect 2041 41491 2099 41497
rect 8294 41460 8300 41472
rect 8255 41432 8300 41460
rect 8294 41420 8300 41432
rect 8352 41420 8358 41472
rect 8496 41460 8524 41500
rect 8864 41460 8892 41568
rect 15102 41556 15108 41568
rect 15160 41556 15166 41608
rect 20180 41472 20208 41636
rect 26237 41633 26249 41667
rect 26283 41633 26295 41667
rect 26510 41664 26516 41676
rect 26471 41636 26516 41664
rect 26237 41627 26295 41633
rect 26252 41596 26280 41627
rect 26510 41624 26516 41636
rect 26568 41624 26574 41676
rect 26602 41624 26608 41676
rect 26660 41673 26666 41676
rect 26660 41664 26668 41673
rect 26660 41636 26705 41664
rect 26660 41627 26668 41636
rect 26660 41624 26666 41627
rect 27632 41596 27660 41772
rect 31110 41760 31116 41772
rect 31168 41760 31174 41812
rect 34606 41800 34612 41812
rect 34567 41772 34612 41800
rect 34606 41760 34612 41772
rect 34664 41760 34670 41812
rect 35437 41803 35495 41809
rect 35437 41769 35449 41803
rect 35483 41800 35495 41803
rect 35894 41800 35900 41812
rect 35483 41772 35900 41800
rect 35483 41769 35495 41772
rect 35437 41763 35495 41769
rect 35894 41760 35900 41772
rect 35952 41760 35958 41812
rect 36081 41803 36139 41809
rect 36081 41769 36093 41803
rect 36127 41800 36139 41803
rect 37550 41800 37556 41812
rect 36127 41772 37556 41800
rect 36127 41769 36139 41772
rect 36081 41763 36139 41769
rect 37550 41760 37556 41772
rect 37608 41760 37614 41812
rect 27706 41692 27712 41744
rect 27764 41732 27770 41744
rect 27982 41732 27988 41744
rect 27764 41704 27988 41732
rect 27764 41692 27770 41704
rect 27982 41692 27988 41704
rect 28040 41692 28046 41744
rect 28626 41692 28632 41744
rect 28684 41732 28690 41744
rect 28813 41735 28871 41741
rect 28813 41732 28825 41735
rect 28684 41704 28825 41732
rect 28684 41692 28690 41704
rect 28813 41701 28825 41704
rect 28859 41732 28871 41735
rect 29086 41732 29092 41744
rect 28859 41704 29092 41732
rect 28859 41701 28871 41704
rect 28813 41695 28871 41701
rect 29086 41692 29092 41704
rect 29144 41692 29150 41744
rect 35989 41735 36047 41741
rect 35989 41701 36001 41735
rect 36035 41732 36047 41735
rect 37090 41732 37096 41744
rect 36035 41704 37096 41732
rect 36035 41701 36047 41704
rect 35989 41695 36047 41701
rect 37090 41692 37096 41704
rect 37148 41692 37154 41744
rect 29549 41667 29607 41673
rect 29549 41664 29561 41667
rect 29104 41636 29561 41664
rect 29104 41608 29132 41636
rect 29549 41633 29561 41636
rect 29595 41664 29607 41667
rect 29730 41664 29736 41676
rect 29595 41636 29736 41664
rect 29595 41633 29607 41636
rect 29549 41627 29607 41633
rect 29730 41624 29736 41636
rect 29788 41624 29794 41676
rect 34790 41664 34796 41676
rect 34751 41636 34796 41664
rect 34790 41624 34796 41636
rect 34848 41624 34854 41676
rect 35253 41667 35311 41673
rect 35253 41633 35265 41667
rect 35299 41664 35311 41667
rect 35802 41664 35808 41676
rect 35299 41636 35808 41664
rect 35299 41633 35311 41636
rect 35253 41627 35311 41633
rect 35802 41624 35808 41636
rect 35860 41624 35866 41676
rect 35894 41624 35900 41676
rect 35952 41664 35958 41676
rect 36722 41664 36728 41676
rect 35952 41636 36728 41664
rect 35952 41624 35958 41636
rect 36722 41624 36728 41636
rect 36780 41624 36786 41676
rect 36998 41624 37004 41676
rect 37056 41664 37062 41676
rect 37826 41664 37832 41676
rect 37056 41636 37832 41664
rect 37056 41624 37062 41636
rect 37826 41624 37832 41636
rect 37884 41624 37890 41676
rect 26252 41568 26372 41596
rect 9122 41460 9128 41472
rect 8496 41432 8892 41460
rect 9083 41432 9128 41460
rect 9122 41420 9128 41432
rect 9180 41420 9186 41472
rect 20162 41420 20168 41472
rect 20220 41420 20226 41472
rect 26344 41460 26372 41568
rect 26712 41568 27660 41596
rect 26712 41460 26740 41568
rect 29086 41556 29092 41608
rect 29144 41556 29150 41608
rect 34882 41556 34888 41608
rect 34940 41596 34946 41608
rect 35342 41596 35348 41608
rect 34940 41568 35348 41596
rect 34940 41556 34946 41568
rect 35342 41556 35348 41568
rect 35400 41556 35406 41608
rect 35526 41556 35532 41608
rect 35584 41556 35590 41608
rect 35820 41596 35848 41624
rect 36814 41596 36820 41608
rect 35820 41568 36820 41596
rect 36814 41556 36820 41568
rect 36872 41596 36878 41608
rect 36909 41599 36967 41605
rect 36909 41596 36921 41599
rect 36872 41568 36921 41596
rect 36872 41556 36878 41568
rect 36909 41565 36921 41568
rect 36955 41565 36967 41599
rect 36909 41559 36967 41565
rect 26789 41531 26847 41537
rect 26789 41497 26801 41531
rect 26835 41528 26847 41531
rect 27154 41528 27160 41540
rect 26835 41500 27160 41528
rect 26835 41497 26847 41500
rect 26789 41491 26847 41497
rect 27154 41488 27160 41500
rect 27212 41488 27218 41540
rect 27890 41488 27896 41540
rect 27948 41528 27954 41540
rect 29733 41531 29791 41537
rect 29733 41528 29745 41531
rect 27948 41500 29745 41528
rect 27948 41488 27954 41500
rect 29733 41497 29745 41500
rect 29779 41497 29791 41531
rect 35250 41528 35256 41540
rect 29733 41491 29791 41497
rect 34808 41500 35256 41528
rect 34808 41472 34836 41500
rect 35250 41488 35256 41500
rect 35308 41488 35314 41540
rect 35544 41528 35572 41556
rect 35802 41528 35808 41540
rect 35544 41500 35808 41528
rect 35802 41488 35808 41500
rect 35860 41488 35866 41540
rect 26344 41432 26740 41460
rect 27522 41420 27528 41472
rect 27580 41460 27586 41472
rect 28905 41463 28963 41469
rect 28905 41460 28917 41463
rect 27580 41432 28917 41460
rect 27580 41420 27586 41432
rect 28905 41429 28917 41432
rect 28951 41429 28963 41463
rect 28905 41423 28963 41429
rect 29178 41420 29184 41472
rect 29236 41460 29242 41472
rect 29914 41460 29920 41472
rect 29236 41432 29920 41460
rect 29236 41420 29242 41432
rect 29914 41420 29920 41432
rect 29972 41420 29978 41472
rect 30282 41420 30288 41472
rect 30340 41460 30346 41472
rect 32582 41460 32588 41472
rect 30340 41432 32588 41460
rect 30340 41420 30346 41432
rect 32582 41420 32588 41432
rect 32640 41420 32646 41472
rect 34790 41420 34796 41472
rect 34848 41420 34854 41472
rect 35526 41420 35532 41472
rect 35584 41460 35590 41472
rect 37366 41460 37372 41472
rect 35584 41432 37372 41460
rect 35584 41420 35590 41432
rect 37366 41420 37372 41432
rect 37424 41420 37430 41472
rect 1104 41370 38824 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 38824 41370
rect 1104 41296 38824 41318
rect 22830 41216 22836 41268
rect 22888 41256 22894 41268
rect 27065 41259 27123 41265
rect 22888 41228 27016 41256
rect 22888 41216 22894 41228
rect 2041 41191 2099 41197
rect 2041 41157 2053 41191
rect 2087 41188 2099 41191
rect 2130 41188 2136 41200
rect 2087 41160 2136 41188
rect 2087 41157 2099 41160
rect 2041 41151 2099 41157
rect 2130 41148 2136 41160
rect 2188 41148 2194 41200
rect 23106 41148 23112 41200
rect 23164 41188 23170 41200
rect 26988 41188 27016 41228
rect 27065 41225 27077 41259
rect 27111 41256 27123 41259
rect 27430 41256 27436 41268
rect 27111 41228 27436 41256
rect 27111 41225 27123 41228
rect 27065 41219 27123 41225
rect 27430 41216 27436 41228
rect 27488 41216 27494 41268
rect 34054 41216 34060 41268
rect 34112 41256 34118 41268
rect 34793 41259 34851 41265
rect 34793 41256 34805 41259
rect 34112 41228 34805 41256
rect 34112 41216 34118 41228
rect 34793 41225 34805 41228
rect 34839 41225 34851 41259
rect 34793 41219 34851 41225
rect 36173 41259 36231 41265
rect 36173 41225 36185 41259
rect 36219 41256 36231 41259
rect 38102 41256 38108 41268
rect 36219 41228 38108 41256
rect 36219 41225 36231 41228
rect 36173 41219 36231 41225
rect 38102 41216 38108 41228
rect 38160 41216 38166 41268
rect 36722 41188 36728 41200
rect 23164 41160 26740 41188
rect 26988 41160 36728 41188
rect 23164 41148 23170 41160
rect 6454 41080 6460 41132
rect 6512 41120 6518 41132
rect 6512 41092 8064 41120
rect 6512 41080 6518 41092
rect 1854 41052 1860 41064
rect 1815 41024 1860 41052
rect 1854 41012 1860 41024
rect 1912 41012 1918 41064
rect 7926 41052 7932 41064
rect 7887 41024 7932 41052
rect 7926 41012 7932 41024
rect 7984 41012 7990 41064
rect 8036 41061 8064 41092
rect 8202 41080 8208 41132
rect 8260 41120 8266 41132
rect 9493 41123 9551 41129
rect 9493 41120 9505 41123
rect 8260 41092 9505 41120
rect 8260 41080 8266 41092
rect 9493 41089 9505 41092
rect 9539 41089 9551 41123
rect 26712 41120 26740 41160
rect 36722 41148 36728 41160
rect 36780 41148 36786 41200
rect 37366 41148 37372 41200
rect 37424 41148 37430 41200
rect 9493 41083 9551 41089
rect 22066 41092 26648 41120
rect 26712 41092 36584 41120
rect 8021 41055 8079 41061
rect 8021 41021 8033 41055
rect 8067 41021 8079 41055
rect 8021 41015 8079 41021
rect 9582 41012 9588 41064
rect 9640 41052 9646 41064
rect 9677 41055 9735 41061
rect 9677 41052 9689 41055
rect 9640 41024 9689 41052
rect 9640 41012 9646 41024
rect 9677 41021 9689 41024
rect 9723 41021 9735 41055
rect 9677 41015 9735 41021
rect 10962 40944 10968 40996
rect 11020 40984 11026 40996
rect 22066 40984 22094 41092
rect 22370 41012 22376 41064
rect 22428 41052 22434 41064
rect 23106 41052 23112 41064
rect 22428 41024 23112 41052
rect 22428 41012 22434 41024
rect 23106 41012 23112 41024
rect 23164 41012 23170 41064
rect 26510 41052 26516 41064
rect 26471 41024 26516 41052
rect 26510 41012 26516 41024
rect 26568 41012 26574 41064
rect 26620 41052 26648 41092
rect 26886 41055 26944 41061
rect 26886 41052 26898 41055
rect 26620 41024 26898 41052
rect 26886 41021 26898 41024
rect 26932 41021 26944 41055
rect 34606 41052 34612 41064
rect 34567 41024 34612 41052
rect 26886 41015 26944 41021
rect 34606 41012 34612 41024
rect 34664 41012 34670 41064
rect 36173 41055 36231 41061
rect 36173 41021 36185 41055
rect 36219 41052 36231 41055
rect 36265 41055 36323 41061
rect 36265 41052 36277 41055
rect 36219 41024 36277 41052
rect 36219 41021 36231 41024
rect 36173 41015 36231 41021
rect 36265 41021 36277 41024
rect 36311 41021 36323 41055
rect 36265 41015 36323 41021
rect 36358 41055 36416 41061
rect 36358 41021 36370 41055
rect 36404 41021 36416 41055
rect 36556 41052 36584 41092
rect 36630 41080 36636 41132
rect 36688 41120 36694 41132
rect 37384 41120 37412 41148
rect 36688 41092 36860 41120
rect 37384 41092 37872 41120
rect 36688 41080 36694 41092
rect 36730 41055 36788 41061
rect 36730 41052 36742 41055
rect 36556 41024 36742 41052
rect 36358 41015 36416 41021
rect 36730 41021 36742 41024
rect 36776 41021 36788 41055
rect 36832 41052 36860 41092
rect 37366 41052 37372 41064
rect 36832 41024 37372 41052
rect 36730 41015 36788 41021
rect 11020 40956 22094 40984
rect 11020 40944 11026 40956
rect 26418 40944 26424 40996
rect 26476 40984 26482 40996
rect 26697 40987 26755 40993
rect 26697 40984 26709 40987
rect 26476 40956 26709 40984
rect 26476 40944 26482 40956
rect 26697 40953 26709 40956
rect 26743 40953 26755 40987
rect 26697 40947 26755 40953
rect 26786 40944 26792 40996
rect 26844 40984 26850 40996
rect 28721 40987 28779 40993
rect 26844 40956 26889 40984
rect 26844 40944 26850 40956
rect 28721 40953 28733 40987
rect 28767 40984 28779 40987
rect 29086 40984 29092 40996
rect 28767 40956 29092 40984
rect 28767 40953 28779 40956
rect 28721 40947 28779 40953
rect 29086 40944 29092 40956
rect 29144 40944 29150 40996
rect 30742 40944 30748 40996
rect 30800 40984 30806 40996
rect 31570 40984 31576 40996
rect 30800 40956 31576 40984
rect 30800 40944 30806 40956
rect 31570 40944 31576 40956
rect 31628 40944 31634 40996
rect 34146 40944 34152 40996
rect 34204 40984 34210 40996
rect 34790 40984 34796 40996
rect 34204 40956 34796 40984
rect 34204 40944 34210 40956
rect 34790 40944 34796 40956
rect 34848 40944 34854 40996
rect 35342 40944 35348 40996
rect 35400 40984 35406 40996
rect 36372 40984 36400 41015
rect 37366 41012 37372 41024
rect 37424 41012 37430 41064
rect 37550 41052 37556 41064
rect 37511 41024 37556 41052
rect 37550 41012 37556 41024
rect 37608 41012 37614 41064
rect 37844 41061 37872 41092
rect 37829 41055 37887 41061
rect 37829 41021 37841 41055
rect 37875 41021 37887 41055
rect 37829 41015 37887 41021
rect 37921 41055 37979 41061
rect 37921 41021 37933 41055
rect 37967 41052 37979 41055
rect 38838 41052 38844 41064
rect 37967 41024 38844 41052
rect 37967 41021 37979 41024
rect 37921 41015 37979 41021
rect 38838 41012 38844 41024
rect 38896 41012 38902 41064
rect 36538 40984 36544 40996
rect 35400 40956 36400 40984
rect 36499 40956 36544 40984
rect 35400 40944 35406 40956
rect 36538 40944 36544 40956
rect 36596 40944 36602 40996
rect 36630 40944 36636 40996
rect 36688 40984 36694 40996
rect 36688 40956 36733 40984
rect 36688 40944 36694 40956
rect 37458 40944 37464 40996
rect 37516 40984 37522 40996
rect 37737 40987 37795 40993
rect 37737 40984 37749 40987
rect 37516 40956 37749 40984
rect 37516 40944 37522 40956
rect 37737 40953 37749 40956
rect 37783 40953 37795 40987
rect 37737 40947 37795 40953
rect 7466 40876 7472 40928
rect 7524 40916 7530 40928
rect 8205 40919 8263 40925
rect 8205 40916 8217 40919
rect 7524 40888 8217 40916
rect 7524 40876 7530 40888
rect 8205 40885 8217 40888
rect 8251 40885 8263 40919
rect 8205 40879 8263 40885
rect 9861 40919 9919 40925
rect 9861 40885 9873 40919
rect 9907 40916 9919 40919
rect 9950 40916 9956 40928
rect 9907 40888 9956 40916
rect 9907 40885 9919 40888
rect 9861 40879 9919 40885
rect 9950 40876 9956 40888
rect 10008 40876 10014 40928
rect 27890 40876 27896 40928
rect 27948 40916 27954 40928
rect 28813 40919 28871 40925
rect 28813 40916 28825 40919
rect 27948 40888 28825 40916
rect 27948 40876 27954 40888
rect 28813 40885 28825 40888
rect 28859 40885 28871 40919
rect 28813 40879 28871 40885
rect 34330 40876 34336 40928
rect 34388 40916 34394 40928
rect 35434 40916 35440 40928
rect 34388 40888 35440 40916
rect 34388 40876 34394 40888
rect 35434 40876 35440 40888
rect 35492 40876 35498 40928
rect 36906 40916 36912 40928
rect 36867 40888 36912 40916
rect 36906 40876 36912 40888
rect 36964 40876 36970 40928
rect 37090 40876 37096 40928
rect 37148 40916 37154 40928
rect 38105 40919 38163 40925
rect 38105 40916 38117 40919
rect 37148 40888 38117 40916
rect 37148 40876 37154 40888
rect 38105 40885 38117 40888
rect 38151 40885 38163 40919
rect 38105 40879 38163 40885
rect 1104 40826 38824 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 38824 40826
rect 1104 40752 38824 40774
rect 1578 40672 1584 40724
rect 1636 40712 1642 40724
rect 24854 40712 24860 40724
rect 1636 40684 8892 40712
rect 24815 40684 24860 40712
rect 1636 40672 1642 40684
rect 4890 40604 4896 40656
rect 4948 40644 4954 40656
rect 4948 40616 6914 40644
rect 4948 40604 4954 40616
rect 6886 40576 6914 40616
rect 8021 40579 8079 40585
rect 8021 40576 8033 40579
rect 6886 40548 8033 40576
rect 8021 40545 8033 40548
rect 8067 40545 8079 40579
rect 8021 40539 8079 40545
rect 8202 40536 8208 40588
rect 8260 40576 8266 40588
rect 8864 40585 8892 40684
rect 24854 40672 24860 40684
rect 24912 40672 24918 40724
rect 26510 40672 26516 40724
rect 26568 40712 26574 40724
rect 34054 40712 34060 40724
rect 26568 40684 34060 40712
rect 26568 40672 26574 40684
rect 34054 40672 34060 40684
rect 34112 40672 34118 40724
rect 35621 40715 35679 40721
rect 35621 40681 35633 40715
rect 35667 40712 35679 40715
rect 36998 40712 37004 40724
rect 35667 40684 36216 40712
rect 35667 40681 35679 40684
rect 35621 40675 35679 40681
rect 24213 40647 24271 40653
rect 24213 40613 24225 40647
rect 24259 40644 24271 40647
rect 24302 40644 24308 40656
rect 24259 40616 24308 40644
rect 24259 40613 24271 40616
rect 24213 40607 24271 40613
rect 24302 40604 24308 40616
rect 24360 40604 24366 40656
rect 28994 40653 29000 40656
rect 28988 40644 29000 40653
rect 28955 40616 29000 40644
rect 28988 40607 29000 40616
rect 28994 40604 29000 40607
rect 29052 40604 29058 40656
rect 8665 40579 8723 40585
rect 8665 40576 8677 40579
rect 8260 40548 8677 40576
rect 8260 40536 8266 40548
rect 8665 40545 8677 40548
rect 8711 40545 8723 40579
rect 8665 40539 8723 40545
rect 8849 40579 8907 40585
rect 8849 40545 8861 40579
rect 8895 40545 8907 40579
rect 8849 40539 8907 40545
rect 22557 40579 22615 40585
rect 22557 40545 22569 40579
rect 22603 40576 22615 40579
rect 24670 40576 24676 40588
rect 22603 40548 23060 40576
rect 24583 40548 24676 40576
rect 22603 40545 22615 40548
rect 22557 40539 22615 40545
rect 7837 40511 7895 40517
rect 7837 40477 7849 40511
rect 7883 40508 7895 40511
rect 7926 40508 7932 40520
rect 7883 40480 7932 40508
rect 7883 40477 7895 40480
rect 7837 40471 7895 40477
rect 7926 40468 7932 40480
rect 7984 40468 7990 40520
rect 8220 40440 8248 40536
rect 23032 40520 23060 40548
rect 24670 40536 24676 40548
rect 24728 40536 24734 40588
rect 26510 40536 26516 40588
rect 26568 40576 26574 40588
rect 28810 40576 28816 40588
rect 26568 40548 28816 40576
rect 26568 40536 26574 40548
rect 28810 40536 28816 40548
rect 28868 40536 28874 40588
rect 29270 40536 29276 40588
rect 29328 40576 29334 40588
rect 30006 40576 30012 40588
rect 29328 40548 30012 40576
rect 29328 40536 29334 40548
rect 30006 40536 30012 40548
rect 30064 40536 30070 40588
rect 35158 40576 35164 40588
rect 35119 40548 35164 40576
rect 35158 40536 35164 40548
rect 35216 40536 35222 40588
rect 35802 40576 35808 40588
rect 35763 40548 35808 40576
rect 35802 40536 35808 40548
rect 35860 40536 35866 40588
rect 22830 40508 22836 40520
rect 22791 40480 22836 40508
rect 22830 40468 22836 40480
rect 22888 40468 22894 40520
rect 23014 40468 23020 40520
rect 23072 40468 23078 40520
rect 7944 40412 8248 40440
rect 7944 40384 7972 40412
rect 8570 40400 8576 40452
rect 8628 40440 8634 40452
rect 21542 40440 21548 40452
rect 8628 40412 21548 40440
rect 8628 40400 8634 40412
rect 21542 40400 21548 40412
rect 21600 40400 21606 40452
rect 7926 40332 7932 40384
rect 7984 40332 7990 40384
rect 8110 40332 8116 40384
rect 8168 40372 8174 40384
rect 8205 40375 8263 40381
rect 8205 40372 8217 40375
rect 8168 40344 8217 40372
rect 8168 40332 8174 40344
rect 8205 40341 8217 40344
rect 8251 40341 8263 40375
rect 8205 40335 8263 40341
rect 9033 40375 9091 40381
rect 9033 40341 9045 40375
rect 9079 40372 9091 40375
rect 13538 40372 13544 40384
rect 9079 40344 13544 40372
rect 9079 40341 9091 40344
rect 9033 40335 9091 40341
rect 13538 40332 13544 40344
rect 13596 40332 13602 40384
rect 21358 40332 21364 40384
rect 21416 40372 21422 40384
rect 24688 40372 24716 40536
rect 27430 40468 27436 40520
rect 27488 40508 27494 40520
rect 28721 40511 28779 40517
rect 28721 40508 28733 40511
rect 27488 40480 28733 40508
rect 27488 40468 27494 40480
rect 28721 40477 28733 40480
rect 28767 40477 28779 40511
rect 28721 40471 28779 40477
rect 34882 40468 34888 40520
rect 34940 40508 34946 40520
rect 35434 40508 35440 40520
rect 34940 40480 35440 40508
rect 34940 40468 34946 40480
rect 35434 40468 35440 40480
rect 35492 40468 35498 40520
rect 36188 40508 36216 40684
rect 36280 40684 37004 40712
rect 36280 40585 36308 40684
rect 36998 40672 37004 40684
rect 37056 40672 37062 40724
rect 36538 40644 36544 40656
rect 36499 40616 36544 40644
rect 36538 40604 36544 40616
rect 36596 40604 36602 40656
rect 36265 40579 36323 40585
rect 36265 40545 36277 40579
rect 36311 40545 36323 40579
rect 36265 40539 36323 40545
rect 36354 40536 36360 40588
rect 36412 40576 36418 40588
rect 36630 40576 36636 40588
rect 36412 40548 36457 40576
rect 36591 40548 36636 40576
rect 36412 40536 36418 40548
rect 36630 40536 36636 40548
rect 36688 40536 36694 40588
rect 36722 40536 36728 40588
rect 36780 40585 36786 40588
rect 36780 40576 36788 40585
rect 36780 40548 36825 40576
rect 36780 40539 36788 40548
rect 36780 40536 36786 40539
rect 38562 40508 38568 40520
rect 36188 40480 38568 40508
rect 38562 40468 38568 40480
rect 38620 40468 38626 40520
rect 29730 40400 29736 40452
rect 29788 40440 29794 40452
rect 33962 40440 33968 40452
rect 29788 40412 33968 40440
rect 29788 40400 29794 40412
rect 33962 40400 33968 40412
rect 34020 40400 34026 40452
rect 34977 40443 35035 40449
rect 34977 40409 34989 40443
rect 35023 40440 35035 40443
rect 36078 40440 36084 40452
rect 35023 40412 36084 40440
rect 35023 40409 35035 40412
rect 34977 40403 35035 40409
rect 36078 40400 36084 40412
rect 36136 40400 36142 40452
rect 21416 40344 24716 40372
rect 30101 40375 30159 40381
rect 21416 40332 21422 40344
rect 30101 40341 30113 40375
rect 30147 40372 30159 40375
rect 30650 40372 30656 40384
rect 30147 40344 30656 40372
rect 30147 40341 30159 40344
rect 30101 40335 30159 40341
rect 30650 40332 30656 40344
rect 30708 40332 30714 40384
rect 32950 40332 32956 40384
rect 33008 40372 33014 40384
rect 36909 40375 36967 40381
rect 36909 40372 36921 40375
rect 33008 40344 36921 40372
rect 33008 40332 33014 40344
rect 36909 40341 36921 40344
rect 36955 40341 36967 40375
rect 36909 40335 36967 40341
rect 1104 40282 38824 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 38824 40282
rect 1104 40208 38824 40230
rect 20254 40128 20260 40180
rect 20312 40168 20318 40180
rect 37550 40168 37556 40180
rect 20312 40140 37556 40168
rect 20312 40128 20318 40140
rect 37550 40128 37556 40140
rect 37608 40128 37614 40180
rect 37826 40128 37832 40180
rect 37884 40168 37890 40180
rect 38562 40168 38568 40180
rect 37884 40140 38568 40168
rect 37884 40128 37890 40140
rect 38562 40128 38568 40140
rect 38620 40128 38626 40180
rect 26786 40060 26792 40112
rect 26844 40100 26850 40112
rect 27798 40100 27804 40112
rect 26844 40072 27804 40100
rect 26844 40060 26850 40072
rect 27798 40060 27804 40072
rect 27856 40060 27862 40112
rect 29270 40060 29276 40112
rect 29328 40100 29334 40112
rect 32214 40100 32220 40112
rect 29328 40072 32220 40100
rect 29328 40060 29334 40072
rect 32214 40060 32220 40072
rect 32272 40060 32278 40112
rect 36173 40103 36231 40109
rect 36173 40069 36185 40103
rect 36219 40100 36231 40103
rect 36219 40072 36768 40100
rect 36219 40069 36231 40072
rect 36173 40063 36231 40069
rect 2038 40032 2044 40044
rect 1999 40004 2044 40032
rect 2038 39992 2044 40004
rect 2096 39992 2102 40044
rect 8018 40032 8024 40044
rect 7979 40004 8024 40032
rect 8018 39992 8024 40004
rect 8076 39992 8082 40044
rect 9858 39992 9864 40044
rect 9916 40032 9922 40044
rect 11698 40032 11704 40044
rect 9916 40004 11704 40032
rect 9916 39992 9922 40004
rect 11698 39992 11704 40004
rect 11756 39992 11762 40044
rect 17310 39992 17316 40044
rect 17368 40032 17374 40044
rect 22462 40032 22468 40044
rect 17368 40004 22468 40032
rect 17368 39992 17374 40004
rect 22462 39992 22468 40004
rect 22520 39992 22526 40044
rect 32674 40032 32680 40044
rect 31726 40004 32680 40032
rect 1854 39964 1860 39976
rect 1815 39936 1860 39964
rect 1854 39924 1860 39936
rect 1912 39924 1918 39976
rect 7926 39924 7932 39976
rect 7984 39964 7990 39976
rect 8205 39967 8263 39973
rect 8205 39964 8217 39967
rect 7984 39936 8217 39964
rect 7984 39924 7990 39936
rect 8205 39933 8217 39936
rect 8251 39933 8263 39967
rect 8205 39927 8263 39933
rect 27430 39924 27436 39976
rect 27488 39964 27494 39976
rect 27798 39964 27804 39976
rect 27488 39936 27804 39964
rect 27488 39924 27494 39936
rect 27798 39924 27804 39936
rect 27856 39964 27862 39976
rect 28077 39967 28135 39973
rect 28077 39964 28089 39967
rect 27856 39936 28089 39964
rect 27856 39924 27862 39936
rect 28077 39933 28089 39936
rect 28123 39933 28135 39967
rect 28077 39927 28135 39933
rect 28344 39967 28402 39973
rect 28344 39933 28356 39967
rect 28390 39964 28402 39967
rect 29546 39964 29552 39976
rect 28390 39936 29552 39964
rect 28390 39933 28402 39936
rect 28344 39927 28402 39933
rect 29546 39924 29552 39936
rect 29604 39924 29610 39976
rect 28810 39856 28816 39908
rect 28868 39896 28874 39908
rect 31726 39896 31754 40004
rect 32674 39992 32680 40004
rect 32732 39992 32738 40044
rect 35710 39992 35716 40044
rect 35768 40032 35774 40044
rect 36740 40032 36768 40072
rect 37274 40032 37280 40044
rect 35768 40004 36676 40032
rect 36740 40004 37280 40032
rect 35768 39992 35774 40004
rect 34606 39964 34612 39976
rect 34567 39936 34612 39964
rect 34606 39924 34612 39936
rect 34664 39924 34670 39976
rect 36078 39964 36084 39976
rect 34716 39936 36084 39964
rect 28868 39868 31754 39896
rect 28868 39856 28874 39868
rect 32214 39856 32220 39908
rect 32272 39896 32278 39908
rect 34716 39896 34744 39936
rect 36078 39924 36084 39936
rect 36136 39924 36142 39976
rect 36173 39967 36231 39973
rect 36173 39933 36185 39967
rect 36219 39964 36231 39967
rect 36265 39967 36323 39973
rect 36265 39964 36277 39967
rect 36219 39936 36277 39964
rect 36219 39933 36231 39936
rect 36173 39927 36231 39933
rect 36265 39933 36277 39936
rect 36311 39933 36323 39967
rect 36265 39927 36323 39933
rect 36358 39967 36416 39973
rect 36358 39933 36370 39967
rect 36404 39933 36416 39967
rect 36538 39964 36544 39976
rect 36499 39936 36544 39964
rect 36358 39927 36416 39933
rect 32272 39868 34744 39896
rect 32272 39856 32278 39868
rect 35802 39856 35808 39908
rect 35860 39896 35866 39908
rect 36372 39896 36400 39927
rect 36538 39924 36544 39936
rect 36596 39924 36602 39976
rect 36648 39964 36676 40004
rect 37274 39992 37280 40004
rect 37332 39992 37338 40044
rect 38286 40032 38292 40044
rect 37752 40004 38292 40032
rect 37752 39976 37780 40004
rect 38286 39992 38292 40004
rect 38344 39992 38350 40044
rect 36730 39967 36788 39973
rect 36730 39964 36742 39967
rect 36648 39936 36742 39964
rect 36730 39933 36742 39936
rect 36776 39933 36788 39967
rect 36730 39927 36788 39933
rect 37553 39967 37611 39973
rect 37553 39933 37565 39967
rect 37599 39933 37611 39967
rect 37734 39964 37740 39976
rect 37647 39936 37740 39964
rect 37553 39927 37611 39933
rect 36630 39896 36636 39908
rect 35860 39868 36400 39896
rect 36591 39868 36636 39896
rect 35860 39856 35866 39868
rect 36630 39856 36636 39868
rect 36688 39856 36694 39908
rect 37568 39896 37596 39927
rect 37734 39924 37740 39936
rect 37792 39924 37798 39976
rect 37921 39967 37979 39973
rect 37921 39933 37933 39967
rect 37967 39964 37979 39967
rect 38102 39964 38108 39976
rect 37967 39936 38108 39964
rect 37967 39933 37979 39936
rect 37921 39927 37979 39933
rect 38102 39924 38108 39936
rect 38160 39924 38166 39976
rect 36740 39868 37596 39896
rect 37829 39899 37887 39905
rect 8386 39828 8392 39840
rect 8347 39800 8392 39828
rect 8386 39788 8392 39800
rect 8444 39788 8450 39840
rect 29457 39831 29515 39837
rect 29457 39797 29469 39831
rect 29503 39828 29515 39831
rect 29546 39828 29552 39840
rect 29503 39800 29552 39828
rect 29503 39797 29515 39800
rect 29457 39791 29515 39797
rect 29546 39788 29552 39800
rect 29604 39788 29610 39840
rect 31294 39788 31300 39840
rect 31352 39828 31358 39840
rect 34793 39831 34851 39837
rect 34793 39828 34805 39831
rect 31352 39800 34805 39828
rect 31352 39788 31358 39800
rect 34793 39797 34805 39800
rect 34839 39797 34851 39831
rect 34793 39791 34851 39797
rect 34882 39788 34888 39840
rect 34940 39828 34946 39840
rect 36740 39828 36768 39868
rect 37829 39865 37841 39899
rect 37875 39896 37887 39899
rect 38010 39896 38016 39908
rect 37875 39868 38016 39896
rect 37875 39865 37887 39868
rect 37829 39859 37887 39865
rect 38010 39856 38016 39868
rect 38068 39856 38074 39908
rect 36906 39828 36912 39840
rect 34940 39800 36768 39828
rect 36867 39800 36912 39828
rect 34940 39788 34946 39800
rect 36906 39788 36912 39800
rect 36964 39788 36970 39840
rect 37550 39788 37556 39840
rect 37608 39828 37614 39840
rect 38105 39831 38163 39837
rect 38105 39828 38117 39831
rect 37608 39800 38117 39828
rect 37608 39788 37614 39800
rect 38105 39797 38117 39800
rect 38151 39797 38163 39831
rect 38105 39791 38163 39797
rect 1104 39738 38824 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 38824 39738
rect 1104 39664 38824 39686
rect 1949 39627 2007 39633
rect 1949 39593 1961 39627
rect 1995 39624 2007 39627
rect 2682 39624 2688 39636
rect 1995 39596 2688 39624
rect 1995 39593 2007 39596
rect 1949 39587 2007 39593
rect 2682 39584 2688 39596
rect 2740 39584 2746 39636
rect 18966 39584 18972 39636
rect 19024 39624 19030 39636
rect 34882 39624 34888 39636
rect 19024 39596 34888 39624
rect 19024 39584 19030 39596
rect 34882 39584 34888 39596
rect 34940 39584 34946 39636
rect 35069 39627 35127 39633
rect 35069 39593 35081 39627
rect 35115 39624 35127 39627
rect 35526 39624 35532 39636
rect 35115 39596 35532 39624
rect 35115 39593 35127 39596
rect 35069 39587 35127 39593
rect 35526 39584 35532 39596
rect 35584 39584 35590 39636
rect 36722 39624 36728 39636
rect 36428 39596 36728 39624
rect 2130 39516 2136 39568
rect 2188 39556 2194 39568
rect 10962 39556 10968 39568
rect 2188 39528 10968 39556
rect 2188 39516 2194 39528
rect 10962 39516 10968 39528
rect 11020 39516 11026 39568
rect 28436 39559 28494 39565
rect 28436 39525 28448 39559
rect 28482 39556 28494 39559
rect 28902 39556 28908 39568
rect 28482 39528 28908 39556
rect 28482 39525 28494 39528
rect 28436 39519 28494 39525
rect 28902 39516 28908 39528
rect 28960 39516 28966 39568
rect 29546 39516 29552 39568
rect 29604 39556 29610 39568
rect 30190 39556 30196 39568
rect 29604 39528 30196 39556
rect 29604 39516 29610 39528
rect 30190 39516 30196 39528
rect 30248 39516 30254 39568
rect 30374 39565 30380 39568
rect 30368 39556 30380 39565
rect 30335 39528 30380 39556
rect 30368 39519 30380 39528
rect 30374 39516 30380 39519
rect 30432 39516 30438 39568
rect 31294 39516 31300 39568
rect 31352 39556 31358 39568
rect 32306 39556 32312 39568
rect 31352 39528 32312 39556
rect 31352 39516 31358 39528
rect 32306 39516 32312 39528
rect 32364 39516 32370 39568
rect 32674 39516 32680 39568
rect 32732 39556 32738 39568
rect 36078 39556 36084 39568
rect 32732 39528 36084 39556
rect 32732 39516 32738 39528
rect 36078 39516 36084 39528
rect 36136 39516 36142 39568
rect 1854 39488 1860 39500
rect 1815 39460 1860 39488
rect 1854 39448 1860 39460
rect 1912 39448 1918 39500
rect 8202 39448 8208 39500
rect 8260 39488 8266 39500
rect 17494 39488 17500 39500
rect 8260 39460 17500 39488
rect 8260 39448 8266 39460
rect 17494 39448 17500 39460
rect 17552 39448 17558 39500
rect 30101 39491 30159 39497
rect 30101 39488 30113 39491
rect 28184 39460 30113 39488
rect 2038 39380 2044 39432
rect 2096 39420 2102 39432
rect 9490 39420 9496 39432
rect 2096 39392 9496 39420
rect 2096 39380 2102 39392
rect 9490 39380 9496 39392
rect 9548 39380 9554 39432
rect 16850 39420 16856 39432
rect 9600 39392 16856 39420
rect 9214 39312 9220 39364
rect 9272 39352 9278 39364
rect 9600 39352 9628 39392
rect 16850 39380 16856 39392
rect 16908 39380 16914 39432
rect 27798 39380 27804 39432
rect 27856 39420 27862 39432
rect 28184 39429 28212 39460
rect 30101 39457 30113 39460
rect 30147 39457 30159 39491
rect 30101 39451 30159 39457
rect 34425 39491 34483 39497
rect 34425 39457 34437 39491
rect 34471 39488 34483 39491
rect 34514 39488 34520 39500
rect 34471 39460 34520 39488
rect 34471 39457 34483 39460
rect 34425 39451 34483 39457
rect 34514 39448 34520 39460
rect 34572 39448 34578 39500
rect 34885 39491 34943 39497
rect 34885 39457 34897 39491
rect 34931 39488 34943 39491
rect 35526 39488 35532 39500
rect 34931 39460 35532 39488
rect 34931 39457 34943 39460
rect 34885 39451 34943 39457
rect 35526 39448 35532 39460
rect 35584 39448 35590 39500
rect 35621 39491 35679 39497
rect 35621 39457 35633 39491
rect 35667 39488 35679 39491
rect 35894 39488 35900 39500
rect 35667 39460 35900 39488
rect 35667 39457 35679 39460
rect 35621 39451 35679 39457
rect 35894 39448 35900 39460
rect 35952 39448 35958 39500
rect 36262 39488 36268 39500
rect 36223 39460 36268 39488
rect 36262 39448 36268 39460
rect 36320 39448 36326 39500
rect 36428 39497 36456 39596
rect 36722 39584 36728 39596
rect 36780 39584 36786 39636
rect 36538 39556 36544 39568
rect 36499 39528 36544 39556
rect 36538 39516 36544 39528
rect 36596 39516 36602 39568
rect 36413 39491 36471 39497
rect 36413 39457 36425 39491
rect 36459 39457 36471 39491
rect 36630 39488 36636 39500
rect 36591 39460 36636 39488
rect 36413 39451 36471 39457
rect 36630 39448 36636 39460
rect 36688 39448 36694 39500
rect 36730 39491 36788 39497
rect 36730 39457 36742 39491
rect 36776 39457 36788 39491
rect 36730 39451 36788 39457
rect 28169 39423 28227 39429
rect 28169 39420 28181 39423
rect 27856 39392 28181 39420
rect 27856 39380 27862 39392
rect 28169 39389 28181 39392
rect 28215 39389 28227 39423
rect 28169 39383 28227 39389
rect 35250 39380 35256 39432
rect 35308 39420 35314 39432
rect 36745 39420 36773 39451
rect 35308 39392 36773 39420
rect 35308 39380 35314 39392
rect 9272 39324 9628 39352
rect 9272 39312 9278 39324
rect 12342 39312 12348 39364
rect 12400 39352 12406 39364
rect 22554 39352 22560 39364
rect 12400 39324 22560 39352
rect 12400 39312 12406 39324
rect 22554 39312 22560 39324
rect 22612 39312 22618 39364
rect 23382 39312 23388 39364
rect 23440 39352 23446 39364
rect 24026 39352 24032 39364
rect 23440 39324 24032 39352
rect 23440 39312 23446 39324
rect 24026 39312 24032 39324
rect 24084 39312 24090 39364
rect 31478 39352 31484 39364
rect 31439 39324 31484 39352
rect 31478 39312 31484 39324
rect 31536 39312 31542 39364
rect 34241 39355 34299 39361
rect 34241 39321 34253 39355
rect 34287 39352 34299 39355
rect 35986 39352 35992 39364
rect 34287 39324 35992 39352
rect 34287 39321 34299 39324
rect 34241 39315 34299 39321
rect 35986 39312 35992 39324
rect 36044 39312 36050 39364
rect 36078 39312 36084 39364
rect 36136 39352 36142 39364
rect 36909 39355 36967 39361
rect 36909 39352 36921 39355
rect 36136 39324 36921 39352
rect 36136 39312 36142 39324
rect 36909 39321 36921 39324
rect 36955 39321 36967 39355
rect 36909 39315 36967 39321
rect 23290 39244 23296 39296
rect 23348 39284 23354 39296
rect 28902 39284 28908 39296
rect 23348 39256 28908 39284
rect 23348 39244 23354 39256
rect 28902 39244 28908 39256
rect 28960 39244 28966 39296
rect 29546 39284 29552 39296
rect 29507 39256 29552 39284
rect 29546 39244 29552 39256
rect 29604 39244 29610 39296
rect 35713 39287 35771 39293
rect 35713 39253 35725 39287
rect 35759 39284 35771 39287
rect 36262 39284 36268 39296
rect 35759 39256 36268 39284
rect 35759 39253 35771 39256
rect 35713 39247 35771 39253
rect 36262 39244 36268 39256
rect 36320 39244 36326 39296
rect 1104 39194 38824 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 38824 39194
rect 1104 39120 38824 39142
rect 22830 39040 22836 39092
rect 22888 39080 22894 39092
rect 23569 39083 23627 39089
rect 23569 39080 23581 39083
rect 22888 39052 23581 39080
rect 22888 39040 22894 39052
rect 23569 39049 23581 39052
rect 23615 39049 23627 39083
rect 23569 39043 23627 39049
rect 25406 39040 25412 39092
rect 25464 39080 25470 39092
rect 29457 39083 29515 39089
rect 29457 39080 29469 39083
rect 25464 39052 29469 39080
rect 25464 39040 25470 39052
rect 29457 39049 29469 39052
rect 29503 39049 29515 39083
rect 29457 39043 29515 39049
rect 30558 39040 30564 39092
rect 30616 39080 30622 39092
rect 31478 39080 31484 39092
rect 30616 39052 31484 39080
rect 30616 39040 30622 39052
rect 31478 39040 31484 39052
rect 31536 39040 31542 39092
rect 32858 39040 32864 39092
rect 32916 39080 32922 39092
rect 34793 39083 34851 39089
rect 34793 39080 34805 39083
rect 32916 39052 34805 39080
rect 32916 39040 32922 39052
rect 34793 39049 34805 39052
rect 34839 39049 34851 39083
rect 34793 39043 34851 39049
rect 35526 39040 35532 39092
rect 35584 39080 35590 39092
rect 35986 39080 35992 39092
rect 35584 39052 35992 39080
rect 35584 39040 35590 39052
rect 35986 39040 35992 39052
rect 36044 39040 36050 39092
rect 36173 39083 36231 39089
rect 36173 39049 36185 39083
rect 36219 39080 36231 39083
rect 37090 39080 37096 39092
rect 36219 39052 36860 39080
rect 36219 39049 36231 39052
rect 36173 39043 36231 39049
rect 22281 39015 22339 39021
rect 22281 38981 22293 39015
rect 22327 39012 22339 39015
rect 28074 39012 28080 39024
rect 22327 38984 28080 39012
rect 22327 38981 22339 38984
rect 22281 38975 22339 38981
rect 28074 38972 28080 38984
rect 28132 38972 28138 39024
rect 35250 38972 35256 39024
rect 35308 39012 35314 39024
rect 36078 39012 36084 39024
rect 35308 38984 36084 39012
rect 35308 38972 35314 38984
rect 36078 38972 36084 38984
rect 36136 38972 36142 39024
rect 36465 38984 36773 39012
rect 6270 38904 6276 38956
rect 6328 38944 6334 38956
rect 23474 38944 23480 38956
rect 6328 38916 21956 38944
rect 6328 38904 6334 38916
rect 17678 38836 17684 38888
rect 17736 38876 17742 38888
rect 21818 38885 21824 38888
rect 21637 38879 21695 38885
rect 21637 38876 21649 38879
rect 17736 38848 21649 38876
rect 17736 38836 17742 38848
rect 21637 38845 21649 38848
rect 21683 38845 21695 38879
rect 21637 38839 21695 38845
rect 21785 38879 21824 38885
rect 21785 38845 21797 38879
rect 21785 38839 21824 38845
rect 21818 38836 21824 38839
rect 21876 38836 21882 38888
rect 21928 38876 21956 38916
rect 23124 38916 23480 38944
rect 22102 38879 22160 38885
rect 22102 38876 22114 38879
rect 21928 38848 22114 38876
rect 22102 38845 22114 38848
rect 22148 38845 22160 38879
rect 23014 38876 23020 38888
rect 22975 38848 23020 38876
rect 22102 38839 22160 38845
rect 23014 38836 23020 38848
rect 23072 38836 23078 38888
rect 21910 38808 21916 38820
rect 21871 38780 21916 38808
rect 21910 38768 21916 38780
rect 21968 38768 21974 38820
rect 22005 38811 22063 38817
rect 22005 38777 22017 38811
rect 22051 38808 22063 38811
rect 23124 38808 23152 38916
rect 23474 38904 23480 38916
rect 23532 38904 23538 38956
rect 24026 38904 24032 38956
rect 24084 38944 24090 38956
rect 36465 38944 36493 38984
rect 24084 38916 36493 38944
rect 24084 38904 24090 38916
rect 36538 38904 36544 38956
rect 36596 38904 36602 38956
rect 23385 38879 23443 38885
rect 23385 38845 23397 38879
rect 23431 38876 23443 38879
rect 24302 38876 24308 38888
rect 23431 38848 24308 38876
rect 23431 38845 23443 38848
rect 23385 38839 23443 38845
rect 24302 38836 24308 38848
rect 24360 38836 24366 38888
rect 25222 38876 25228 38888
rect 25183 38848 25228 38876
rect 25222 38836 25228 38848
rect 25280 38836 25286 38888
rect 25409 38879 25467 38885
rect 25409 38845 25421 38879
rect 25455 38876 25467 38879
rect 25498 38876 25504 38888
rect 25455 38848 25504 38876
rect 25455 38845 25467 38848
rect 25409 38839 25467 38845
rect 22051 38780 23152 38808
rect 23201 38811 23259 38817
rect 22051 38777 22063 38780
rect 22005 38771 22063 38777
rect 23201 38777 23213 38811
rect 23247 38777 23259 38811
rect 23201 38771 23259 38777
rect 23293 38811 23351 38817
rect 23293 38777 23305 38811
rect 23339 38808 23351 38811
rect 24394 38808 24400 38820
rect 23339 38780 24400 38808
rect 23339 38777 23351 38780
rect 23293 38771 23351 38777
rect 23216 38740 23244 38771
rect 24394 38768 24400 38780
rect 24452 38808 24458 38820
rect 25424 38808 25452 38839
rect 25498 38836 25504 38848
rect 25556 38836 25562 38888
rect 28626 38876 28632 38888
rect 28587 38848 28632 38876
rect 28626 38836 28632 38848
rect 28684 38836 28690 38888
rect 29086 38836 29092 38888
rect 29144 38876 29150 38888
rect 29365 38879 29423 38885
rect 29365 38876 29377 38879
rect 29144 38848 29377 38876
rect 29144 38836 29150 38848
rect 29365 38845 29377 38848
rect 29411 38845 29423 38879
rect 29365 38839 29423 38845
rect 34609 38879 34667 38885
rect 34609 38845 34621 38879
rect 34655 38876 34667 38879
rect 34790 38876 34796 38888
rect 34655 38848 34796 38876
rect 34655 38845 34667 38848
rect 34609 38839 34667 38845
rect 34790 38836 34796 38848
rect 34848 38836 34854 38888
rect 36173 38879 36231 38885
rect 36173 38845 36185 38879
rect 36219 38876 36231 38879
rect 36265 38879 36323 38885
rect 36265 38876 36277 38879
rect 36219 38848 36277 38876
rect 36219 38845 36231 38848
rect 36173 38839 36231 38845
rect 36265 38845 36277 38848
rect 36311 38845 36323 38879
rect 36265 38839 36323 38845
rect 36413 38879 36471 38885
rect 36413 38845 36425 38879
rect 36459 38876 36471 38879
rect 36556 38876 36584 38904
rect 36745 38885 36773 38984
rect 36832 38944 36860 39052
rect 37016 39052 37096 39080
rect 37016 38944 37044 39052
rect 37090 39040 37096 39052
rect 37148 39040 37154 39092
rect 38102 39080 38108 39092
rect 37752 39052 38108 39080
rect 36832 38916 37044 38944
rect 37274 38904 37280 38956
rect 37332 38944 37338 38956
rect 37332 38916 37596 38944
rect 37332 38904 37338 38916
rect 36459 38848 36584 38876
rect 36730 38879 36788 38885
rect 36459 38845 36471 38848
rect 36413 38839 36471 38845
rect 36730 38845 36742 38879
rect 36776 38845 36788 38879
rect 37458 38876 37464 38888
rect 36730 38839 36788 38845
rect 36832 38848 37464 38876
rect 24452 38780 25452 38808
rect 24452 38768 24458 38780
rect 34514 38768 34520 38820
rect 34572 38808 34578 38820
rect 35250 38808 35256 38820
rect 34572 38780 35256 38808
rect 34572 38768 34578 38780
rect 35250 38768 35256 38780
rect 35308 38768 35314 38820
rect 35526 38768 35532 38820
rect 35584 38808 35590 38820
rect 36541 38811 36599 38817
rect 36541 38808 36553 38811
rect 35584 38780 36553 38808
rect 35584 38768 35590 38780
rect 36541 38777 36553 38780
rect 36587 38777 36599 38811
rect 36541 38771 36599 38777
rect 36630 38768 36636 38820
rect 36688 38808 36694 38820
rect 36832 38808 36860 38848
rect 37458 38836 37464 38848
rect 37516 38836 37522 38888
rect 37568 38885 37596 38916
rect 37553 38879 37611 38885
rect 37553 38845 37565 38879
rect 37599 38845 37611 38879
rect 37752 38876 37780 39052
rect 38102 39040 38108 39052
rect 38160 39040 38166 39092
rect 38010 38972 38016 39024
rect 38068 39012 38074 39024
rect 38068 38984 38240 39012
rect 38068 38972 38074 38984
rect 37921 38879 37979 38885
rect 37921 38876 37933 38879
rect 37752 38848 37933 38876
rect 37553 38839 37611 38845
rect 37921 38845 37933 38848
rect 37967 38845 37979 38879
rect 37921 38839 37979 38845
rect 37734 38808 37740 38820
rect 36688 38780 36860 38808
rect 37695 38780 37740 38808
rect 36688 38768 36694 38780
rect 37734 38768 37740 38780
rect 37792 38768 37798 38820
rect 37829 38811 37887 38817
rect 37829 38777 37841 38811
rect 37875 38808 37887 38811
rect 38212 38808 38240 38984
rect 37875 38780 38240 38808
rect 37875 38777 37887 38780
rect 37829 38771 37887 38777
rect 24026 38740 24032 38752
rect 23216 38712 24032 38740
rect 24026 38700 24032 38712
rect 24084 38700 24090 38752
rect 25314 38740 25320 38752
rect 25275 38712 25320 38740
rect 25314 38700 25320 38712
rect 25372 38700 25378 38752
rect 25498 38700 25504 38752
rect 25556 38740 25562 38752
rect 28721 38743 28779 38749
rect 28721 38740 28733 38743
rect 25556 38712 28733 38740
rect 25556 38700 25562 38712
rect 28721 38709 28733 38712
rect 28767 38709 28779 38743
rect 28721 38703 28779 38709
rect 30374 38700 30380 38752
rect 30432 38740 30438 38752
rect 31938 38740 31944 38752
rect 30432 38712 31944 38740
rect 30432 38700 30438 38712
rect 31938 38700 31944 38712
rect 31996 38700 32002 38752
rect 36909 38743 36967 38749
rect 36909 38709 36921 38743
rect 36955 38740 36967 38743
rect 37090 38740 37096 38752
rect 36955 38712 37096 38740
rect 36955 38709 36967 38712
rect 36909 38703 36967 38709
rect 37090 38700 37096 38712
rect 37148 38700 37154 38752
rect 37274 38700 37280 38752
rect 37332 38740 37338 38752
rect 38105 38743 38163 38749
rect 38105 38740 38117 38743
rect 37332 38712 38117 38740
rect 37332 38700 37338 38712
rect 38105 38709 38117 38712
rect 38151 38709 38163 38743
rect 38105 38703 38163 38709
rect 1104 38650 38824 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 38824 38650
rect 1104 38576 38824 38598
rect 22094 38496 22100 38548
rect 22152 38536 22158 38548
rect 22738 38536 22744 38548
rect 22152 38508 22744 38536
rect 22152 38496 22158 38508
rect 22738 38496 22744 38508
rect 22796 38496 22802 38548
rect 22941 38508 23152 38536
rect 1854 38468 1860 38480
rect 1815 38440 1860 38468
rect 1854 38428 1860 38440
rect 1912 38428 1918 38480
rect 2038 38468 2044 38480
rect 1999 38440 2044 38468
rect 2038 38428 2044 38440
rect 2096 38428 2102 38480
rect 17770 38428 17776 38480
rect 17828 38468 17834 38480
rect 22278 38468 22284 38480
rect 17828 38440 22284 38468
rect 17828 38428 17834 38440
rect 22278 38428 22284 38440
rect 22336 38428 22342 38480
rect 22941 38477 22969 38508
rect 22833 38471 22891 38477
rect 22833 38468 22845 38471
rect 22388 38440 22845 38468
rect 22002 38360 22008 38412
rect 22060 38400 22066 38412
rect 22388 38400 22416 38440
rect 22833 38437 22845 38440
rect 22879 38437 22891 38471
rect 22833 38431 22891 38437
rect 22925 38471 22983 38477
rect 22925 38437 22937 38471
rect 22971 38437 22983 38471
rect 23124 38468 23152 38508
rect 23382 38496 23388 38548
rect 23440 38536 23446 38548
rect 23440 38508 31754 38536
rect 23440 38496 23446 38508
rect 23474 38468 23480 38480
rect 23124 38440 23480 38468
rect 22925 38431 22983 38437
rect 23474 38428 23480 38440
rect 23532 38428 23538 38480
rect 24112 38471 24170 38477
rect 24112 38437 24124 38471
rect 24158 38468 24170 38471
rect 25314 38468 25320 38480
rect 24158 38440 25320 38468
rect 24158 38437 24170 38440
rect 24112 38431 24170 38437
rect 25314 38428 25320 38440
rect 25372 38428 25378 38480
rect 26418 38468 26424 38480
rect 26331 38440 26424 38468
rect 26418 38428 26424 38440
rect 26476 38468 26482 38480
rect 26476 38440 26740 38468
rect 26476 38428 26482 38440
rect 22554 38400 22560 38412
rect 22060 38372 22416 38400
rect 22515 38372 22560 38400
rect 22060 38360 22066 38372
rect 22554 38360 22560 38372
rect 22612 38360 22618 38412
rect 22695 38403 22753 38409
rect 22695 38369 22707 38403
rect 22741 38369 22753 38403
rect 22695 38363 22753 38369
rect 23063 38403 23121 38409
rect 23063 38369 23075 38403
rect 23109 38400 23121 38403
rect 23198 38400 23204 38412
rect 23109 38372 23204 38400
rect 23109 38369 23121 38372
rect 23063 38363 23121 38369
rect 6362 38292 6368 38344
rect 6420 38332 6426 38344
rect 22278 38332 22284 38344
rect 6420 38304 22284 38332
rect 6420 38292 6426 38304
rect 22278 38292 22284 38304
rect 22336 38292 22342 38344
rect 22720 38276 22748 38363
rect 23198 38360 23204 38372
rect 23256 38360 23262 38412
rect 23382 38360 23388 38412
rect 23440 38400 23446 38412
rect 24486 38400 24492 38412
rect 23440 38372 24492 38400
rect 23440 38360 23446 38372
rect 24486 38360 24492 38372
rect 24544 38360 24550 38412
rect 25866 38360 25872 38412
rect 25924 38400 25930 38412
rect 26237 38403 26295 38409
rect 26237 38400 26249 38403
rect 25924 38372 26249 38400
rect 25924 38360 25930 38372
rect 26237 38369 26249 38372
rect 26283 38369 26295 38403
rect 26510 38400 26516 38412
rect 26471 38372 26516 38400
rect 26237 38363 26295 38369
rect 26510 38360 26516 38372
rect 26568 38360 26574 38412
rect 26610 38403 26668 38409
rect 26610 38369 26622 38403
rect 26656 38369 26668 38403
rect 26712 38400 26740 38440
rect 27338 38428 27344 38480
rect 27396 38468 27402 38480
rect 31478 38468 31484 38480
rect 27396 38440 31484 38468
rect 27396 38428 27402 38440
rect 31478 38428 31484 38440
rect 31536 38428 31542 38480
rect 31726 38468 31754 38508
rect 34606 38496 34612 38548
rect 34664 38536 34670 38548
rect 34793 38539 34851 38545
rect 34793 38536 34805 38539
rect 34664 38508 34805 38536
rect 34664 38496 34670 38508
rect 34793 38505 34805 38508
rect 34839 38505 34851 38539
rect 34793 38499 34851 38505
rect 35437 38539 35495 38545
rect 35437 38505 35449 38539
rect 35483 38536 35495 38539
rect 35618 38536 35624 38548
rect 35483 38508 35624 38536
rect 35483 38505 35495 38508
rect 35437 38499 35495 38505
rect 35618 38496 35624 38508
rect 35676 38496 35682 38548
rect 36265 38539 36323 38545
rect 36265 38505 36277 38539
rect 36311 38536 36323 38539
rect 38010 38536 38016 38548
rect 36311 38508 38016 38536
rect 36311 38505 36323 38508
rect 36265 38499 36323 38505
rect 37001 38471 37059 38477
rect 37001 38468 37013 38471
rect 31726 38440 37013 38468
rect 37001 38437 37013 38440
rect 37047 38437 37059 38471
rect 37001 38431 37059 38437
rect 27890 38400 27896 38412
rect 26712 38372 27896 38400
rect 26610 38363 26668 38369
rect 23290 38292 23296 38344
rect 23348 38332 23354 38344
rect 23845 38335 23903 38341
rect 23845 38332 23857 38335
rect 23348 38304 23857 38332
rect 23348 38292 23354 38304
rect 23845 38301 23857 38304
rect 23891 38301 23903 38335
rect 26625 38332 26653 38363
rect 27890 38360 27896 38372
rect 27948 38360 27954 38412
rect 28810 38360 28816 38412
rect 28868 38400 28874 38412
rect 28905 38403 28963 38409
rect 28905 38400 28917 38403
rect 28868 38372 28917 38400
rect 28868 38360 28874 38372
rect 28905 38369 28917 38372
rect 28951 38369 28963 38403
rect 28905 38363 28963 38369
rect 29089 38403 29147 38409
rect 29089 38369 29101 38403
rect 29135 38400 29147 38403
rect 29270 38400 29276 38412
rect 29135 38372 29276 38400
rect 29135 38369 29147 38372
rect 29089 38363 29147 38369
rect 29270 38360 29276 38372
rect 29328 38360 29334 38412
rect 29365 38403 29423 38409
rect 29365 38369 29377 38403
rect 29411 38400 29423 38403
rect 29454 38400 29460 38412
rect 29411 38372 29460 38400
rect 29411 38369 29423 38372
rect 29365 38363 29423 38369
rect 29454 38360 29460 38372
rect 29512 38360 29518 38412
rect 34977 38403 35035 38409
rect 34977 38369 34989 38403
rect 35023 38400 35035 38403
rect 35342 38400 35348 38412
rect 35023 38372 35348 38400
rect 35023 38369 35035 38372
rect 34977 38363 35035 38369
rect 35342 38360 35348 38372
rect 35400 38360 35406 38412
rect 35621 38403 35679 38409
rect 35621 38369 35633 38403
rect 35667 38400 35679 38403
rect 35710 38400 35716 38412
rect 35667 38372 35716 38400
rect 35667 38369 35679 38372
rect 35621 38363 35679 38369
rect 35710 38360 35716 38372
rect 35768 38360 35774 38412
rect 35986 38360 35992 38412
rect 36044 38400 36050 38412
rect 36173 38403 36231 38409
rect 36173 38400 36185 38403
rect 36044 38372 36185 38400
rect 36044 38360 36050 38372
rect 36173 38369 36185 38372
rect 36219 38369 36231 38403
rect 36173 38363 36231 38369
rect 36538 38360 36544 38412
rect 36596 38400 36602 38412
rect 36722 38400 36728 38412
rect 36596 38372 36728 38400
rect 36596 38360 36602 38372
rect 36722 38360 36728 38372
rect 36780 38360 36786 38412
rect 36817 38403 36875 38409
rect 36817 38369 36829 38403
rect 36863 38400 36875 38403
rect 36906 38400 36912 38412
rect 36863 38372 36912 38400
rect 36863 38369 36875 38372
rect 36817 38363 36875 38369
rect 36906 38360 36912 38372
rect 36964 38360 36970 38412
rect 37200 38409 37228 38508
rect 38010 38496 38016 38508
rect 38068 38496 38074 38548
rect 37093 38403 37151 38409
rect 37093 38369 37105 38403
rect 37139 38369 37151 38403
rect 37093 38363 37151 38369
rect 37185 38403 37243 38409
rect 37185 38369 37197 38403
rect 37231 38369 37243 38403
rect 37185 38363 37243 38369
rect 23845 38295 23903 38301
rect 24872 38304 26653 38332
rect 1578 38224 1584 38276
rect 1636 38264 1642 38276
rect 1636 38236 19334 38264
rect 22720 38236 22744 38276
rect 1636 38224 1642 38236
rect 19306 38196 19334 38236
rect 22738 38224 22744 38236
rect 22796 38224 22802 38276
rect 23201 38267 23259 38273
rect 23201 38233 23213 38267
rect 23247 38264 23259 38267
rect 23382 38264 23388 38276
rect 23247 38236 23388 38264
rect 23247 38233 23259 38236
rect 23201 38227 23259 38233
rect 23382 38224 23388 38236
rect 23440 38224 23446 38276
rect 24872 38196 24900 38304
rect 29178 38292 29184 38344
rect 29236 38332 29242 38344
rect 29236 38304 29281 38332
rect 29236 38292 29242 38304
rect 35526 38292 35532 38344
rect 35584 38332 35590 38344
rect 37108 38332 37136 38363
rect 37366 38332 37372 38344
rect 35584 38304 37136 38332
rect 37200 38304 37372 38332
rect 35584 38292 35590 38304
rect 26326 38224 26332 38276
rect 26384 38264 26390 38276
rect 26789 38267 26847 38273
rect 26789 38264 26801 38267
rect 26384 38236 26801 38264
rect 26384 38224 26390 38236
rect 26789 38233 26801 38236
rect 26835 38233 26847 38267
rect 26789 38227 26847 38233
rect 28997 38267 29055 38273
rect 28997 38233 29009 38267
rect 29043 38264 29055 38267
rect 29730 38264 29736 38276
rect 29043 38236 29736 38264
rect 29043 38233 29055 38236
rect 28997 38227 29055 38233
rect 29730 38224 29736 38236
rect 29788 38224 29794 38276
rect 34606 38224 34612 38276
rect 34664 38264 34670 38276
rect 34974 38264 34980 38276
rect 34664 38236 34980 38264
rect 34664 38224 34670 38236
rect 34974 38224 34980 38236
rect 35032 38224 35038 38276
rect 35986 38224 35992 38276
rect 36044 38264 36050 38276
rect 37200 38264 37228 38304
rect 37366 38292 37372 38304
rect 37424 38292 37430 38344
rect 36044 38236 37228 38264
rect 36044 38224 36050 38236
rect 25222 38196 25228 38208
rect 19306 38168 24900 38196
rect 25183 38168 25228 38196
rect 25222 38156 25228 38168
rect 25280 38156 25286 38208
rect 25314 38156 25320 38208
rect 25372 38196 25378 38208
rect 27154 38196 27160 38208
rect 25372 38168 27160 38196
rect 25372 38156 25378 38168
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 27890 38156 27896 38208
rect 27948 38196 27954 38208
rect 28721 38199 28779 38205
rect 28721 38196 28733 38199
rect 27948 38168 28733 38196
rect 27948 38156 27954 38168
rect 28721 38165 28733 38168
rect 28767 38165 28779 38199
rect 28721 38159 28779 38165
rect 36630 38156 36636 38208
rect 36688 38196 36694 38208
rect 37369 38199 37427 38205
rect 37369 38196 37381 38199
rect 36688 38168 37381 38196
rect 36688 38156 36694 38168
rect 37369 38165 37381 38168
rect 37415 38165 37427 38199
rect 37369 38159 37427 38165
rect 1104 38106 38824 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 38824 38106
rect 1104 38032 38824 38054
rect 2498 37952 2504 38004
rect 2556 37992 2562 38004
rect 26602 37992 26608 38004
rect 2556 37964 26608 37992
rect 2556 37952 2562 37964
rect 26602 37952 26608 37964
rect 26660 37952 26666 38004
rect 26786 37992 26792 38004
rect 26747 37964 26792 37992
rect 26786 37952 26792 37964
rect 26844 37952 26850 38004
rect 28442 37952 28448 38004
rect 28500 37992 28506 38004
rect 28500 37964 30512 37992
rect 28500 37952 28506 37964
rect 2041 37927 2099 37933
rect 2041 37893 2053 37927
rect 2087 37924 2099 37927
rect 2130 37924 2136 37936
rect 2087 37896 2136 37924
rect 2087 37893 2099 37896
rect 2041 37887 2099 37893
rect 2130 37884 2136 37896
rect 2188 37884 2194 37936
rect 21910 37924 21916 37936
rect 6886 37896 21916 37924
rect 1670 37816 1676 37868
rect 1728 37856 1734 37868
rect 6886 37856 6914 37896
rect 21910 37884 21916 37896
rect 21968 37884 21974 37936
rect 22373 37927 22431 37933
rect 22373 37924 22385 37927
rect 22296 37896 22385 37924
rect 22296 37868 22324 37896
rect 22373 37893 22385 37896
rect 22419 37893 22431 37927
rect 22373 37887 22431 37893
rect 23477 37927 23535 37933
rect 23477 37893 23489 37927
rect 23523 37893 23535 37927
rect 23477 37887 23535 37893
rect 1728 37828 6914 37856
rect 1728 37816 1734 37828
rect 18046 37816 18052 37868
rect 18104 37856 18110 37868
rect 18104 37828 22094 37856
rect 18104 37816 18110 37828
rect 21726 37788 21732 37800
rect 21687 37760 21732 37788
rect 21726 37748 21732 37760
rect 21784 37748 21790 37800
rect 21910 37797 21916 37800
rect 21877 37791 21916 37797
rect 21877 37757 21889 37791
rect 21877 37751 21916 37757
rect 21910 37748 21916 37751
rect 21968 37748 21974 37800
rect 22066 37788 22094 37828
rect 22278 37816 22284 37868
rect 22336 37816 22342 37868
rect 23492 37856 23520 37887
rect 24210 37884 24216 37936
rect 24268 37924 24274 37936
rect 24268 37896 26653 37924
rect 24268 37884 24274 37896
rect 25314 37856 25320 37868
rect 22388 37828 22969 37856
rect 23492 37828 25320 37856
rect 22388 37800 22416 37828
rect 22194 37791 22252 37797
rect 22194 37788 22206 37791
rect 22066 37760 22206 37788
rect 22194 37757 22206 37760
rect 22240 37757 22252 37791
rect 22194 37751 22252 37757
rect 22370 37748 22376 37800
rect 22428 37748 22434 37800
rect 22462 37748 22468 37800
rect 22520 37788 22526 37800
rect 22941 37797 22969 37828
rect 25314 37816 25320 37828
rect 25372 37816 25378 37868
rect 26326 37856 26332 37868
rect 26252 37828 26332 37856
rect 22833 37791 22891 37797
rect 22833 37788 22845 37791
rect 22520 37760 22845 37788
rect 22520 37748 22526 37760
rect 22833 37757 22845 37760
rect 22879 37757 22891 37791
rect 22833 37751 22891 37757
rect 22926 37791 22984 37797
rect 22926 37757 22938 37791
rect 22972 37757 22984 37791
rect 22926 37751 22984 37757
rect 23290 37748 23296 37800
rect 23348 37797 23354 37800
rect 23348 37788 23356 37797
rect 23348 37760 23393 37788
rect 23348 37751 23356 37760
rect 23348 37748 23354 37751
rect 23474 37748 23480 37800
rect 23532 37788 23538 37800
rect 24121 37791 24179 37797
rect 24121 37788 24133 37791
rect 23532 37760 24133 37788
rect 23532 37748 23538 37760
rect 24121 37757 24133 37760
rect 24167 37757 24179 37791
rect 24121 37751 24179 37757
rect 24305 37791 24363 37797
rect 24305 37757 24317 37791
rect 24351 37788 24363 37791
rect 24394 37788 24400 37800
rect 24351 37760 24400 37788
rect 24351 37757 24363 37760
rect 24305 37751 24363 37757
rect 24394 37748 24400 37760
rect 24452 37748 24458 37800
rect 26252 37797 26280 37828
rect 26326 37816 26332 37828
rect 26384 37816 26390 37868
rect 26237 37791 26295 37797
rect 26237 37757 26249 37791
rect 26283 37757 26295 37791
rect 26510 37788 26516 37800
rect 26471 37760 26516 37788
rect 26237 37751 26295 37757
rect 26510 37748 26516 37760
rect 26568 37748 26574 37800
rect 26625 37797 26653 37896
rect 28626 37884 28632 37936
rect 28684 37924 28690 37936
rect 28813 37927 28871 37933
rect 28813 37924 28825 37927
rect 28684 37896 28825 37924
rect 28684 37884 28690 37896
rect 28813 37893 28825 37896
rect 28859 37893 28871 37927
rect 30374 37924 30380 37936
rect 28813 37887 28871 37893
rect 28920 37896 30380 37924
rect 28442 37816 28448 37868
rect 28500 37856 28506 37868
rect 28920 37865 28948 37896
rect 30374 37884 30380 37896
rect 30432 37884 30438 37936
rect 28905 37859 28963 37865
rect 28500 37828 28764 37856
rect 28500 37816 28506 37828
rect 26610 37791 26668 37797
rect 26610 37757 26622 37791
rect 26656 37757 26668 37791
rect 26610 37751 26668 37757
rect 28258 37748 28264 37800
rect 28316 37788 28322 37800
rect 28626 37788 28632 37800
rect 28316 37760 28632 37788
rect 28316 37748 28322 37760
rect 28626 37748 28632 37760
rect 28684 37748 28690 37800
rect 28736 37797 28764 37828
rect 28905 37825 28917 37859
rect 28951 37825 28963 37859
rect 28905 37819 28963 37825
rect 28997 37859 29055 37865
rect 28997 37825 29009 37859
rect 29043 37856 29055 37859
rect 29270 37856 29276 37868
rect 29043 37828 29276 37856
rect 29043 37825 29055 37828
rect 28997 37819 29055 37825
rect 29270 37816 29276 37828
rect 29328 37816 29334 37868
rect 29914 37816 29920 37868
rect 29972 37856 29978 37868
rect 30282 37856 30288 37868
rect 29972 37828 30288 37856
rect 29972 37816 29978 37828
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 28721 37791 28779 37797
rect 28721 37757 28733 37791
rect 28767 37757 28779 37791
rect 28721 37751 28779 37757
rect 29086 37748 29092 37800
rect 29144 37788 29150 37800
rect 29181 37791 29239 37797
rect 29181 37788 29193 37791
rect 29144 37760 29193 37788
rect 29144 37748 29150 37760
rect 29181 37757 29193 37760
rect 29227 37788 29239 37791
rect 29454 37788 29460 37800
rect 29227 37760 29460 37788
rect 29227 37757 29239 37760
rect 29181 37751 29239 37757
rect 29454 37748 29460 37760
rect 29512 37748 29518 37800
rect 1854 37720 1860 37732
rect 1815 37692 1860 37720
rect 1854 37680 1860 37692
rect 1912 37680 1918 37732
rect 22002 37720 22008 37732
rect 21915 37692 22008 37720
rect 22002 37680 22008 37692
rect 22060 37680 22066 37732
rect 22097 37723 22155 37729
rect 22097 37689 22109 37723
rect 22143 37720 22155 37723
rect 22278 37720 22284 37732
rect 22143 37692 22284 37720
rect 22143 37689 22155 37692
rect 22097 37683 22155 37689
rect 22278 37680 22284 37692
rect 22336 37680 22342 37732
rect 23109 37723 23167 37729
rect 23109 37720 23121 37723
rect 22388 37692 23121 37720
rect 22020 37652 22048 37680
rect 22388 37652 22416 37692
rect 23109 37689 23121 37692
rect 23155 37689 23167 37723
rect 23109 37683 23167 37689
rect 23201 37723 23259 37729
rect 23201 37689 23213 37723
rect 23247 37720 23259 37723
rect 23382 37720 23388 37732
rect 23247 37692 23388 37720
rect 23247 37689 23259 37692
rect 23201 37683 23259 37689
rect 22020 37624 22416 37652
rect 22554 37612 22560 37664
rect 22612 37652 22618 37664
rect 22830 37652 22836 37664
rect 22612 37624 22836 37652
rect 22612 37612 22618 37624
rect 22830 37612 22836 37624
rect 22888 37612 22894 37664
rect 23124 37652 23152 37683
rect 23382 37680 23388 37692
rect 23440 37680 23446 37732
rect 24854 37720 24860 37732
rect 23492 37692 24860 37720
rect 23492 37652 23520 37692
rect 24854 37680 24860 37692
rect 24912 37680 24918 37732
rect 26418 37720 26424 37732
rect 26379 37692 26424 37720
rect 26418 37680 26424 37692
rect 26476 37680 26482 37732
rect 30282 37720 30288 37732
rect 26611 37692 30288 37720
rect 24210 37652 24216 37664
rect 23124 37624 23520 37652
rect 24171 37624 24216 37652
rect 24210 37612 24216 37624
rect 24268 37612 24274 37664
rect 24670 37612 24676 37664
rect 24728 37652 24734 37664
rect 26611 37652 26639 37692
rect 30282 37680 30288 37692
rect 30340 37680 30346 37732
rect 24728 37624 26639 37652
rect 24728 37612 24734 37624
rect 28442 37612 28448 37664
rect 28500 37652 28506 37664
rect 28537 37655 28595 37661
rect 28537 37652 28549 37655
rect 28500 37624 28549 37652
rect 28500 37612 28506 37624
rect 28537 37621 28549 37624
rect 28583 37621 28595 37655
rect 28537 37615 28595 37621
rect 28902 37612 28908 37664
rect 28960 37652 28966 37664
rect 30374 37652 30380 37664
rect 28960 37624 30380 37652
rect 28960 37612 28966 37624
rect 30374 37612 30380 37624
rect 30432 37612 30438 37664
rect 30484 37652 30512 37964
rect 30834 37952 30840 38004
rect 30892 37952 30898 38004
rect 36357 37995 36415 38001
rect 36357 37961 36369 37995
rect 36403 37992 36415 37995
rect 36906 37992 36912 38004
rect 36403 37964 36912 37992
rect 36403 37961 36415 37964
rect 36357 37955 36415 37961
rect 36906 37952 36912 37964
rect 36964 37952 36970 38004
rect 30650 37680 30656 37732
rect 30708 37720 30714 37732
rect 30852 37720 30880 37952
rect 35710 37884 35716 37936
rect 35768 37924 35774 37936
rect 38105 37927 38163 37933
rect 38105 37924 38117 37927
rect 35768 37896 38117 37924
rect 35768 37884 35774 37896
rect 38105 37893 38117 37896
rect 38151 37893 38163 37927
rect 38105 37887 38163 37893
rect 31478 37816 31484 37868
rect 31536 37856 31542 37868
rect 38470 37856 38476 37868
rect 31536 37828 37596 37856
rect 31536 37816 31542 37828
rect 36170 37788 36176 37800
rect 36131 37760 36176 37788
rect 36170 37748 36176 37760
rect 36228 37748 36234 37800
rect 37568 37797 37596 37828
rect 37660 37828 38476 37856
rect 36909 37791 36967 37797
rect 36909 37757 36921 37791
rect 36955 37788 36967 37791
rect 37553 37791 37611 37797
rect 36955 37760 37504 37788
rect 36955 37757 36967 37760
rect 36909 37751 36967 37757
rect 37090 37720 37096 37732
rect 30708 37692 30880 37720
rect 37051 37692 37096 37720
rect 30708 37680 30714 37692
rect 37090 37680 37096 37692
rect 37148 37680 37154 37732
rect 37476 37720 37504 37760
rect 37553 37757 37565 37791
rect 37599 37757 37611 37791
rect 37553 37751 37611 37757
rect 37660 37720 37688 37828
rect 38470 37816 38476 37828
rect 38528 37816 38534 37868
rect 37734 37748 37740 37800
rect 37792 37788 37798 37800
rect 37921 37791 37979 37797
rect 37792 37760 37837 37788
rect 37792 37748 37798 37760
rect 37921 37757 37933 37791
rect 37967 37788 37979 37791
rect 38286 37788 38292 37800
rect 37967 37760 38292 37788
rect 37967 37757 37979 37760
rect 37921 37751 37979 37757
rect 38286 37748 38292 37760
rect 38344 37748 38350 37800
rect 37476 37692 37688 37720
rect 37829 37723 37887 37729
rect 37829 37689 37841 37723
rect 37875 37689 37887 37723
rect 37829 37683 37887 37689
rect 35158 37652 35164 37664
rect 30484 37624 35164 37652
rect 35158 37612 35164 37624
rect 35216 37612 35222 37664
rect 35342 37612 35348 37664
rect 35400 37652 35406 37664
rect 35526 37652 35532 37664
rect 35400 37624 35532 37652
rect 35400 37612 35406 37624
rect 35526 37612 35532 37624
rect 35584 37612 35590 37664
rect 35986 37612 35992 37664
rect 36044 37652 36050 37664
rect 36170 37652 36176 37664
rect 36044 37624 36176 37652
rect 36044 37612 36050 37624
rect 36170 37612 36176 37624
rect 36228 37612 36234 37664
rect 37366 37612 37372 37664
rect 37424 37652 37430 37664
rect 37844 37652 37872 37683
rect 37424 37624 37872 37652
rect 37424 37612 37430 37624
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 24670 37448 24676 37460
rect 19306 37420 24676 37448
rect 17862 37272 17868 37324
rect 17920 37312 17926 37324
rect 19306 37312 19334 37420
rect 24670 37408 24676 37420
rect 24728 37408 24734 37460
rect 24780 37420 28028 37448
rect 21542 37340 21548 37392
rect 21600 37380 21606 37392
rect 21600 37352 23980 37380
rect 21600 37340 21606 37352
rect 17920 37284 19334 37312
rect 17920 37272 17926 37284
rect 22830 37272 22836 37324
rect 22888 37312 22894 37324
rect 22925 37315 22983 37321
rect 22925 37312 22937 37315
rect 22888 37284 22937 37312
rect 22888 37272 22894 37284
rect 22925 37281 22937 37284
rect 22971 37281 22983 37315
rect 22925 37275 22983 37281
rect 23201 37315 23259 37321
rect 23201 37281 23213 37315
rect 23247 37312 23259 37315
rect 23382 37312 23388 37324
rect 23247 37284 23388 37312
rect 23247 37281 23259 37284
rect 23201 37275 23259 37281
rect 23382 37272 23388 37284
rect 23440 37272 23446 37324
rect 21726 37204 21732 37256
rect 21784 37244 21790 37256
rect 23566 37244 23572 37256
rect 21784 37216 23336 37244
rect 23527 37216 23572 37244
rect 21784 37204 21790 37216
rect 20346 37136 20352 37188
rect 20404 37176 20410 37188
rect 22554 37176 22560 37188
rect 20404 37148 22560 37176
rect 20404 37136 20410 37148
rect 22554 37136 22560 37148
rect 22612 37136 22618 37188
rect 23017 37179 23075 37185
rect 23017 37145 23029 37179
rect 23063 37176 23075 37179
rect 23198 37176 23204 37188
rect 23063 37148 23204 37176
rect 23063 37145 23075 37148
rect 23017 37139 23075 37145
rect 23198 37136 23204 37148
rect 23256 37136 23262 37188
rect 23308 37176 23336 37216
rect 23566 37204 23572 37216
rect 23624 37204 23630 37256
rect 23952 37244 23980 37352
rect 24026 37340 24032 37392
rect 24084 37380 24090 37392
rect 24121 37383 24179 37389
rect 24121 37380 24133 37383
rect 24084 37352 24133 37380
rect 24084 37340 24090 37352
rect 24121 37349 24133 37352
rect 24167 37349 24179 37383
rect 24121 37343 24179 37349
rect 24302 37340 24308 37392
rect 24360 37389 24366 37392
rect 24360 37383 24384 37389
rect 24372 37349 24384 37383
rect 24360 37343 24384 37349
rect 24360 37340 24366 37343
rect 24780 37312 24808 37420
rect 26418 37380 26424 37392
rect 26379 37352 26424 37380
rect 26418 37340 26424 37352
rect 26476 37340 26482 37392
rect 26513 37383 26571 37389
rect 26513 37349 26525 37383
rect 26559 37349 26571 37383
rect 28000 37380 28028 37420
rect 28074 37408 28080 37460
rect 28132 37448 28138 37460
rect 28353 37451 28411 37457
rect 28353 37448 28365 37451
rect 28132 37420 28365 37448
rect 28132 37408 28138 37420
rect 28353 37417 28365 37420
rect 28399 37417 28411 37451
rect 29454 37448 29460 37460
rect 28353 37411 28411 37417
rect 28644 37420 29460 37448
rect 28644 37380 28672 37420
rect 29454 37408 29460 37420
rect 29512 37408 29518 37460
rect 30374 37408 30380 37460
rect 30432 37448 30438 37460
rect 32306 37448 32312 37460
rect 30432 37420 32312 37448
rect 30432 37408 30438 37420
rect 32306 37408 32312 37420
rect 32364 37408 32370 37460
rect 35158 37408 35164 37460
rect 35216 37448 35222 37460
rect 35713 37451 35771 37457
rect 35713 37448 35725 37451
rect 35216 37420 35725 37448
rect 35216 37408 35222 37420
rect 35713 37417 35725 37420
rect 35759 37417 35771 37451
rect 35713 37411 35771 37417
rect 36173 37451 36231 37457
rect 36173 37417 36185 37451
rect 36219 37448 36231 37451
rect 36354 37448 36360 37460
rect 36219 37420 36360 37448
rect 36219 37417 36231 37420
rect 36173 37411 36231 37417
rect 36354 37408 36360 37420
rect 36412 37408 36418 37460
rect 28000 37352 28672 37380
rect 28736 37352 30236 37380
rect 26513 37343 26571 37349
rect 24228 37284 24808 37312
rect 26237 37315 26295 37321
rect 24228 37244 24256 37284
rect 26237 37281 26249 37315
rect 26283 37281 26295 37315
rect 26237 37275 26295 37281
rect 23952 37216 24256 37244
rect 24489 37179 24547 37185
rect 24489 37176 24501 37179
rect 23308 37148 24501 37176
rect 24489 37145 24501 37148
rect 24535 37145 24547 37179
rect 24489 37139 24547 37145
rect 23566 37068 23572 37120
rect 23624 37108 23630 37120
rect 24305 37111 24363 37117
rect 24305 37108 24317 37111
rect 23624 37080 24317 37108
rect 23624 37068 23630 37080
rect 24305 37077 24317 37080
rect 24351 37077 24363 37111
rect 26252 37108 26280 37275
rect 26528 37274 26556 37343
rect 26528 37256 26557 37274
rect 26602 37272 26608 37324
rect 26660 37321 26666 37324
rect 26660 37312 26668 37321
rect 26878 37312 26884 37324
rect 26660 37284 26705 37312
rect 26804 37284 26884 37312
rect 26660 37275 26668 37284
rect 26660 37272 26666 37275
rect 26510 37204 26516 37256
rect 26568 37204 26574 37256
rect 26804 37185 26832 37284
rect 26878 37272 26884 37284
rect 26936 37272 26942 37324
rect 28736 37321 28764 37352
rect 28537 37315 28595 37321
rect 28537 37281 28549 37315
rect 28583 37281 28595 37315
rect 28537 37275 28595 37281
rect 28721 37315 28779 37321
rect 28721 37281 28733 37315
rect 28767 37281 28779 37315
rect 28721 37275 28779 37281
rect 28813 37315 28871 37321
rect 28813 37281 28825 37315
rect 28859 37312 28871 37315
rect 28902 37312 28908 37324
rect 28859 37284 28908 37312
rect 28859 37281 28871 37284
rect 28813 37275 28871 37281
rect 28552 37244 28580 37275
rect 28902 37272 28908 37284
rect 28960 37272 28966 37324
rect 28997 37315 29055 37321
rect 28997 37281 29009 37315
rect 29043 37312 29055 37315
rect 29086 37312 29092 37324
rect 29043 37284 29092 37312
rect 29043 37281 29055 37284
rect 28997 37275 29055 37281
rect 29086 37272 29092 37284
rect 29144 37272 29150 37324
rect 29454 37272 29460 37324
rect 29512 37312 29518 37324
rect 29641 37315 29699 37321
rect 29641 37312 29653 37315
rect 29512 37284 29653 37312
rect 29512 37272 29518 37284
rect 29641 37281 29653 37284
rect 29687 37281 29699 37315
rect 29822 37312 29828 37324
rect 29783 37284 29828 37312
rect 29641 37275 29699 37281
rect 29822 37272 29828 37284
rect 29880 37272 29886 37324
rect 30006 37272 30012 37324
rect 30064 37312 30070 37324
rect 30101 37315 30159 37321
rect 30101 37312 30113 37315
rect 30064 37284 30113 37312
rect 30064 37272 30070 37284
rect 30101 37281 30113 37284
rect 30147 37281 30159 37315
rect 30101 37275 30159 37281
rect 29730 37244 29736 37256
rect 26896 37216 28580 37244
rect 29691 37216 29736 37244
rect 26896 37188 26924 37216
rect 29730 37204 29736 37216
rect 29788 37204 29794 37256
rect 29917 37247 29975 37253
rect 29917 37213 29929 37247
rect 29963 37213 29975 37247
rect 30208 37244 30236 37352
rect 30282 37340 30288 37392
rect 30340 37380 30346 37392
rect 37093 37383 37151 37389
rect 30340 37352 31432 37380
rect 30340 37340 30346 37352
rect 31404 37312 31432 37352
rect 31588 37352 36860 37380
rect 31588 37312 31616 37352
rect 35526 37312 35532 37324
rect 31404 37284 31616 37312
rect 35487 37284 35532 37312
rect 35526 37272 35532 37284
rect 35584 37272 35590 37324
rect 36354 37312 36360 37324
rect 36315 37284 36360 37312
rect 36354 37272 36360 37284
rect 36412 37272 36418 37324
rect 36832 37321 36860 37352
rect 37093 37349 37105 37383
rect 37139 37380 37151 37383
rect 37366 37380 37372 37392
rect 37139 37352 37372 37380
rect 37139 37349 37151 37352
rect 37093 37343 37151 37349
rect 37366 37340 37372 37352
rect 37424 37340 37430 37392
rect 36817 37315 36875 37321
rect 36817 37281 36829 37315
rect 36863 37281 36875 37315
rect 36817 37275 36875 37281
rect 37001 37315 37059 37321
rect 37001 37281 37013 37315
rect 37047 37281 37059 37315
rect 37001 37275 37059 37281
rect 37185 37315 37243 37321
rect 37185 37281 37197 37315
rect 37231 37312 37243 37315
rect 38470 37312 38476 37324
rect 37231 37284 38476 37312
rect 37231 37281 37243 37284
rect 37185 37275 37243 37281
rect 31846 37244 31852 37256
rect 30208 37216 31852 37244
rect 29917 37207 29975 37213
rect 26789 37179 26847 37185
rect 26789 37145 26801 37179
rect 26835 37145 26847 37179
rect 26789 37139 26847 37145
rect 26878 37136 26884 37188
rect 26936 37136 26942 37188
rect 27706 37136 27712 37188
rect 27764 37176 27770 37188
rect 28629 37179 28687 37185
rect 28629 37176 28641 37179
rect 27764 37148 28641 37176
rect 27764 37136 27770 37148
rect 28629 37145 28641 37148
rect 28675 37145 28687 37179
rect 29932 37176 29960 37207
rect 31846 37204 31852 37216
rect 31904 37204 31910 37256
rect 35618 37204 35624 37256
rect 35676 37244 35682 37256
rect 37016 37244 37044 37275
rect 38470 37272 38476 37284
rect 38528 37272 38534 37324
rect 37734 37244 37740 37256
rect 35676 37216 37740 37244
rect 35676 37204 35682 37216
rect 37734 37204 37740 37216
rect 37792 37204 37798 37256
rect 28629 37139 28687 37145
rect 29748 37148 29960 37176
rect 29748 37120 29776 37148
rect 35986 37136 35992 37188
rect 36044 37176 36050 37188
rect 38746 37176 38752 37188
rect 36044 37148 38752 37176
rect 36044 37136 36050 37148
rect 38746 37136 38752 37148
rect 38804 37136 38810 37188
rect 27338 37108 27344 37120
rect 26252 37080 27344 37108
rect 24305 37071 24363 37077
rect 27338 37068 27344 37080
rect 27396 37068 27402 37120
rect 28258 37068 28264 37120
rect 28316 37108 28322 37120
rect 29457 37111 29515 37117
rect 29457 37108 29469 37111
rect 28316 37080 29469 37108
rect 28316 37068 28322 37080
rect 29457 37077 29469 37080
rect 29503 37077 29515 37111
rect 29457 37071 29515 37077
rect 29730 37068 29736 37120
rect 29788 37068 29794 37120
rect 36906 37068 36912 37120
rect 36964 37108 36970 37120
rect 37369 37111 37427 37117
rect 37369 37108 37381 37111
rect 36964 37080 37381 37108
rect 36964 37068 36970 37080
rect 37369 37077 37381 37080
rect 37415 37077 37427 37111
rect 37369 37071 37427 37077
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 1578 36904 1584 36916
rect 1539 36876 1584 36904
rect 1578 36864 1584 36876
rect 1636 36864 1642 36916
rect 23474 36904 23480 36916
rect 23435 36876 23480 36904
rect 23474 36864 23480 36876
rect 23532 36864 23538 36916
rect 23566 36864 23572 36916
rect 23624 36904 23630 36916
rect 25222 36904 25228 36916
rect 23624 36876 25228 36904
rect 23624 36864 23630 36876
rect 25222 36864 25228 36876
rect 25280 36864 25286 36916
rect 26326 36864 26332 36916
rect 26384 36904 26390 36916
rect 26602 36904 26608 36916
rect 26384 36876 26608 36904
rect 26384 36864 26390 36876
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 26694 36864 26700 36916
rect 26752 36904 26758 36916
rect 26789 36907 26847 36913
rect 26789 36904 26801 36907
rect 26752 36876 26801 36904
rect 26752 36864 26758 36876
rect 26789 36873 26801 36876
rect 26835 36873 26847 36907
rect 26789 36867 26847 36873
rect 29454 36864 29460 36916
rect 29512 36904 29518 36916
rect 31386 36904 31392 36916
rect 29512 36876 31392 36904
rect 29512 36864 29518 36876
rect 31386 36864 31392 36876
rect 31444 36864 31450 36916
rect 35713 36907 35771 36913
rect 35713 36873 35725 36907
rect 35759 36904 35771 36907
rect 35894 36904 35900 36916
rect 35759 36876 35900 36904
rect 35759 36873 35771 36876
rect 35713 36867 35771 36873
rect 35894 36864 35900 36876
rect 35952 36864 35958 36916
rect 36170 36864 36176 36916
rect 36228 36904 36234 36916
rect 38105 36907 38163 36913
rect 38105 36904 38117 36907
rect 36228 36876 38117 36904
rect 36228 36864 36234 36876
rect 38105 36873 38117 36876
rect 38151 36873 38163 36907
rect 38105 36867 38163 36873
rect 22554 36796 22560 36848
rect 22612 36836 22618 36848
rect 22612 36808 37596 36836
rect 22612 36796 22618 36808
rect 7098 36728 7104 36780
rect 7156 36768 7162 36780
rect 15930 36768 15936 36780
rect 7156 36740 15936 36768
rect 7156 36728 7162 36740
rect 15930 36728 15936 36740
rect 15988 36728 15994 36780
rect 21545 36771 21603 36777
rect 21545 36737 21557 36771
rect 21591 36768 21603 36771
rect 21726 36768 21732 36780
rect 21591 36740 21732 36768
rect 21591 36737 21603 36740
rect 21545 36731 21603 36737
rect 21726 36728 21732 36740
rect 21784 36728 21790 36780
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 23937 36771 23995 36777
rect 23532 36740 23888 36768
rect 23532 36728 23538 36740
rect 1394 36700 1400 36712
rect 1355 36672 1400 36700
rect 1394 36660 1400 36672
rect 1452 36660 1458 36712
rect 21269 36703 21327 36709
rect 21269 36669 21281 36703
rect 21315 36700 21327 36703
rect 22462 36700 22468 36712
rect 21315 36672 22468 36700
rect 21315 36669 21327 36672
rect 21269 36663 21327 36669
rect 22462 36660 22468 36672
rect 22520 36660 22526 36712
rect 23566 36660 23572 36712
rect 23624 36700 23630 36712
rect 23661 36703 23719 36709
rect 23661 36700 23673 36703
rect 23624 36672 23673 36700
rect 23624 36660 23630 36672
rect 23661 36669 23673 36672
rect 23707 36669 23719 36703
rect 23661 36663 23719 36669
rect 23753 36703 23811 36709
rect 23753 36669 23765 36703
rect 23799 36669 23811 36703
rect 23860 36700 23888 36740
rect 23937 36737 23949 36771
rect 23983 36768 23995 36771
rect 24394 36768 24400 36780
rect 23983 36740 24400 36768
rect 23983 36737 23995 36740
rect 23937 36731 23995 36737
rect 24394 36728 24400 36740
rect 24452 36728 24458 36780
rect 25884 36740 26832 36768
rect 24029 36703 24087 36709
rect 24029 36700 24041 36703
rect 23860 36672 24041 36700
rect 23753 36663 23811 36669
rect 24029 36669 24041 36672
rect 24075 36669 24087 36703
rect 24029 36663 24087 36669
rect 20162 36632 20168 36644
rect 12406 36604 20168 36632
rect 8754 36524 8760 36576
rect 8812 36564 8818 36576
rect 12406 36564 12434 36604
rect 20162 36592 20168 36604
rect 20220 36592 20226 36644
rect 23198 36592 23204 36644
rect 23256 36632 23262 36644
rect 23768 36632 23796 36663
rect 25884 36632 25912 36740
rect 26234 36700 26240 36712
rect 26195 36672 26240 36700
rect 26234 36660 26240 36672
rect 26292 36660 26298 36712
rect 26510 36700 26516 36712
rect 26471 36672 26516 36700
rect 26510 36660 26516 36672
rect 26568 36660 26574 36712
rect 26602 36660 26608 36712
rect 26660 36709 26666 36712
rect 26660 36700 26668 36709
rect 26804 36700 26832 36740
rect 27982 36728 27988 36780
rect 28040 36768 28046 36780
rect 28445 36771 28503 36777
rect 28445 36768 28457 36771
rect 28040 36740 28457 36768
rect 28040 36728 28046 36740
rect 28445 36737 28457 36740
rect 28491 36737 28503 36771
rect 28445 36731 28503 36737
rect 28537 36771 28595 36777
rect 28537 36737 28549 36771
rect 28583 36768 28595 36771
rect 29914 36768 29920 36780
rect 28583 36740 29920 36768
rect 28583 36737 28595 36740
rect 28537 36731 28595 36737
rect 29914 36728 29920 36740
rect 29972 36728 29978 36780
rect 28353 36703 28411 36709
rect 28353 36700 28365 36703
rect 26660 36672 26705 36700
rect 26804 36672 28365 36700
rect 26660 36663 26668 36672
rect 28353 36669 28365 36672
rect 28399 36669 28411 36703
rect 28353 36663 28411 36669
rect 28629 36703 28687 36709
rect 28629 36669 28641 36703
rect 28675 36669 28687 36703
rect 28629 36663 28687 36669
rect 28813 36703 28871 36709
rect 28813 36669 28825 36703
rect 28859 36700 28871 36703
rect 29086 36700 29092 36712
rect 28859 36672 29092 36700
rect 28859 36669 28871 36672
rect 28813 36663 28871 36669
rect 26660 36660 26666 36663
rect 26418 36632 26424 36644
rect 23256 36604 23796 36632
rect 23860 36604 25912 36632
rect 26379 36604 26424 36632
rect 23256 36592 23262 36604
rect 8812 36536 12434 36564
rect 8812 36524 8818 36536
rect 22278 36524 22284 36576
rect 22336 36564 22342 36576
rect 22649 36567 22707 36573
rect 22649 36564 22661 36567
rect 22336 36536 22661 36564
rect 22336 36524 22342 36536
rect 22649 36533 22661 36536
rect 22695 36533 22707 36567
rect 22649 36527 22707 36533
rect 23290 36524 23296 36576
rect 23348 36564 23354 36576
rect 23860 36564 23888 36604
rect 26418 36592 26424 36604
rect 26476 36592 26482 36644
rect 27982 36592 27988 36644
rect 28040 36632 28046 36644
rect 28644 36632 28672 36663
rect 29086 36660 29092 36672
rect 29144 36700 29150 36712
rect 30006 36700 30012 36712
rect 29144 36672 30012 36700
rect 29144 36660 29150 36672
rect 30006 36660 30012 36672
rect 30064 36660 30070 36712
rect 35713 36703 35771 36709
rect 35713 36669 35725 36703
rect 35759 36700 35771 36703
rect 35897 36703 35955 36709
rect 35897 36700 35909 36703
rect 35759 36672 35909 36700
rect 35759 36669 35771 36672
rect 35713 36663 35771 36669
rect 35897 36669 35909 36672
rect 35943 36669 35955 36703
rect 35897 36663 35955 36669
rect 36078 36660 36084 36712
rect 36136 36700 36142 36712
rect 36354 36700 36360 36712
rect 36136 36672 36360 36700
rect 36136 36660 36142 36672
rect 36354 36660 36360 36672
rect 36412 36660 36418 36712
rect 36446 36660 36452 36712
rect 36504 36700 36510 36712
rect 36998 36709 37004 36712
rect 36541 36703 36599 36709
rect 36541 36700 36553 36703
rect 36504 36672 36553 36700
rect 36504 36660 36510 36672
rect 36541 36669 36553 36672
rect 36587 36669 36599 36703
rect 36541 36663 36599 36669
rect 36955 36703 37004 36709
rect 36955 36669 36967 36703
rect 37001 36669 37004 36703
rect 36955 36663 37004 36669
rect 36998 36660 37004 36663
rect 37056 36660 37062 36712
rect 37568 36709 37596 36808
rect 37553 36703 37611 36709
rect 37553 36669 37565 36703
rect 37599 36669 37611 36703
rect 37918 36700 37924 36712
rect 37879 36672 37924 36700
rect 37553 36663 37611 36669
rect 37918 36660 37924 36672
rect 37976 36660 37982 36712
rect 28040 36604 28672 36632
rect 28040 36592 28046 36604
rect 35618 36592 35624 36644
rect 35676 36632 35682 36644
rect 36725 36635 36783 36641
rect 36725 36632 36737 36635
rect 35676 36604 36737 36632
rect 35676 36592 35682 36604
rect 36725 36601 36737 36604
rect 36771 36601 36783 36635
rect 36725 36595 36783 36601
rect 36817 36635 36875 36641
rect 36817 36601 36829 36635
rect 36863 36632 36875 36635
rect 37366 36632 37372 36644
rect 36863 36604 37372 36632
rect 36863 36601 36875 36604
rect 36817 36595 36875 36601
rect 37366 36592 37372 36604
rect 37424 36632 37430 36644
rect 37734 36632 37740 36644
rect 37424 36604 37504 36632
rect 37695 36604 37740 36632
rect 37424 36592 37430 36604
rect 23348 36536 23888 36564
rect 23348 36524 23354 36536
rect 26326 36524 26332 36576
rect 26384 36564 26390 36576
rect 26694 36564 26700 36576
rect 26384 36536 26700 36564
rect 26384 36524 26390 36536
rect 26694 36524 26700 36536
rect 26752 36524 26758 36576
rect 27706 36524 27712 36576
rect 27764 36564 27770 36576
rect 28169 36567 28227 36573
rect 28169 36564 28181 36567
rect 27764 36536 28181 36564
rect 27764 36524 27770 36536
rect 28169 36533 28181 36536
rect 28215 36533 28227 36567
rect 35986 36564 35992 36576
rect 35947 36536 35992 36564
rect 28169 36527 28227 36533
rect 35986 36524 35992 36536
rect 36044 36524 36050 36576
rect 36078 36524 36084 36576
rect 36136 36564 36142 36576
rect 37093 36567 37151 36573
rect 37093 36564 37105 36567
rect 36136 36536 37105 36564
rect 36136 36524 36142 36536
rect 37093 36533 37105 36536
rect 37139 36533 37151 36567
rect 37476 36564 37504 36604
rect 37734 36592 37740 36604
rect 37792 36592 37798 36644
rect 37826 36592 37832 36644
rect 37884 36632 37890 36644
rect 37884 36604 37929 36632
rect 37884 36592 37890 36604
rect 37844 36564 37872 36592
rect 37476 36536 37872 36564
rect 37093 36527 37151 36533
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 1581 36363 1639 36369
rect 1581 36329 1593 36363
rect 1627 36360 1639 36363
rect 1670 36360 1676 36372
rect 1627 36332 1676 36360
rect 1627 36329 1639 36332
rect 1581 36323 1639 36329
rect 1670 36320 1676 36332
rect 1728 36320 1734 36372
rect 1762 36320 1768 36372
rect 1820 36360 1826 36372
rect 26602 36360 26608 36372
rect 1820 36332 26608 36360
rect 1820 36320 1826 36332
rect 26602 36320 26608 36332
rect 26660 36320 26666 36372
rect 27154 36320 27160 36372
rect 27212 36360 27218 36372
rect 33042 36360 33048 36372
rect 27212 36332 33048 36360
rect 27212 36320 27218 36332
rect 33042 36320 33048 36332
rect 33100 36320 33106 36372
rect 34790 36360 34796 36372
rect 34751 36332 34796 36360
rect 34790 36320 34796 36332
rect 34848 36320 34854 36372
rect 35253 36363 35311 36369
rect 35253 36329 35265 36363
rect 35299 36360 35311 36363
rect 35894 36360 35900 36372
rect 35299 36332 35900 36360
rect 35299 36329 35311 36332
rect 35253 36323 35311 36329
rect 35894 36320 35900 36332
rect 35952 36320 35958 36372
rect 36814 36360 36820 36372
rect 36060 36332 36820 36360
rect 2038 36252 2044 36304
rect 2096 36292 2102 36304
rect 2096 36264 26653 36292
rect 2096 36252 2102 36264
rect 1394 36224 1400 36236
rect 1355 36196 1400 36224
rect 1394 36184 1400 36196
rect 1452 36184 1458 36236
rect 21450 36224 21456 36236
rect 21363 36196 21456 36224
rect 21450 36184 21456 36196
rect 21508 36184 21514 36236
rect 21545 36227 21603 36233
rect 21545 36193 21557 36227
rect 21591 36224 21603 36227
rect 22830 36224 22836 36236
rect 21591 36196 22836 36224
rect 21591 36193 21603 36196
rect 21545 36187 21603 36193
rect 22830 36184 22836 36196
rect 22888 36184 22894 36236
rect 23376 36227 23434 36233
rect 23376 36193 23388 36227
rect 23422 36224 23434 36227
rect 24210 36224 24216 36236
rect 23422 36196 24216 36224
rect 23422 36193 23434 36196
rect 23376 36187 23434 36193
rect 24210 36184 24216 36196
rect 24268 36184 24274 36236
rect 26237 36227 26295 36233
rect 26237 36193 26249 36227
rect 26283 36193 26295 36227
rect 26237 36187 26295 36193
rect 21468 36156 21496 36184
rect 22278 36156 22284 36168
rect 21468 36128 22284 36156
rect 22278 36116 22284 36128
rect 22336 36116 22342 36168
rect 22462 36116 22468 36168
rect 22520 36156 22526 36168
rect 23109 36159 23167 36165
rect 23109 36156 23121 36159
rect 22520 36128 23121 36156
rect 22520 36116 22526 36128
rect 23109 36125 23121 36128
rect 23155 36125 23167 36159
rect 26252 36156 26280 36187
rect 26326 36184 26332 36236
rect 26384 36233 26390 36236
rect 26384 36227 26433 36233
rect 26384 36193 26387 36227
rect 26421 36193 26433 36227
rect 26510 36224 26516 36236
rect 26471 36196 26516 36224
rect 26384 36187 26433 36193
rect 26384 36184 26390 36187
rect 26510 36184 26516 36196
rect 26568 36184 26574 36236
rect 26625 36233 26653 36264
rect 27338 36252 27344 36304
rect 27396 36292 27402 36304
rect 31846 36292 31852 36304
rect 27396 36264 31852 36292
rect 27396 36252 27402 36264
rect 31846 36252 31852 36264
rect 31904 36252 31910 36304
rect 26610 36227 26668 36233
rect 26610 36193 26622 36227
rect 26656 36193 26668 36227
rect 26610 36187 26668 36193
rect 26806 36227 26864 36233
rect 26806 36193 26818 36227
rect 26852 36224 26864 36227
rect 26970 36224 26976 36236
rect 26852 36196 26976 36224
rect 26852 36193 26864 36196
rect 26806 36187 26864 36193
rect 26970 36184 26976 36196
rect 27028 36184 27034 36236
rect 34609 36227 34667 36233
rect 34609 36193 34621 36227
rect 34655 36224 34667 36227
rect 34790 36224 34796 36236
rect 34655 36196 34796 36224
rect 34655 36193 34667 36196
rect 34609 36187 34667 36193
rect 34790 36184 34796 36196
rect 34848 36184 34854 36236
rect 35434 36224 35440 36236
rect 35395 36196 35440 36224
rect 35434 36184 35440 36196
rect 35492 36184 35498 36236
rect 35894 36224 35900 36236
rect 35855 36196 35900 36224
rect 35894 36184 35900 36196
rect 35952 36184 35958 36236
rect 36060 36233 36088 36332
rect 36814 36320 36820 36332
rect 36872 36320 36878 36372
rect 38930 36360 38936 36372
rect 37292 36332 38936 36360
rect 36265 36295 36323 36301
rect 36265 36261 36277 36295
rect 36311 36292 36323 36295
rect 37292 36292 37320 36332
rect 38930 36320 38936 36332
rect 38988 36320 38994 36372
rect 36311 36264 37320 36292
rect 37369 36295 37427 36301
rect 36311 36261 36323 36264
rect 36265 36255 36323 36261
rect 37369 36261 37381 36295
rect 37415 36292 37427 36295
rect 37458 36292 37464 36304
rect 37415 36264 37464 36292
rect 37415 36261 37427 36264
rect 37369 36255 37427 36261
rect 37458 36252 37464 36264
rect 37516 36252 37522 36304
rect 36045 36227 36103 36233
rect 36045 36193 36057 36227
rect 36091 36193 36103 36227
rect 36045 36187 36103 36193
rect 36173 36227 36231 36233
rect 36173 36193 36185 36227
rect 36219 36193 36231 36227
rect 36173 36187 36231 36193
rect 27338 36156 27344 36168
rect 26252 36128 27344 36156
rect 23109 36119 23167 36125
rect 27338 36116 27344 36128
rect 27396 36116 27402 36168
rect 35802 36116 35808 36168
rect 35860 36156 35866 36168
rect 36188 36156 36216 36187
rect 36354 36184 36360 36236
rect 36412 36233 36418 36236
rect 36412 36224 36420 36233
rect 37185 36227 37243 36233
rect 36412 36196 36457 36224
rect 36412 36187 36420 36196
rect 37185 36193 37197 36227
rect 37231 36193 37243 36227
rect 37185 36187 37243 36193
rect 36412 36184 36418 36187
rect 35860 36128 36216 36156
rect 35860 36116 35866 36128
rect 24670 36048 24676 36100
rect 24728 36088 24734 36100
rect 36541 36091 36599 36097
rect 36541 36088 36553 36091
rect 24728 36060 36553 36088
rect 24728 36048 24734 36060
rect 36541 36057 36553 36060
rect 36587 36057 36599 36091
rect 36541 36051 36599 36057
rect 23382 35980 23388 36032
rect 23440 36020 23446 36032
rect 24394 36020 24400 36032
rect 23440 35992 24400 36020
rect 23440 35980 23446 35992
rect 24394 35980 24400 35992
rect 24452 36020 24458 36032
rect 24489 36023 24547 36029
rect 24489 36020 24501 36023
rect 24452 35992 24501 36020
rect 24452 35980 24458 35992
rect 24489 35989 24501 35992
rect 24535 35989 24547 36023
rect 24489 35983 24547 35989
rect 27522 35980 27528 36032
rect 27580 36020 27586 36032
rect 27798 36020 27804 36032
rect 27580 35992 27804 36020
rect 27580 35980 27586 35992
rect 27798 35980 27804 35992
rect 27856 35980 27862 36032
rect 30282 35980 30288 36032
rect 30340 36020 30346 36032
rect 34514 36020 34520 36032
rect 30340 35992 34520 36020
rect 30340 35980 30346 35992
rect 34514 35980 34520 35992
rect 34572 35980 34578 36032
rect 34606 35980 34612 36032
rect 34664 36020 34670 36032
rect 37200 36020 37228 36187
rect 34664 35992 37228 36020
rect 34664 35980 34670 35992
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 22741 35819 22799 35825
rect 22741 35785 22753 35819
rect 22787 35816 22799 35819
rect 23198 35816 23204 35828
rect 22787 35788 23204 35816
rect 22787 35785 22799 35788
rect 22741 35779 22799 35785
rect 23198 35776 23204 35788
rect 23256 35776 23262 35828
rect 26326 35776 26332 35828
rect 26384 35816 26390 35828
rect 27154 35816 27160 35828
rect 26384 35788 27160 35816
rect 26384 35776 26390 35788
rect 27154 35776 27160 35788
rect 27212 35776 27218 35828
rect 27798 35776 27804 35828
rect 27856 35816 27862 35828
rect 28718 35816 28724 35828
rect 27856 35788 28724 35816
rect 27856 35776 27862 35788
rect 28718 35776 28724 35788
rect 28776 35776 28782 35828
rect 33318 35776 33324 35828
rect 33376 35816 33382 35828
rect 33962 35816 33968 35828
rect 33376 35788 33968 35816
rect 33376 35776 33382 35788
rect 33962 35776 33968 35788
rect 34020 35776 34026 35828
rect 34609 35819 34667 35825
rect 34609 35785 34621 35819
rect 34655 35816 34667 35819
rect 35250 35816 35256 35828
rect 34655 35788 35256 35816
rect 34655 35785 34667 35788
rect 34609 35779 34667 35785
rect 35250 35776 35256 35788
rect 35308 35776 35314 35828
rect 35894 35776 35900 35828
rect 35952 35816 35958 35828
rect 37550 35816 37556 35828
rect 35952 35788 37556 35816
rect 35952 35776 35958 35788
rect 37550 35776 37556 35788
rect 37608 35776 37614 35828
rect 7834 35708 7840 35760
rect 7892 35748 7898 35760
rect 14826 35748 14832 35760
rect 7892 35720 14832 35748
rect 7892 35708 7898 35720
rect 14826 35708 14832 35720
rect 14884 35708 14890 35760
rect 20530 35708 20536 35760
rect 20588 35748 20594 35760
rect 20588 35720 37412 35748
rect 20588 35708 20594 35720
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 22925 35683 22983 35689
rect 22925 35680 22937 35683
rect 22888 35652 22937 35680
rect 22888 35640 22894 35652
rect 22925 35649 22937 35652
rect 22971 35649 22983 35683
rect 22925 35643 22983 35649
rect 26786 35640 26792 35692
rect 26844 35680 26850 35692
rect 31938 35680 31944 35692
rect 26844 35652 31944 35680
rect 26844 35640 26850 35652
rect 31938 35640 31944 35652
rect 31996 35640 32002 35692
rect 36446 35680 36452 35692
rect 35544 35652 36452 35680
rect 35544 35624 35572 35652
rect 22649 35615 22707 35621
rect 22649 35581 22661 35615
rect 22695 35581 22707 35615
rect 22649 35575 22707 35581
rect 8386 35504 8392 35556
rect 8444 35544 8450 35556
rect 15746 35544 15752 35556
rect 8444 35516 15752 35544
rect 8444 35504 8450 35516
rect 15746 35504 15752 35516
rect 15804 35504 15810 35556
rect 22664 35476 22692 35575
rect 23566 35572 23572 35624
rect 23624 35612 23630 35624
rect 23937 35615 23995 35621
rect 23937 35612 23949 35615
rect 23624 35584 23949 35612
rect 23624 35572 23630 35584
rect 23937 35581 23949 35584
rect 23983 35581 23995 35615
rect 23937 35575 23995 35581
rect 26234 35572 26240 35624
rect 26292 35612 26298 35624
rect 33226 35612 33232 35624
rect 26292 35584 33232 35612
rect 26292 35572 26298 35584
rect 33226 35572 33232 35584
rect 33284 35572 33290 35624
rect 34790 35612 34796 35624
rect 34751 35584 34796 35612
rect 34790 35572 34796 35584
rect 34848 35572 34854 35624
rect 35526 35572 35532 35624
rect 35584 35572 35590 35624
rect 35894 35612 35900 35624
rect 35855 35584 35900 35612
rect 35894 35572 35900 35584
rect 35952 35572 35958 35624
rect 36280 35621 36308 35652
rect 36446 35640 36452 35652
rect 36504 35640 36510 35692
rect 36814 35640 36820 35692
rect 36872 35640 36878 35692
rect 37274 35680 37280 35692
rect 37108 35652 37280 35680
rect 35990 35615 36048 35621
rect 35990 35581 36002 35615
rect 36036 35581 36048 35615
rect 35990 35575 36048 35581
rect 36265 35615 36323 35621
rect 36265 35581 36277 35615
rect 36311 35581 36323 35615
rect 36265 35575 36323 35581
rect 22925 35547 22983 35553
rect 22925 35513 22937 35547
rect 22971 35544 22983 35547
rect 24302 35544 24308 35556
rect 22971 35516 24308 35544
rect 22971 35513 22983 35516
rect 22925 35507 22983 35513
rect 24302 35504 24308 35516
rect 24360 35504 24366 35556
rect 26970 35504 26976 35556
rect 27028 35544 27034 35556
rect 33318 35544 33324 35556
rect 27028 35516 33324 35544
rect 27028 35504 27034 35516
rect 33318 35504 33324 35516
rect 33376 35504 33382 35556
rect 35342 35504 35348 35556
rect 35400 35544 35406 35556
rect 36004 35544 36032 35575
rect 36354 35572 36360 35624
rect 36412 35621 36418 35624
rect 36412 35612 36420 35621
rect 36832 35612 36860 35640
rect 37108 35621 37136 35652
rect 37274 35640 37280 35652
rect 37332 35640 37338 35692
rect 36412 35584 36457 35612
rect 36510 35584 36860 35612
rect 37093 35615 37151 35621
rect 36412 35575 36420 35584
rect 36412 35572 36418 35575
rect 35400 35516 36032 35544
rect 36173 35547 36231 35553
rect 35400 35504 35406 35516
rect 36173 35513 36185 35547
rect 36219 35544 36231 35547
rect 36510 35544 36538 35584
rect 36219 35516 36538 35544
rect 36219 35513 36231 35516
rect 36173 35507 36231 35513
rect 23474 35476 23480 35488
rect 22664 35448 23480 35476
rect 23474 35436 23480 35448
rect 23532 35476 23538 35488
rect 24029 35479 24087 35485
rect 24029 35476 24041 35479
rect 23532 35448 24041 35476
rect 23532 35436 23538 35448
rect 24029 35445 24041 35448
rect 24075 35445 24087 35479
rect 24029 35439 24087 35445
rect 26602 35436 26608 35488
rect 26660 35476 26666 35488
rect 31570 35476 31576 35488
rect 26660 35448 31576 35476
rect 26660 35436 26666 35448
rect 31570 35436 31576 35448
rect 31628 35436 31634 35488
rect 33042 35436 33048 35488
rect 33100 35476 33106 35488
rect 36541 35479 36599 35485
rect 36541 35476 36553 35479
rect 33100 35448 36553 35476
rect 33100 35436 33106 35448
rect 36541 35445 36553 35448
rect 36587 35445 36599 35479
rect 36740 35476 36768 35584
rect 37093 35581 37105 35615
rect 37139 35581 37151 35615
rect 37093 35575 37151 35581
rect 37186 35615 37244 35621
rect 37186 35581 37198 35615
rect 37232 35581 37244 35615
rect 37384 35612 37412 35720
rect 37558 35615 37616 35621
rect 37558 35612 37570 35615
rect 37384 35584 37570 35612
rect 37186 35575 37244 35581
rect 37558 35581 37570 35584
rect 37604 35581 37616 35615
rect 37558 35575 37616 35581
rect 36814 35504 36820 35556
rect 36872 35544 36878 35556
rect 37200 35544 37228 35575
rect 36872 35516 37228 35544
rect 37369 35547 37427 35553
rect 36872 35504 36878 35516
rect 37369 35513 37381 35547
rect 37415 35513 37427 35547
rect 37369 35507 37427 35513
rect 37384 35476 37412 35507
rect 37458 35504 37464 35556
rect 37516 35544 37522 35556
rect 37516 35516 37561 35544
rect 37516 35504 37522 35516
rect 36740 35448 37412 35476
rect 37737 35479 37795 35485
rect 36541 35439 36599 35445
rect 37737 35445 37749 35479
rect 37783 35476 37795 35479
rect 38746 35476 38752 35488
rect 37783 35448 38752 35476
rect 37783 35445 37795 35448
rect 37737 35439 37795 35445
rect 38746 35436 38752 35448
rect 38804 35436 38810 35488
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 2498 35272 2504 35284
rect 1627 35244 2504 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 2498 35232 2504 35244
rect 2556 35232 2562 35284
rect 2608 35244 12848 35272
rect 2406 35164 2412 35216
rect 2464 35204 2470 35216
rect 2608 35204 2636 35244
rect 2464 35176 2636 35204
rect 2464 35164 2470 35176
rect 4798 35164 4804 35216
rect 4856 35204 4862 35216
rect 12820 35204 12848 35244
rect 23198 35232 23204 35284
rect 23256 35272 23262 35284
rect 23477 35275 23535 35281
rect 23477 35272 23489 35275
rect 23256 35244 23489 35272
rect 23256 35232 23262 35244
rect 23477 35241 23489 35244
rect 23523 35241 23535 35275
rect 23477 35235 23535 35241
rect 26234 35232 26240 35284
rect 26292 35272 26298 35284
rect 28626 35272 28632 35284
rect 26292 35244 28632 35272
rect 26292 35232 26298 35244
rect 28626 35232 28632 35244
rect 28684 35232 28690 35284
rect 31386 35232 31392 35284
rect 31444 35272 31450 35284
rect 36725 35275 36783 35281
rect 36725 35272 36737 35275
rect 31444 35244 36737 35272
rect 31444 35232 31450 35244
rect 36725 35241 36737 35244
rect 36771 35241 36783 35275
rect 36725 35235 36783 35241
rect 23106 35204 23112 35216
rect 4856 35176 12434 35204
rect 12820 35176 23112 35204
rect 4856 35164 4862 35176
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 12406 35136 12434 35176
rect 23106 35164 23112 35176
rect 23164 35164 23170 35216
rect 26896 35176 31754 35204
rect 18598 35136 18604 35148
rect 12406 35108 18604 35136
rect 18598 35096 18604 35108
rect 18656 35096 18662 35148
rect 22462 35096 22468 35148
rect 22520 35136 22526 35148
rect 23382 35136 23388 35148
rect 22520 35108 23388 35136
rect 22520 35096 22526 35108
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 26896 35068 26924 35176
rect 27522 35096 27528 35148
rect 27580 35136 27586 35148
rect 27801 35139 27859 35145
rect 27801 35136 27813 35139
rect 27580 35108 27813 35136
rect 27580 35096 27614 35108
rect 27801 35105 27813 35108
rect 27847 35105 27859 35139
rect 27801 35099 27859 35105
rect 28068 35139 28126 35145
rect 28068 35105 28080 35139
rect 28114 35136 28126 35139
rect 28442 35136 28448 35148
rect 28114 35108 28448 35136
rect 28114 35105 28126 35108
rect 28068 35099 28126 35105
rect 28442 35096 28448 35108
rect 28500 35096 28506 35148
rect 31726 35136 31754 35176
rect 34606 35164 34612 35216
rect 34664 35204 34670 35216
rect 35437 35207 35495 35213
rect 35437 35204 35449 35207
rect 34664 35176 35449 35204
rect 34664 35164 34670 35176
rect 35437 35173 35449 35176
rect 35483 35204 35495 35207
rect 35894 35204 35900 35216
rect 35483 35176 35900 35204
rect 35483 35173 35495 35176
rect 35437 35167 35495 35173
rect 35894 35164 35900 35176
rect 35952 35164 35958 35216
rect 36359 35213 36365 35216
rect 36357 35204 36365 35213
rect 36320 35176 36365 35204
rect 36357 35167 36365 35176
rect 36359 35164 36365 35167
rect 36417 35164 36423 35216
rect 34514 35136 34520 35148
rect 31726 35108 34520 35136
rect 34514 35096 34520 35108
rect 34572 35096 34578 35148
rect 35618 35096 35624 35148
rect 35676 35136 35682 35148
rect 36262 35145 36268 35148
rect 36081 35139 36139 35145
rect 36081 35136 36093 35139
rect 35676 35108 36093 35136
rect 35676 35096 35682 35108
rect 36081 35105 36093 35108
rect 36127 35105 36139 35139
rect 36081 35099 36139 35105
rect 36229 35139 36268 35145
rect 36229 35105 36241 35139
rect 36229 35099 36268 35105
rect 36262 35096 36268 35099
rect 36320 35096 36326 35148
rect 36446 35136 36452 35148
rect 36407 35108 36452 35136
rect 36446 35096 36452 35108
rect 36504 35096 36510 35148
rect 36546 35139 36604 35145
rect 36546 35105 36558 35139
rect 36592 35105 36604 35139
rect 36546 35099 36604 35105
rect 37185 35139 37243 35145
rect 37185 35105 37197 35139
rect 37231 35136 37243 35139
rect 37274 35136 37280 35148
rect 37231 35108 37280 35136
rect 37231 35105 37243 35108
rect 37185 35099 37243 35105
rect 20956 35040 26924 35068
rect 20956 35028 20962 35040
rect 22066 34972 23612 35000
rect 18506 34892 18512 34944
rect 18564 34932 18570 34944
rect 22066 34932 22094 34972
rect 18564 34904 22094 34932
rect 23584 34932 23612 34972
rect 25866 34960 25872 35012
rect 25924 35000 25930 35012
rect 27586 35000 27614 35096
rect 29914 35028 29920 35080
rect 29972 35068 29978 35080
rect 30650 35068 30656 35080
rect 29972 35040 30656 35068
rect 29972 35028 29978 35040
rect 30650 35028 30656 35040
rect 30708 35028 30714 35080
rect 36561 35000 36589 35099
rect 37274 35096 37280 35108
rect 37332 35096 37338 35148
rect 25924 34972 27614 35000
rect 28736 34972 36589 35000
rect 25924 34960 25930 34972
rect 28736 34932 28764 34972
rect 23584 34904 28764 34932
rect 29181 34935 29239 34941
rect 18564 34892 18570 34904
rect 29181 34901 29193 34935
rect 29227 34932 29239 34935
rect 29270 34932 29276 34944
rect 29227 34904 29276 34932
rect 29227 34901 29239 34904
rect 29181 34895 29239 34901
rect 29270 34892 29276 34904
rect 29328 34892 29334 34944
rect 35526 34932 35532 34944
rect 35487 34904 35532 34932
rect 35526 34892 35532 34904
rect 35584 34892 35590 34944
rect 35618 34892 35624 34944
rect 35676 34932 35682 34944
rect 36630 34932 36636 34944
rect 35676 34904 36636 34932
rect 35676 34892 35682 34904
rect 36630 34892 36636 34904
rect 36688 34892 36694 34944
rect 37369 34935 37427 34941
rect 37369 34901 37381 34935
rect 37415 34932 37427 34935
rect 37826 34932 37832 34944
rect 37415 34904 37832 34932
rect 37415 34901 37427 34904
rect 37369 34895 37427 34901
rect 37826 34892 37832 34904
rect 37884 34892 37890 34944
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 1762 34728 1768 34740
rect 1627 34700 1768 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 1762 34688 1768 34700
rect 1820 34688 1826 34740
rect 22066 34700 36272 34728
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 22066 34592 22094 34700
rect 22554 34620 22560 34672
rect 22612 34660 22618 34672
rect 24210 34660 24216 34672
rect 22612 34632 24216 34660
rect 22612 34620 22618 34632
rect 24210 34620 24216 34632
rect 24268 34660 24274 34672
rect 25225 34663 25283 34669
rect 25225 34660 25237 34663
rect 24268 34632 25237 34660
rect 24268 34620 24274 34632
rect 25225 34629 25237 34632
rect 25271 34629 25283 34663
rect 25225 34623 25283 34629
rect 20680 34564 22094 34592
rect 25240 34592 25268 34623
rect 27982 34620 27988 34672
rect 28040 34660 28046 34672
rect 28077 34663 28135 34669
rect 28077 34660 28089 34663
rect 28040 34632 28089 34660
rect 28040 34620 28046 34632
rect 28077 34629 28089 34632
rect 28123 34629 28135 34663
rect 28077 34623 28135 34629
rect 28905 34663 28963 34669
rect 28905 34629 28917 34663
rect 28951 34660 28963 34663
rect 28994 34660 29000 34672
rect 28951 34632 29000 34660
rect 28951 34629 28963 34632
rect 28905 34623 28963 34629
rect 28994 34620 29000 34632
rect 29052 34620 29058 34672
rect 29822 34620 29828 34672
rect 29880 34660 29886 34672
rect 34793 34663 34851 34669
rect 34793 34660 34805 34663
rect 29880 34632 34805 34660
rect 29880 34620 29886 34632
rect 34793 34629 34805 34632
rect 34839 34629 34851 34663
rect 36244 34660 36272 34700
rect 36244 34632 36584 34660
rect 34793 34623 34851 34629
rect 26697 34595 26755 34601
rect 26697 34592 26709 34595
rect 25240 34564 26709 34592
rect 20680 34552 20686 34564
rect 26697 34561 26709 34564
rect 26743 34561 26755 34595
rect 26697 34555 26755 34561
rect 1394 34524 1400 34536
rect 1355 34496 1400 34524
rect 1394 34484 1400 34496
rect 1452 34484 1458 34536
rect 10686 34484 10692 34536
rect 10744 34524 10750 34536
rect 11790 34524 11796 34536
rect 10744 34496 11796 34524
rect 10744 34484 10750 34496
rect 11790 34484 11796 34496
rect 11848 34484 11854 34536
rect 11882 34484 11888 34536
rect 11940 34524 11946 34536
rect 17770 34524 17776 34536
rect 11940 34496 17776 34524
rect 11940 34484 11946 34496
rect 17770 34484 17776 34496
rect 17828 34484 17834 34536
rect 22278 34484 22284 34536
rect 22336 34524 22342 34536
rect 22554 34524 22560 34536
rect 22336 34496 22560 34524
rect 22336 34484 22342 34496
rect 22554 34484 22560 34496
rect 22612 34484 22618 34536
rect 25409 34527 25467 34533
rect 25409 34493 25421 34527
rect 25455 34524 25467 34527
rect 26237 34527 26295 34533
rect 26237 34524 26249 34527
rect 25455 34496 26249 34524
rect 25455 34493 25467 34496
rect 25409 34487 25467 34493
rect 26237 34493 26249 34496
rect 26283 34524 26295 34527
rect 26510 34524 26516 34536
rect 26283 34496 26516 34524
rect 26283 34493 26295 34496
rect 26237 34487 26295 34493
rect 26510 34484 26516 34496
rect 26568 34484 26574 34536
rect 25866 34348 25872 34400
rect 25924 34388 25930 34400
rect 26053 34391 26111 34397
rect 26053 34388 26065 34391
rect 25924 34360 26065 34388
rect 25924 34348 25930 34360
rect 26053 34357 26065 34360
rect 26099 34357 26111 34391
rect 26712 34388 26740 34555
rect 28718 34552 28724 34604
rect 28776 34592 28782 34604
rect 29089 34595 29147 34601
rect 29089 34592 29101 34595
rect 28776 34564 29101 34592
rect 28776 34552 28782 34564
rect 29089 34561 29101 34564
rect 29135 34561 29147 34595
rect 29454 34592 29460 34604
rect 29089 34555 29147 34561
rect 29196 34564 29460 34592
rect 26964 34527 27022 34533
rect 26964 34493 26976 34527
rect 27010 34524 27022 34527
rect 27706 34524 27712 34536
rect 27010 34496 27712 34524
rect 27010 34493 27022 34496
rect 26964 34487 27022 34493
rect 27706 34484 27712 34496
rect 27764 34484 27770 34536
rect 28813 34527 28871 34533
rect 28813 34493 28825 34527
rect 28859 34493 28871 34527
rect 28813 34487 28871 34493
rect 28997 34527 29055 34533
rect 28997 34493 29009 34527
rect 29043 34524 29055 34527
rect 29196 34524 29224 34564
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 36556 34592 36584 34632
rect 36630 34620 36636 34672
rect 36688 34660 36694 34672
rect 37550 34660 37556 34672
rect 36688 34632 37556 34660
rect 36688 34620 36694 34632
rect 37550 34620 37556 34632
rect 37608 34620 37614 34672
rect 36556 34564 36589 34592
rect 29043 34496 29224 34524
rect 29273 34527 29331 34533
rect 29043 34493 29055 34496
rect 28997 34487 29055 34493
rect 29273 34493 29285 34527
rect 29319 34493 29331 34527
rect 34606 34524 34612 34536
rect 34567 34496 34612 34524
rect 29273 34487 29331 34493
rect 28828 34400 28856 34487
rect 29086 34416 29092 34468
rect 29144 34456 29150 34468
rect 29288 34456 29316 34487
rect 34606 34484 34612 34496
rect 34664 34484 34670 34536
rect 35526 34484 35532 34536
rect 35584 34524 35590 34536
rect 36081 34527 36139 34533
rect 36081 34524 36093 34527
rect 35584 34496 36093 34524
rect 35584 34484 35590 34496
rect 36081 34493 36093 34496
rect 36127 34493 36139 34527
rect 36081 34487 36139 34493
rect 36174 34527 36232 34533
rect 36174 34493 36186 34527
rect 36220 34493 36232 34527
rect 36174 34487 36232 34493
rect 29144 34428 29316 34456
rect 29144 34416 29150 34428
rect 35618 34416 35624 34468
rect 35676 34456 35682 34468
rect 36189 34456 36217 34487
rect 36354 34484 36360 34536
rect 36412 34524 36418 34536
rect 36561 34533 36589 34564
rect 36546 34527 36604 34533
rect 36412 34496 36457 34524
rect 36412 34484 36418 34496
rect 36546 34493 36558 34527
rect 36592 34493 36604 34527
rect 36546 34487 36604 34493
rect 37553 34527 37611 34533
rect 37553 34493 37565 34527
rect 37599 34524 37611 34527
rect 37642 34524 37648 34536
rect 37599 34496 37648 34524
rect 37599 34493 37611 34496
rect 37553 34487 37611 34493
rect 37642 34484 37648 34496
rect 37700 34484 37706 34536
rect 37826 34524 37832 34536
rect 37787 34496 37832 34524
rect 37826 34484 37832 34496
rect 37884 34484 37890 34536
rect 37921 34527 37979 34533
rect 37921 34493 37933 34527
rect 37967 34524 37979 34527
rect 38562 34524 38568 34536
rect 37967 34496 38568 34524
rect 37967 34493 37979 34496
rect 37921 34487 37979 34493
rect 38562 34484 38568 34496
rect 38620 34484 38626 34536
rect 35676 34428 36217 34456
rect 35676 34416 35682 34428
rect 36447 34416 36453 34468
rect 36505 34456 36511 34468
rect 37734 34456 37740 34468
rect 36505 34428 36549 34456
rect 37695 34428 37740 34456
rect 36505 34416 36511 34428
rect 37734 34416 37740 34428
rect 37792 34416 37798 34468
rect 27706 34388 27712 34400
rect 26712 34360 27712 34388
rect 26053 34351 26111 34357
rect 27706 34348 27712 34360
rect 27764 34348 27770 34400
rect 28626 34388 28632 34400
rect 28587 34360 28632 34388
rect 28626 34348 28632 34360
rect 28684 34348 28690 34400
rect 28810 34348 28816 34400
rect 28868 34348 28874 34400
rect 36722 34388 36728 34400
rect 36683 34360 36728 34388
rect 36722 34348 36728 34360
rect 36780 34348 36786 34400
rect 38102 34388 38108 34400
rect 38063 34360 38108 34388
rect 38102 34348 38108 34360
rect 38160 34348 38166 34400
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 26145 34187 26203 34193
rect 26145 34153 26157 34187
rect 26191 34184 26203 34187
rect 28442 34184 28448 34196
rect 26191 34156 28448 34184
rect 26191 34153 26203 34156
rect 26145 34147 26203 34153
rect 28442 34144 28448 34156
rect 28500 34144 28506 34196
rect 28902 34144 28908 34196
rect 28960 34184 28966 34196
rect 29181 34187 29239 34193
rect 29181 34184 29193 34187
rect 28960 34156 29193 34184
rect 28960 34144 28966 34156
rect 29181 34153 29193 34156
rect 29227 34153 29239 34187
rect 29181 34147 29239 34153
rect 29917 34187 29975 34193
rect 29917 34153 29929 34187
rect 29963 34184 29975 34187
rect 30006 34184 30012 34196
rect 29963 34156 30012 34184
rect 29963 34153 29975 34156
rect 29917 34147 29975 34153
rect 30006 34144 30012 34156
rect 30064 34144 30070 34196
rect 30742 34144 30748 34196
rect 30800 34184 30806 34196
rect 36722 34184 36728 34196
rect 30800 34156 36728 34184
rect 30800 34144 30806 34156
rect 36722 34144 36728 34156
rect 36780 34144 36786 34196
rect 37182 34184 37188 34196
rect 37143 34156 37188 34184
rect 37182 34144 37188 34156
rect 37240 34144 37246 34196
rect 18322 34076 18328 34128
rect 18380 34116 18386 34128
rect 35526 34116 35532 34128
rect 18380 34088 35532 34116
rect 18380 34076 18386 34088
rect 35526 34076 35532 34088
rect 35584 34076 35590 34128
rect 35894 34076 35900 34128
rect 35952 34116 35958 34128
rect 36354 34116 36360 34128
rect 35952 34088 36217 34116
rect 36315 34088 36360 34116
rect 35952 34076 35958 34088
rect 25406 34048 25412 34060
rect 25367 34020 25412 34048
rect 25406 34008 25412 34020
rect 25464 34008 25470 34060
rect 26421 34051 26479 34057
rect 26421 34017 26433 34051
rect 26467 34048 26479 34051
rect 26786 34048 26792 34060
rect 26467 34020 26792 34048
rect 26467 34017 26479 34020
rect 26421 34011 26479 34017
rect 26786 34008 26792 34020
rect 26844 34008 26850 34060
rect 26881 34051 26939 34057
rect 26881 34017 26893 34051
rect 26927 34048 26939 34051
rect 26927 34020 27614 34048
rect 26927 34017 26939 34020
rect 26881 34011 26939 34017
rect 23106 33940 23112 33992
rect 23164 33980 23170 33992
rect 24670 33980 24676 33992
rect 23164 33952 24676 33980
rect 23164 33940 23170 33952
rect 24670 33940 24676 33952
rect 24728 33940 24734 33992
rect 26602 33980 26608 33992
rect 26563 33952 26608 33980
rect 26602 33940 26608 33952
rect 26660 33940 26666 33992
rect 26694 33940 26700 33992
rect 26752 33980 26758 33992
rect 26752 33952 26797 33980
rect 26752 33940 26758 33952
rect 7834 33872 7840 33924
rect 7892 33912 7898 33924
rect 18414 33912 18420 33924
rect 7892 33884 18420 33912
rect 7892 33872 7898 33884
rect 18414 33872 18420 33884
rect 18472 33872 18478 33924
rect 26513 33915 26571 33921
rect 26513 33881 26525 33915
rect 26559 33912 26571 33915
rect 27062 33912 27068 33924
rect 26559 33884 27068 33912
rect 26559 33881 26571 33884
rect 26513 33875 26571 33881
rect 27062 33872 27068 33884
rect 27120 33872 27126 33924
rect 2130 33804 2136 33856
rect 2188 33844 2194 33856
rect 18046 33844 18052 33856
rect 2188 33816 18052 33844
rect 2188 33804 2194 33816
rect 18046 33804 18052 33816
rect 18104 33804 18110 33856
rect 24946 33804 24952 33856
rect 25004 33844 25010 33856
rect 25593 33847 25651 33853
rect 25593 33844 25605 33847
rect 25004 33816 25605 33844
rect 25004 33804 25010 33816
rect 25593 33813 25605 33816
rect 25639 33844 25651 33847
rect 26145 33847 26203 33853
rect 26145 33844 26157 33847
rect 25639 33816 26157 33844
rect 25639 33813 25651 33816
rect 25593 33807 25651 33813
rect 26145 33813 26157 33816
rect 26191 33813 26203 33847
rect 26145 33807 26203 33813
rect 26237 33847 26295 33853
rect 26237 33813 26249 33847
rect 26283 33844 26295 33847
rect 26602 33844 26608 33856
rect 26283 33816 26608 33844
rect 26283 33813 26295 33816
rect 26237 33807 26295 33813
rect 26602 33804 26608 33816
rect 26660 33804 26666 33856
rect 27586 33844 27614 34020
rect 27706 34008 27712 34060
rect 27764 34048 27770 34060
rect 28074 34057 28080 34060
rect 27801 34051 27859 34057
rect 27801 34048 27813 34051
rect 27764 34020 27813 34048
rect 27764 34008 27770 34020
rect 27801 34017 27813 34020
rect 27847 34017 27859 34051
rect 28068 34048 28080 34057
rect 28035 34020 28080 34048
rect 27801 34011 27859 34017
rect 28068 34011 28080 34020
rect 28074 34008 28080 34011
rect 28132 34008 28138 34060
rect 28442 34008 28448 34060
rect 28500 34048 28506 34060
rect 29822 34048 29828 34060
rect 28500 34020 29040 34048
rect 29783 34020 29828 34048
rect 28500 34008 28506 34020
rect 29012 33980 29040 34020
rect 29822 34008 29828 34020
rect 29880 34008 29886 34060
rect 35618 34048 35624 34060
rect 35579 34020 35624 34048
rect 35618 34008 35624 34020
rect 35676 34008 35682 34060
rect 36189 34057 36217 34088
rect 36354 34076 36360 34088
rect 36412 34076 36418 34128
rect 36081 34051 36139 34057
rect 36081 34017 36093 34051
rect 36127 34017 36139 34051
rect 36081 34011 36139 34017
rect 36174 34051 36232 34057
rect 36174 34017 36186 34051
rect 36220 34017 36232 34051
rect 36446 34048 36452 34060
rect 36407 34020 36452 34048
rect 36174 34011 36232 34017
rect 30190 33980 30196 33992
rect 29012 33952 30196 33980
rect 30190 33940 30196 33952
rect 30248 33940 30254 33992
rect 30006 33872 30012 33924
rect 30064 33912 30070 33924
rect 36096 33912 36124 34011
rect 36446 34008 36452 34020
rect 36504 34008 36510 34060
rect 36587 34051 36645 34057
rect 36587 34017 36599 34051
rect 36633 34048 36645 34051
rect 36722 34048 36728 34060
rect 36633 34020 36728 34048
rect 36633 34017 36645 34020
rect 36587 34011 36645 34017
rect 36722 34008 36728 34020
rect 36780 34008 36786 34060
rect 37366 34048 37372 34060
rect 37327 34020 37372 34048
rect 37366 34008 37372 34020
rect 37424 34008 37430 34060
rect 36906 33912 36912 33924
rect 30064 33884 35848 33912
rect 36096 33884 36912 33912
rect 30064 33872 30070 33884
rect 27706 33844 27712 33856
rect 27586 33816 27712 33844
rect 27706 33804 27712 33816
rect 27764 33844 27770 33856
rect 29086 33844 29092 33856
rect 27764 33816 29092 33844
rect 27764 33804 27770 33816
rect 29086 33804 29092 33816
rect 29144 33804 29150 33856
rect 35437 33847 35495 33853
rect 35437 33813 35449 33847
rect 35483 33844 35495 33847
rect 35710 33844 35716 33856
rect 35483 33816 35716 33844
rect 35483 33813 35495 33816
rect 35437 33807 35495 33813
rect 35710 33804 35716 33816
rect 35768 33804 35774 33856
rect 35820 33844 35848 33884
rect 36906 33872 36912 33884
rect 36964 33872 36970 33924
rect 36725 33847 36783 33853
rect 36725 33844 36737 33847
rect 35820 33816 36737 33844
rect 36725 33813 36737 33816
rect 36771 33813 36783 33847
rect 36725 33807 36783 33813
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 25774 33640 25780 33652
rect 25735 33612 25780 33640
rect 25774 33600 25780 33612
rect 25832 33600 25838 33652
rect 38105 33643 38163 33649
rect 25884 33612 27384 33640
rect 2038 33572 2044 33584
rect 1999 33544 2044 33572
rect 2038 33532 2044 33544
rect 2096 33532 2102 33584
rect 18782 33532 18788 33584
rect 18840 33572 18846 33584
rect 25884 33572 25912 33612
rect 18840 33544 25912 33572
rect 18840 33532 18846 33544
rect 25774 33504 25780 33516
rect 25240 33476 25780 33504
rect 1854 33436 1860 33448
rect 1815 33408 1860 33436
rect 1854 33396 1860 33408
rect 1912 33396 1918 33448
rect 1946 33396 1952 33448
rect 2004 33436 2010 33448
rect 25240 33445 25268 33476
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 27356 33504 27384 33612
rect 28368 33612 31754 33640
rect 27982 33532 27988 33584
rect 28040 33572 28046 33584
rect 28261 33575 28319 33581
rect 28261 33572 28273 33575
rect 28040 33544 28273 33572
rect 28040 33532 28046 33544
rect 28261 33541 28273 33544
rect 28307 33541 28319 33575
rect 28261 33535 28319 33541
rect 28368 33504 28396 33612
rect 28442 33532 28448 33584
rect 28500 33532 28506 33584
rect 27356 33476 28396 33504
rect 28460 33504 28488 33532
rect 28537 33507 28595 33513
rect 28537 33504 28549 33507
rect 28460 33476 28549 33504
rect 28537 33473 28549 33476
rect 28583 33473 28595 33507
rect 28537 33467 28595 33473
rect 28721 33507 28779 33513
rect 28721 33473 28733 33507
rect 28767 33504 28779 33507
rect 28994 33504 29000 33516
rect 28767 33476 29000 33504
rect 28767 33473 28779 33476
rect 28721 33467 28779 33473
rect 28994 33464 29000 33476
rect 29052 33464 29058 33516
rect 31726 33504 31754 33612
rect 38105 33609 38117 33643
rect 38151 33640 38163 33643
rect 38194 33640 38200 33652
rect 38151 33612 38200 33640
rect 38151 33609 38163 33612
rect 38105 33603 38163 33609
rect 38194 33600 38200 33612
rect 38252 33600 38258 33652
rect 35894 33532 35900 33584
rect 35952 33572 35958 33584
rect 36170 33572 36176 33584
rect 35952 33544 36176 33572
rect 35952 33532 35958 33544
rect 36170 33532 36176 33544
rect 36228 33532 36234 33584
rect 37277 33575 37335 33581
rect 37277 33541 37289 33575
rect 37323 33572 37335 33575
rect 39022 33572 39028 33584
rect 37323 33544 39028 33572
rect 37323 33541 37335 33544
rect 37277 33535 37335 33541
rect 39022 33532 39028 33544
rect 39080 33532 39086 33584
rect 31726 33476 36400 33504
rect 25225 33439 25283 33445
rect 2004 33408 6914 33436
rect 2004 33396 2010 33408
rect 6886 33368 6914 33408
rect 25225 33405 25237 33439
rect 25271 33405 25283 33439
rect 25598 33439 25656 33445
rect 25598 33436 25610 33439
rect 25225 33399 25283 33405
rect 25332 33408 25610 33436
rect 25332 33368 25360 33408
rect 25598 33405 25610 33408
rect 25644 33405 25656 33439
rect 25598 33399 25656 33405
rect 25866 33396 25872 33448
rect 25924 33436 25930 33448
rect 26329 33439 26387 33445
rect 26329 33436 26341 33439
rect 25924 33408 26341 33436
rect 25924 33396 25930 33408
rect 26329 33405 26341 33408
rect 26375 33405 26387 33439
rect 26329 33399 26387 33405
rect 26596 33439 26654 33445
rect 26596 33405 26608 33439
rect 26642 33436 26654 33439
rect 26878 33436 26884 33448
rect 26642 33408 26884 33436
rect 26642 33405 26654 33408
rect 26596 33399 26654 33405
rect 6886 33340 25360 33368
rect 25409 33371 25467 33377
rect 25409 33337 25421 33371
rect 25455 33337 25467 33371
rect 25409 33331 25467 33337
rect 10134 33260 10140 33312
rect 10192 33300 10198 33312
rect 14458 33300 14464 33312
rect 10192 33272 14464 33300
rect 10192 33260 10198 33272
rect 14458 33260 14464 33272
rect 14516 33260 14522 33312
rect 25314 33260 25320 33312
rect 25372 33300 25378 33312
rect 25424 33300 25452 33331
rect 25498 33328 25504 33380
rect 25556 33368 25562 33380
rect 25556 33340 25601 33368
rect 25556 33328 25562 33340
rect 25372 33272 25452 33300
rect 26344 33300 26372 33399
rect 26878 33396 26884 33408
rect 26936 33396 26942 33448
rect 28350 33396 28356 33448
rect 28408 33436 28414 33448
rect 28445 33439 28503 33445
rect 28445 33436 28457 33439
rect 28408 33408 28457 33436
rect 28408 33396 28414 33408
rect 28445 33405 28457 33408
rect 28491 33405 28503 33439
rect 28445 33399 28503 33405
rect 28629 33439 28687 33445
rect 28629 33405 28641 33439
rect 28675 33405 28687 33439
rect 28896 33439 28954 33445
rect 28896 33436 28908 33439
rect 28629 33399 28687 33405
rect 28828 33408 28908 33436
rect 26510 33328 26516 33380
rect 26568 33368 26574 33380
rect 27062 33368 27068 33380
rect 26568 33340 27068 33368
rect 26568 33328 26574 33340
rect 27062 33328 27068 33340
rect 27120 33328 27126 33380
rect 28534 33328 28540 33380
rect 28592 33368 28598 33380
rect 28644 33368 28672 33399
rect 28592 33340 28672 33368
rect 28828 33368 28856 33408
rect 28896 33405 28908 33408
rect 28942 33405 28954 33439
rect 36078 33436 36084 33448
rect 36039 33408 36084 33436
rect 28896 33399 28954 33405
rect 36078 33396 36084 33408
rect 36136 33396 36142 33448
rect 36170 33396 36176 33448
rect 36228 33436 36234 33448
rect 36372 33436 36400 33476
rect 36546 33439 36604 33445
rect 36546 33436 36558 33439
rect 36228 33408 36273 33436
rect 36372 33408 36558 33436
rect 36228 33396 36234 33408
rect 36546 33405 36558 33408
rect 36592 33405 36604 33439
rect 37458 33436 37464 33448
rect 37419 33408 37464 33436
rect 36546 33399 36604 33405
rect 37458 33396 37464 33408
rect 37516 33396 37522 33448
rect 37921 33439 37979 33445
rect 37921 33405 37933 33439
rect 37967 33436 37979 33439
rect 38010 33436 38016 33448
rect 37967 33408 38016 33436
rect 37967 33405 37979 33408
rect 37921 33399 37979 33405
rect 38010 33396 38016 33408
rect 38068 33396 38074 33448
rect 29086 33368 29092 33380
rect 28828 33340 29092 33368
rect 28592 33328 28598 33340
rect 29086 33328 29092 33340
rect 29144 33328 29150 33380
rect 36354 33368 36360 33380
rect 36315 33340 36360 33368
rect 36354 33328 36360 33340
rect 36412 33328 36418 33380
rect 36446 33328 36452 33380
rect 36504 33368 36510 33380
rect 36504 33340 36549 33368
rect 36504 33328 36510 33340
rect 26878 33300 26884 33312
rect 26344 33272 26884 33300
rect 25372 33260 25378 33272
rect 26878 33260 26884 33272
rect 26936 33260 26942 33312
rect 27614 33260 27620 33312
rect 27672 33300 27678 33312
rect 27709 33303 27767 33309
rect 27709 33300 27721 33303
rect 27672 33272 27721 33300
rect 27672 33260 27678 33272
rect 27709 33269 27721 33272
rect 27755 33300 27767 33303
rect 29730 33300 29736 33312
rect 27755 33272 29736 33300
rect 27755 33269 27767 33272
rect 27709 33263 27767 33269
rect 29730 33260 29736 33272
rect 29788 33260 29794 33312
rect 35618 33260 35624 33312
rect 35676 33300 35682 33312
rect 36725 33303 36783 33309
rect 36725 33300 36737 33303
rect 35676 33272 36737 33300
rect 35676 33260 35682 33272
rect 36725 33269 36737 33272
rect 36771 33269 36783 33303
rect 36725 33263 36783 33269
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 1581 33099 1639 33105
rect 1581 33065 1593 33099
rect 1627 33096 1639 33099
rect 1946 33096 1952 33108
rect 1627 33068 1952 33096
rect 1627 33065 1639 33068
rect 1581 33059 1639 33065
rect 1946 33056 1952 33068
rect 2004 33056 2010 33108
rect 24670 33056 24676 33108
rect 24728 33096 24734 33108
rect 24728 33068 25641 33096
rect 24728 33056 24734 33068
rect 1854 32988 1860 33040
rect 1912 33028 1918 33040
rect 22830 33028 22836 33040
rect 1912 33000 22836 33028
rect 1912 32988 1918 33000
rect 22830 32988 22836 33000
rect 22888 32988 22894 33040
rect 25613 33028 25641 33068
rect 26878 33056 26884 33108
rect 26936 33096 26942 33108
rect 29178 33096 29184 33108
rect 26936 33068 27200 33096
rect 29139 33068 29184 33096
rect 26936 33056 26942 33068
rect 22940 33000 25549 33028
rect 25613 33000 27108 33028
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 1578 32852 1584 32904
rect 1636 32892 1642 32904
rect 22940 32892 22968 33000
rect 24854 32920 24860 32972
rect 24912 32960 24918 32972
rect 25133 32963 25191 32969
rect 25133 32960 25145 32963
rect 24912 32932 25145 32960
rect 24912 32920 24918 32932
rect 25133 32929 25145 32932
rect 25179 32929 25191 32963
rect 25314 32960 25320 32972
rect 25275 32932 25320 32960
rect 25133 32923 25191 32929
rect 25314 32920 25320 32932
rect 25372 32920 25378 32972
rect 25521 32969 25549 33000
rect 25409 32963 25467 32969
rect 25409 32929 25421 32963
rect 25455 32929 25467 32963
rect 25409 32923 25467 32929
rect 25506 32963 25564 32969
rect 25506 32929 25518 32963
rect 25552 32929 25564 32963
rect 26418 32960 26424 32972
rect 26379 32932 26424 32960
rect 25506 32923 25564 32929
rect 1636 32864 22968 32892
rect 25424 32892 25452 32923
rect 26418 32920 26424 32932
rect 26476 32920 26482 32972
rect 26510 32920 26516 32972
rect 26568 32960 26574 32972
rect 26697 32963 26755 32969
rect 26697 32960 26709 32963
rect 26568 32932 26709 32960
rect 26568 32920 26574 32932
rect 26697 32929 26709 32932
rect 26743 32929 26755 32963
rect 26697 32923 26755 32929
rect 26881 32963 26939 32969
rect 26881 32929 26893 32963
rect 26927 32929 26939 32963
rect 26881 32923 26939 32929
rect 25424 32864 25544 32892
rect 1636 32852 1642 32864
rect 25516 32836 25544 32864
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26605 32895 26663 32901
rect 26384 32864 26556 32892
rect 26384 32852 26390 32864
rect 25498 32784 25504 32836
rect 25556 32784 25562 32836
rect 25682 32824 25688 32836
rect 25643 32796 25688 32824
rect 25682 32784 25688 32796
rect 25740 32784 25746 32836
rect 26528 32833 26556 32864
rect 26605 32861 26617 32895
rect 26651 32861 26663 32895
rect 26605 32855 26663 32861
rect 26513 32827 26571 32833
rect 26513 32793 26525 32827
rect 26559 32793 26571 32827
rect 26513 32787 26571 32793
rect 26237 32759 26295 32765
rect 26237 32725 26249 32759
rect 26283 32756 26295 32759
rect 26326 32756 26332 32768
rect 26283 32728 26332 32756
rect 26283 32725 26295 32728
rect 26237 32719 26295 32725
rect 26326 32716 26332 32728
rect 26384 32716 26390 32768
rect 26620 32756 26648 32855
rect 26896 32824 26924 32923
rect 27080 32892 27108 33000
rect 27172 32960 27200 33068
rect 29178 33056 29184 33068
rect 29236 33056 29242 33108
rect 32858 33096 32864 33108
rect 31726 33068 32864 33096
rect 27890 32988 27896 33040
rect 27948 33028 27954 33040
rect 28046 33031 28104 33037
rect 28046 33028 28058 33031
rect 27948 33000 28058 33028
rect 27948 32988 27954 33000
rect 28046 32997 28058 33000
rect 28092 32997 28104 33031
rect 28046 32991 28104 32997
rect 27801 32963 27859 32969
rect 27801 32960 27813 32963
rect 27172 32932 27813 32960
rect 27801 32929 27813 32932
rect 27847 32929 27859 32963
rect 31726 32960 31754 33068
rect 32858 33056 32864 33068
rect 32916 33056 32922 33108
rect 33962 33056 33968 33108
rect 34020 33096 34026 33108
rect 35621 33099 35679 33105
rect 35621 33096 35633 33099
rect 34020 33068 35633 33096
rect 34020 33056 34026 33068
rect 35621 33065 35633 33068
rect 35667 33065 35679 33099
rect 35621 33059 35679 33065
rect 36538 33056 36544 33108
rect 36596 33096 36602 33108
rect 37185 33099 37243 33105
rect 37185 33096 37197 33099
rect 36596 33068 37197 33096
rect 36596 33056 36602 33068
rect 37185 33065 37197 33068
rect 37231 33065 37243 33099
rect 37185 33059 37243 33065
rect 36354 33028 36360 33040
rect 36315 33000 36360 33028
rect 36354 32988 36360 33000
rect 36412 32988 36418 33040
rect 27801 32923 27859 32929
rect 27908 32932 31754 32960
rect 27908 32892 27936 32932
rect 33962 32920 33968 32972
rect 34020 32960 34026 32972
rect 34146 32960 34152 32972
rect 34020 32932 34152 32960
rect 34020 32920 34026 32932
rect 34146 32920 34152 32932
rect 34204 32920 34210 32972
rect 35434 32960 35440 32972
rect 35395 32932 35440 32960
rect 35434 32920 35440 32932
rect 35492 32920 35498 32972
rect 36078 32960 36084 32972
rect 36039 32932 36084 32960
rect 36078 32920 36084 32932
rect 36136 32920 36142 32972
rect 36229 32963 36287 32969
rect 36229 32929 36241 32963
rect 36275 32929 36287 32963
rect 36446 32960 36452 32972
rect 36407 32932 36452 32960
rect 36229 32923 36287 32929
rect 27080 32864 27936 32892
rect 36244 32892 36272 32923
rect 36446 32920 36452 32932
rect 36504 32920 36510 32972
rect 36538 32920 36544 32972
rect 36596 32969 36602 32972
rect 36596 32960 36604 32969
rect 37366 32960 37372 32972
rect 36596 32932 36641 32960
rect 37327 32932 37372 32960
rect 36596 32923 36604 32932
rect 36596 32920 36602 32923
rect 37366 32920 37372 32932
rect 37424 32920 37430 32972
rect 37642 32892 37648 32904
rect 36244 32864 37648 32892
rect 37642 32852 37648 32864
rect 37700 32852 37706 32904
rect 27706 32824 27712 32836
rect 26896 32796 27712 32824
rect 27706 32784 27712 32796
rect 27764 32784 27770 32836
rect 29914 32824 29920 32836
rect 28966 32796 29920 32824
rect 26970 32756 26976 32768
rect 26620 32728 26976 32756
rect 26970 32716 26976 32728
rect 27028 32716 27034 32768
rect 27982 32716 27988 32768
rect 28040 32756 28046 32768
rect 28966 32756 28994 32796
rect 29914 32784 29920 32796
rect 29972 32784 29978 32836
rect 35250 32784 35256 32836
rect 35308 32824 35314 32836
rect 36725 32827 36783 32833
rect 36725 32824 36737 32827
rect 35308 32796 36737 32824
rect 35308 32784 35314 32796
rect 36725 32793 36737 32796
rect 36771 32793 36783 32827
rect 36725 32787 36783 32793
rect 28040 32728 28994 32756
rect 28040 32716 28046 32728
rect 29270 32716 29276 32768
rect 29328 32756 29334 32768
rect 30650 32756 30656 32768
rect 29328 32728 30656 32756
rect 29328 32716 29334 32728
rect 30650 32716 30656 32728
rect 30708 32716 30714 32768
rect 36354 32716 36360 32768
rect 36412 32756 36418 32768
rect 37182 32756 37188 32768
rect 36412 32728 37188 32756
rect 36412 32716 36418 32728
rect 37182 32716 37188 32728
rect 37240 32716 37246 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 25961 32555 26019 32561
rect 19306 32524 25825 32552
rect 19306 32416 19334 32524
rect 23845 32487 23903 32493
rect 23845 32453 23857 32487
rect 23891 32484 23903 32487
rect 24026 32484 24032 32496
rect 23891 32456 24032 32484
rect 23891 32453 23903 32456
rect 23845 32447 23903 32453
rect 24026 32444 24032 32456
rect 24084 32444 24090 32496
rect 25222 32444 25228 32496
rect 25280 32444 25286 32496
rect 25498 32444 25504 32496
rect 25556 32484 25562 32496
rect 25682 32484 25688 32496
rect 25556 32456 25688 32484
rect 25556 32444 25562 32456
rect 25682 32444 25688 32456
rect 25740 32444 25746 32496
rect 6886 32388 19334 32416
rect 25240 32416 25268 32444
rect 25240 32388 25452 32416
rect 4706 32308 4712 32360
rect 4764 32348 4770 32360
rect 6886 32348 6914 32388
rect 4764 32320 6914 32348
rect 4764 32308 4770 32320
rect 25314 32308 25320 32360
rect 25372 32308 25378 32360
rect 25424 32357 25452 32388
rect 25797 32357 25825 32524
rect 25961 32521 25973 32555
rect 26007 32552 26019 32555
rect 26050 32552 26056 32564
rect 26007 32524 26056 32552
rect 26007 32521 26019 32524
rect 25961 32515 26019 32521
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 26970 32552 26976 32564
rect 26897 32524 26976 32552
rect 26897 32425 26925 32524
rect 26970 32512 26976 32524
rect 27028 32512 27034 32564
rect 27706 32552 27712 32564
rect 27172 32524 27712 32552
rect 26881 32419 26939 32425
rect 26881 32385 26893 32419
rect 26927 32385 26939 32419
rect 26881 32379 26939 32385
rect 26970 32376 26976 32428
rect 27028 32416 27034 32428
rect 27028 32388 27073 32416
rect 27028 32376 27034 32388
rect 27172 32357 27200 32524
rect 27706 32512 27712 32524
rect 27764 32512 27770 32564
rect 28166 32552 28172 32564
rect 28127 32524 28172 32552
rect 28166 32512 28172 32524
rect 28224 32512 28230 32564
rect 36265 32555 36323 32561
rect 36265 32521 36277 32555
rect 36311 32552 36323 32555
rect 36446 32552 36452 32564
rect 36311 32524 36452 32552
rect 36311 32521 36323 32524
rect 36265 32515 36323 32521
rect 36446 32512 36452 32524
rect 36504 32512 36510 32564
rect 36538 32512 36544 32564
rect 36596 32512 36602 32564
rect 36722 32512 36728 32564
rect 36780 32552 36786 32564
rect 37093 32555 37151 32561
rect 37093 32552 37105 32555
rect 36780 32524 37105 32552
rect 36780 32512 36786 32524
rect 37093 32521 37105 32524
rect 37139 32521 37151 32555
rect 37093 32515 37151 32521
rect 27356 32456 27844 32484
rect 25409 32351 25467 32357
rect 25409 32317 25421 32351
rect 25455 32317 25467 32351
rect 25409 32311 25467 32317
rect 25782 32351 25840 32357
rect 25782 32317 25794 32351
rect 25828 32317 25840 32351
rect 25782 32311 25840 32317
rect 26697 32351 26755 32357
rect 26697 32317 26709 32351
rect 26743 32317 26755 32351
rect 26697 32311 26755 32317
rect 26789 32351 26847 32357
rect 26789 32317 26801 32351
rect 26835 32348 26847 32351
rect 27157 32351 27215 32357
rect 26835 32317 26849 32348
rect 26789 32311 26849 32317
rect 27157 32317 27169 32351
rect 27203 32317 27215 32351
rect 27157 32311 27215 32317
rect 22830 32240 22836 32292
rect 22888 32280 22894 32292
rect 23661 32283 23719 32289
rect 23661 32280 23673 32283
rect 22888 32252 23673 32280
rect 22888 32240 22894 32252
rect 23661 32249 23673 32252
rect 23707 32280 23719 32283
rect 24302 32280 24308 32292
rect 23707 32252 24308 32280
rect 23707 32249 23719 32252
rect 23661 32243 23719 32249
rect 24302 32240 24308 32252
rect 24360 32240 24366 32292
rect 25332 32280 25360 32308
rect 25593 32283 25651 32289
rect 25593 32280 25605 32283
rect 25332 32252 25605 32280
rect 25593 32249 25605 32252
rect 25639 32249 25651 32283
rect 25593 32243 25651 32249
rect 25682 32240 25688 32292
rect 25740 32280 25746 32292
rect 25740 32252 25785 32280
rect 25740 32240 25746 32252
rect 25314 32172 25320 32224
rect 25372 32212 25378 32224
rect 26513 32215 26571 32221
rect 26513 32212 26525 32215
rect 25372 32184 26525 32212
rect 25372 32172 25378 32184
rect 26513 32181 26525 32184
rect 26559 32181 26571 32215
rect 26712 32212 26740 32311
rect 26821 32280 26849 32311
rect 27356 32280 27384 32456
rect 27430 32376 27436 32428
rect 27488 32416 27494 32428
rect 27816 32416 27844 32456
rect 27890 32444 27896 32496
rect 27948 32484 27954 32496
rect 36556 32484 36584 32512
rect 39482 32484 39488 32496
rect 27948 32456 36584 32484
rect 37016 32456 39488 32484
rect 27948 32444 27954 32456
rect 31754 32416 31760 32428
rect 27488 32388 27752 32416
rect 27816 32388 31760 32416
rect 27488 32376 27494 32388
rect 27617 32351 27675 32357
rect 27617 32317 27629 32351
rect 27663 32348 27675 32351
rect 27724 32348 27752 32388
rect 31754 32376 31760 32388
rect 31812 32376 31818 32428
rect 36538 32376 36544 32428
rect 36596 32416 36602 32428
rect 37016 32416 37044 32456
rect 39482 32444 39488 32456
rect 39540 32444 39546 32496
rect 38378 32416 38384 32428
rect 36596 32388 37044 32416
rect 37568 32388 38384 32416
rect 36596 32376 36602 32388
rect 27801 32351 27859 32357
rect 27801 32348 27813 32351
rect 27663 32317 27680 32348
rect 27724 32320 27813 32348
rect 27617 32311 27680 32317
rect 27801 32317 27813 32320
rect 27847 32317 27859 32351
rect 27982 32348 27988 32360
rect 28040 32357 28046 32360
rect 27948 32320 27988 32348
rect 27801 32311 27859 32317
rect 26821 32252 27384 32280
rect 27338 32212 27344 32224
rect 26712 32184 27344 32212
rect 26513 32175 26571 32181
rect 27338 32172 27344 32184
rect 27396 32172 27402 32224
rect 27652 32212 27680 32311
rect 27982 32308 27988 32320
rect 28040 32311 28048 32357
rect 28040 32308 28046 32311
rect 28258 32308 28264 32360
rect 28316 32348 28322 32360
rect 28626 32348 28632 32360
rect 28316 32320 28632 32348
rect 28316 32308 28322 32320
rect 28626 32308 28632 32320
rect 28684 32308 28690 32360
rect 35894 32308 35900 32360
rect 35952 32348 35958 32360
rect 36081 32351 36139 32357
rect 36081 32348 36093 32351
rect 35952 32320 36093 32348
rect 35952 32308 35958 32320
rect 36081 32317 36093 32320
rect 36127 32348 36139 32351
rect 36722 32348 36728 32360
rect 36127 32320 36728 32348
rect 36127 32317 36139 32320
rect 36081 32311 36139 32317
rect 36722 32308 36728 32320
rect 36780 32308 36786 32360
rect 36906 32348 36912 32360
rect 36867 32320 36912 32348
rect 36906 32308 36912 32320
rect 36964 32308 36970 32360
rect 37568 32357 37596 32388
rect 38378 32376 38384 32388
rect 38436 32376 38442 32428
rect 37553 32351 37611 32357
rect 37553 32317 37565 32351
rect 37599 32317 37611 32351
rect 37553 32311 37611 32317
rect 37921 32351 37979 32357
rect 37921 32317 37933 32351
rect 37967 32348 37979 32351
rect 38930 32348 38936 32360
rect 37967 32320 38936 32348
rect 37967 32317 37979 32320
rect 37921 32311 37979 32317
rect 38930 32308 38936 32320
rect 38988 32308 38994 32360
rect 27890 32240 27896 32292
rect 27948 32280 27954 32292
rect 31570 32280 31576 32292
rect 27948 32252 27993 32280
rect 28966 32252 31576 32280
rect 27948 32240 27954 32252
rect 27982 32212 27988 32224
rect 27652 32184 27988 32212
rect 27982 32172 27988 32184
rect 28040 32172 28046 32224
rect 28626 32172 28632 32224
rect 28684 32212 28690 32224
rect 28966 32212 28994 32252
rect 31570 32240 31576 32252
rect 31628 32240 31634 32292
rect 37734 32280 37740 32292
rect 37695 32252 37740 32280
rect 37734 32240 37740 32252
rect 37792 32240 37798 32292
rect 37826 32240 37832 32292
rect 37884 32280 37890 32292
rect 37884 32252 37929 32280
rect 37884 32240 37890 32252
rect 28684 32184 28994 32212
rect 28684 32172 28690 32184
rect 37458 32172 37464 32224
rect 37516 32212 37522 32224
rect 38105 32215 38163 32221
rect 38105 32212 38117 32215
rect 37516 32184 38117 32212
rect 37516 32172 37522 32184
rect 38105 32181 38117 32184
rect 38151 32181 38163 32215
rect 38105 32175 38163 32181
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 1578 32008 1584 32020
rect 1539 31980 1584 32008
rect 1578 31968 1584 31980
rect 1636 31968 1642 32020
rect 12406 31980 25360 32008
rect 2774 31900 2780 31952
rect 2832 31940 2838 31952
rect 2832 31912 6914 31940
rect 2832 31900 2838 31912
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 6886 31804 6914 31912
rect 12406 31804 12434 31980
rect 15286 31900 15292 31952
rect 15344 31940 15350 31952
rect 23382 31940 23388 31952
rect 15344 31912 23388 31940
rect 15344 31900 15350 31912
rect 23382 31900 23388 31912
rect 23440 31900 23446 31952
rect 24765 31943 24823 31949
rect 24765 31909 24777 31943
rect 24811 31940 24823 31943
rect 24946 31940 24952 31952
rect 24811 31912 24952 31940
rect 24811 31909 24823 31912
rect 24765 31903 24823 31909
rect 24946 31900 24952 31912
rect 25004 31900 25010 31952
rect 22094 31832 22100 31884
rect 22152 31872 22158 31884
rect 22557 31875 22615 31881
rect 22557 31872 22569 31875
rect 22152 31844 22569 31872
rect 22152 31832 22158 31844
rect 22557 31841 22569 31844
rect 22603 31841 22615 31875
rect 22557 31835 22615 31841
rect 22649 31875 22707 31881
rect 22649 31841 22661 31875
rect 22695 31872 22707 31875
rect 22830 31872 22836 31884
rect 22695 31844 22836 31872
rect 22695 31841 22707 31844
rect 22649 31835 22707 31841
rect 22830 31832 22836 31844
rect 22888 31832 22894 31884
rect 24670 31832 24676 31884
rect 24728 31872 24734 31884
rect 24857 31875 24915 31881
rect 24857 31872 24869 31875
rect 24728 31844 24869 31872
rect 24728 31832 24734 31844
rect 24857 31841 24869 31844
rect 24903 31841 24915 31875
rect 25041 31875 25099 31881
rect 25041 31872 25053 31875
rect 24857 31835 24915 31841
rect 24964 31844 25053 31872
rect 6886 31776 12434 31804
rect 24765 31671 24823 31677
rect 24765 31637 24777 31671
rect 24811 31668 24823 31671
rect 24854 31668 24860 31680
rect 24811 31640 24860 31668
rect 24811 31637 24823 31640
rect 24765 31631 24823 31637
rect 24854 31628 24860 31640
rect 24912 31628 24918 31680
rect 24964 31668 24992 31844
rect 25041 31841 25053 31844
rect 25087 31841 25099 31875
rect 25041 31835 25099 31841
rect 25133 31875 25191 31881
rect 25133 31841 25145 31875
rect 25179 31841 25191 31875
rect 25133 31835 25191 31841
rect 25230 31875 25288 31881
rect 25230 31841 25242 31875
rect 25276 31872 25288 31875
rect 25332 31872 25360 31980
rect 25682 31968 25688 32020
rect 25740 32008 25746 32020
rect 26050 32008 26056 32020
rect 25740 31980 26056 32008
rect 25740 31968 25746 31980
rect 26050 31968 26056 31980
rect 26108 31968 26114 32020
rect 27522 31968 27528 32020
rect 27580 32008 27586 32020
rect 27890 32008 27896 32020
rect 27580 31980 27896 32008
rect 27580 31968 27586 31980
rect 27890 31968 27896 31980
rect 27948 32008 27954 32020
rect 28350 32008 28356 32020
rect 28408 32017 28414 32020
rect 27948 31980 28120 32008
rect 28319 31980 28356 32008
rect 27948 31968 27954 31980
rect 25498 31900 25504 31952
rect 25556 31940 25562 31952
rect 26237 31943 26295 31949
rect 26237 31940 26249 31943
rect 25556 31912 26249 31940
rect 25556 31900 25562 31912
rect 26237 31909 26249 31912
rect 26283 31909 26295 31943
rect 26237 31903 26295 31909
rect 27430 31900 27436 31952
rect 27488 31940 27494 31952
rect 28092 31949 28120 31980
rect 28350 31968 28356 31980
rect 28408 31971 28419 32017
rect 28408 31968 28414 31971
rect 30926 31968 30932 32020
rect 30984 32008 30990 32020
rect 35713 32011 35771 32017
rect 35713 32008 35725 32011
rect 30984 31980 35725 32008
rect 30984 31968 30990 31980
rect 35713 31977 35725 31980
rect 35759 31977 35771 32011
rect 35713 31971 35771 31977
rect 36357 32011 36415 32017
rect 36357 31977 36369 32011
rect 36403 31977 36415 32011
rect 37182 32008 37188 32020
rect 36357 31971 36415 31977
rect 37016 31980 37188 32008
rect 27985 31943 28043 31949
rect 27985 31940 27997 31943
rect 27488 31912 27997 31940
rect 27488 31900 27494 31912
rect 27985 31909 27997 31912
rect 28031 31909 28043 31943
rect 27985 31903 28043 31909
rect 28077 31943 28135 31949
rect 28077 31909 28089 31943
rect 28123 31909 28135 31943
rect 28077 31903 28135 31909
rect 25276 31844 25360 31872
rect 25961 31875 26019 31881
rect 25276 31841 25288 31844
rect 25230 31835 25288 31841
rect 25961 31841 25973 31875
rect 26007 31872 26019 31875
rect 26050 31872 26056 31884
rect 26007 31844 26056 31872
rect 26007 31841 26019 31844
rect 25961 31835 26019 31841
rect 25148 31804 25176 31835
rect 26050 31832 26056 31844
rect 26108 31832 26114 31884
rect 26145 31875 26203 31881
rect 26145 31841 26157 31875
rect 26191 31841 26203 31875
rect 26145 31835 26203 31841
rect 26381 31875 26439 31881
rect 26381 31841 26393 31875
rect 26427 31872 26439 31875
rect 26878 31872 26884 31884
rect 26427 31844 26884 31872
rect 26427 31841 26439 31844
rect 26381 31835 26439 31841
rect 25498 31804 25504 31816
rect 25148 31776 25504 31804
rect 25498 31764 25504 31776
rect 25556 31764 25562 31816
rect 25038 31696 25044 31748
rect 25096 31736 25102 31748
rect 25409 31739 25467 31745
rect 25409 31736 25421 31739
rect 25096 31708 25421 31736
rect 25096 31696 25102 31708
rect 25409 31705 25421 31708
rect 25455 31705 25467 31739
rect 26160 31736 26188 31835
rect 26878 31832 26884 31844
rect 26936 31832 26942 31884
rect 27798 31872 27804 31884
rect 27759 31844 27804 31872
rect 27798 31832 27804 31844
rect 27856 31832 27862 31884
rect 27890 31832 27896 31884
rect 27948 31872 27954 31884
rect 28174 31875 28232 31881
rect 28174 31872 28186 31875
rect 27948 31844 28186 31872
rect 27948 31832 27954 31844
rect 28174 31841 28186 31844
rect 28220 31841 28232 31875
rect 28174 31835 28232 31841
rect 34146 31832 34152 31884
rect 34204 31872 34210 31884
rect 34514 31872 34520 31884
rect 34204 31844 34520 31872
rect 34204 31832 34210 31844
rect 34514 31832 34520 31844
rect 34572 31832 34578 31884
rect 35526 31872 35532 31884
rect 35487 31844 35532 31872
rect 35526 31832 35532 31844
rect 35584 31832 35590 31884
rect 36170 31872 36176 31884
rect 36131 31844 36176 31872
rect 36170 31832 36176 31844
rect 36228 31832 36234 31884
rect 36372 31872 36400 31971
rect 36446 31900 36452 31952
rect 36504 31940 36510 31952
rect 37016 31949 37044 31980
rect 37182 31968 37188 31980
rect 37240 31968 37246 32020
rect 37001 31943 37059 31949
rect 37001 31940 37013 31943
rect 36504 31912 37013 31940
rect 36504 31900 36510 31912
rect 37001 31909 37013 31912
rect 37047 31909 37059 31943
rect 37001 31903 37059 31909
rect 37093 31943 37151 31949
rect 37093 31909 37105 31943
rect 37139 31940 37151 31943
rect 37826 31940 37832 31952
rect 37139 31912 37832 31940
rect 37139 31909 37151 31912
rect 37093 31903 37151 31909
rect 37826 31900 37832 31912
rect 37884 31900 37890 31952
rect 36372 31844 36492 31872
rect 33318 31764 33324 31816
rect 33376 31804 33382 31816
rect 34330 31804 34336 31816
rect 33376 31776 34336 31804
rect 33376 31764 33382 31776
rect 34330 31764 34336 31776
rect 34388 31764 34394 31816
rect 36464 31804 36492 31844
rect 36538 31832 36544 31884
rect 36596 31872 36602 31884
rect 36817 31875 36875 31881
rect 36817 31872 36829 31875
rect 36596 31844 36829 31872
rect 36596 31832 36602 31844
rect 36817 31841 36829 31844
rect 36863 31841 36875 31875
rect 37182 31872 37188 31884
rect 37143 31844 37188 31872
rect 36817 31835 36875 31841
rect 37182 31832 37188 31844
rect 37240 31832 37246 31884
rect 38838 31804 38844 31816
rect 36464 31776 38844 31804
rect 38838 31764 38844 31776
rect 38896 31764 38902 31816
rect 25409 31699 25467 31705
rect 25507 31708 26188 31736
rect 25222 31668 25228 31680
rect 24964 31640 25228 31668
rect 25222 31628 25228 31640
rect 25280 31668 25286 31680
rect 25507 31668 25535 31708
rect 26234 31696 26240 31748
rect 26292 31736 26298 31748
rect 26513 31739 26571 31745
rect 26513 31736 26525 31739
rect 26292 31708 26525 31736
rect 26292 31696 26298 31708
rect 26513 31705 26525 31708
rect 26559 31705 26571 31739
rect 26513 31699 26571 31705
rect 26970 31696 26976 31748
rect 27028 31736 27034 31748
rect 27338 31736 27344 31748
rect 27028 31708 27344 31736
rect 27028 31696 27034 31708
rect 27338 31696 27344 31708
rect 27396 31696 27402 31748
rect 34146 31696 34152 31748
rect 34204 31736 34210 31748
rect 34790 31736 34796 31748
rect 34204 31708 34796 31736
rect 34204 31696 34210 31708
rect 34790 31696 34796 31708
rect 34848 31696 34854 31748
rect 35894 31696 35900 31748
rect 35952 31736 35958 31748
rect 36722 31736 36728 31748
rect 35952 31708 36728 31736
rect 35952 31696 35958 31708
rect 36722 31696 36728 31708
rect 36780 31696 36786 31748
rect 25280 31640 25535 31668
rect 25280 31628 25286 31640
rect 36538 31628 36544 31680
rect 36596 31668 36602 31680
rect 36998 31668 37004 31680
rect 36596 31640 37004 31668
rect 36596 31628 36602 31640
rect 36998 31628 37004 31640
rect 37056 31628 37062 31680
rect 37366 31668 37372 31680
rect 37327 31640 37372 31668
rect 37366 31628 37372 31640
rect 37424 31628 37430 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 1581 31467 1639 31473
rect 1581 31433 1593 31467
rect 1627 31464 1639 31467
rect 1854 31464 1860 31476
rect 1627 31436 1860 31464
rect 1627 31433 1639 31436
rect 1581 31427 1639 31433
rect 1854 31424 1860 31436
rect 1912 31424 1918 31476
rect 27617 31467 27675 31473
rect 26252 31436 27568 31464
rect 26252 31405 26280 31436
rect 26237 31399 26295 31405
rect 26237 31365 26249 31399
rect 26283 31365 26295 31399
rect 26878 31396 26884 31408
rect 26237 31359 26295 31365
rect 26344 31368 26884 31396
rect 2038 31288 2044 31340
rect 2096 31328 2102 31340
rect 23566 31328 23572 31340
rect 2096 31300 23572 31328
rect 2096 31288 2102 31300
rect 23566 31288 23572 31300
rect 23624 31288 23630 31340
rect 26344 31337 26372 31368
rect 26878 31356 26884 31368
rect 26936 31356 26942 31408
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31297 26387 31331
rect 26329 31291 26387 31297
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31328 26479 31331
rect 26786 31328 26792 31340
rect 26467 31300 26792 31328
rect 26467 31297 26479 31300
rect 26421 31291 26479 31297
rect 26786 31288 26792 31300
rect 26844 31288 26850 31340
rect 27338 31328 27344 31340
rect 27080 31300 27344 31328
rect 1394 31260 1400 31272
rect 1355 31232 1400 31260
rect 1394 31220 1400 31232
rect 1452 31220 1458 31272
rect 26145 31263 26203 31269
rect 26145 31260 26157 31263
rect 22066 31232 26157 31260
rect 21726 31152 21732 31204
rect 21784 31192 21790 31204
rect 22066 31192 22094 31232
rect 26145 31229 26157 31232
rect 26191 31229 26203 31263
rect 26145 31223 26203 31229
rect 26605 31263 26663 31269
rect 26605 31229 26617 31263
rect 26651 31260 26663 31263
rect 26878 31260 26884 31272
rect 26651 31232 26884 31260
rect 26651 31229 26663 31232
rect 26605 31223 26663 31229
rect 26878 31220 26884 31232
rect 26936 31220 26942 31272
rect 27080 31269 27108 31300
rect 27338 31288 27344 31300
rect 27396 31288 27402 31340
rect 27540 31328 27568 31436
rect 27617 31433 27629 31467
rect 27663 31464 27675 31467
rect 27706 31464 27712 31476
rect 27663 31436 27712 31464
rect 27663 31433 27675 31436
rect 27617 31427 27675 31433
rect 27706 31424 27712 31436
rect 27764 31424 27770 31476
rect 28353 31467 28411 31473
rect 28353 31433 28365 31467
rect 28399 31464 28411 31467
rect 28534 31464 28540 31476
rect 28399 31436 28540 31464
rect 28399 31433 28411 31436
rect 28353 31427 28411 31433
rect 28534 31424 28540 31436
rect 28592 31424 28598 31476
rect 36446 31464 36452 31476
rect 36359 31436 36452 31464
rect 36446 31424 36452 31436
rect 36504 31464 36510 31476
rect 37734 31464 37740 31476
rect 36504 31436 37740 31464
rect 36504 31424 36510 31436
rect 37734 31424 37740 31436
rect 37792 31424 37798 31476
rect 27890 31356 27896 31408
rect 27948 31396 27954 31408
rect 31018 31396 31024 31408
rect 27948 31368 31024 31396
rect 27948 31356 27954 31368
rect 31018 31356 31024 31368
rect 31076 31356 31082 31408
rect 31110 31328 31116 31340
rect 27540 31300 31116 31328
rect 31110 31288 31116 31300
rect 31168 31288 31174 31340
rect 27522 31269 27528 31272
rect 27065 31263 27123 31269
rect 27065 31229 27077 31263
rect 27111 31229 27123 31263
rect 27065 31223 27123 31229
rect 27485 31263 27528 31269
rect 27485 31229 27497 31263
rect 27485 31223 27528 31229
rect 27522 31220 27528 31223
rect 27580 31220 27586 31272
rect 27890 31220 27896 31272
rect 27948 31260 27954 31272
rect 28169 31263 28227 31269
rect 28169 31260 28181 31263
rect 27948 31232 28181 31260
rect 27948 31220 27954 31232
rect 28169 31229 28181 31232
rect 28215 31260 28227 31263
rect 29822 31260 29828 31272
rect 28215 31232 29828 31260
rect 28215 31229 28227 31232
rect 28169 31223 28227 31229
rect 29822 31220 29828 31232
rect 29880 31220 29886 31272
rect 25314 31192 25320 31204
rect 21784 31164 22094 31192
rect 25275 31164 25320 31192
rect 21784 31152 21790 31164
rect 25314 31152 25320 31164
rect 25372 31152 25378 31204
rect 27249 31195 27307 31201
rect 27249 31161 27261 31195
rect 27295 31161 27307 31195
rect 27249 31155 27307 31161
rect 9306 31084 9312 31136
rect 9364 31124 9370 31136
rect 20070 31124 20076 31136
rect 9364 31096 20076 31124
rect 9364 31084 9370 31096
rect 20070 31084 20076 31096
rect 20128 31084 20134 31136
rect 24946 31084 24952 31136
rect 25004 31124 25010 31136
rect 25409 31127 25467 31133
rect 25409 31124 25421 31127
rect 25004 31096 25421 31124
rect 25004 31084 25010 31096
rect 25409 31093 25421 31096
rect 25455 31093 25467 31127
rect 25409 31087 25467 31093
rect 25498 31084 25504 31136
rect 25556 31124 25562 31136
rect 25961 31127 26019 31133
rect 25961 31124 25973 31127
rect 25556 31096 25973 31124
rect 25556 31084 25562 31096
rect 25961 31093 25973 31096
rect 26007 31093 26019 31127
rect 27264 31124 27292 31155
rect 27338 31152 27344 31204
rect 27396 31192 27402 31204
rect 36464 31192 36492 31424
rect 38654 31396 38660 31408
rect 36740 31368 38660 31396
rect 36541 31263 36599 31269
rect 36541 31229 36553 31263
rect 36587 31260 36599 31263
rect 36740 31260 36768 31368
rect 38654 31356 38660 31368
rect 38712 31356 38718 31408
rect 39114 31328 39120 31340
rect 37568 31300 39120 31328
rect 36906 31260 36912 31272
rect 36587 31232 36768 31260
rect 36867 31232 36912 31260
rect 36587 31229 36599 31232
rect 36541 31223 36599 31229
rect 36906 31220 36912 31232
rect 36964 31220 36970 31272
rect 37568 31269 37596 31300
rect 39114 31288 39120 31300
rect 39172 31288 39178 31340
rect 37553 31263 37611 31269
rect 37553 31229 37565 31263
rect 37599 31229 37611 31263
rect 37826 31260 37832 31272
rect 37553 31223 37611 31229
rect 37660 31232 37832 31260
rect 36725 31195 36783 31201
rect 36725 31192 36737 31195
rect 27396 31164 27441 31192
rect 36464 31164 36737 31192
rect 27396 31152 27402 31164
rect 36725 31161 36737 31164
rect 36771 31161 36783 31195
rect 36725 31155 36783 31161
rect 36817 31195 36875 31201
rect 36817 31161 36829 31195
rect 36863 31192 36875 31195
rect 37274 31192 37280 31204
rect 36863 31164 37280 31192
rect 36863 31161 36875 31164
rect 36817 31155 36875 31161
rect 37274 31152 37280 31164
rect 37332 31192 37338 31204
rect 37660 31192 37688 31232
rect 37826 31220 37832 31232
rect 37884 31220 37890 31272
rect 37921 31263 37979 31269
rect 37921 31229 37933 31263
rect 37967 31260 37979 31263
rect 38010 31260 38016 31272
rect 37967 31232 38016 31260
rect 37967 31229 37979 31232
rect 37921 31223 37979 31229
rect 38010 31220 38016 31232
rect 38068 31220 38074 31272
rect 37332 31164 37688 31192
rect 37332 31152 37338 31164
rect 37734 31152 37740 31204
rect 37792 31192 37798 31204
rect 37792 31164 37837 31192
rect 37792 31152 37798 31164
rect 32490 31124 32496 31136
rect 27264 31096 32496 31124
rect 25961 31087 26019 31093
rect 32490 31084 32496 31096
rect 32548 31084 32554 31136
rect 36998 31084 37004 31136
rect 37056 31124 37062 31136
rect 37093 31127 37151 31133
rect 37093 31124 37105 31127
rect 37056 31096 37105 31124
rect 37056 31084 37062 31096
rect 37093 31093 37105 31096
rect 37139 31093 37151 31127
rect 37093 31087 37151 31093
rect 37182 31084 37188 31136
rect 37240 31124 37246 31136
rect 38105 31127 38163 31133
rect 38105 31124 38117 31127
rect 37240 31096 38117 31124
rect 37240 31084 37246 31096
rect 38105 31093 38117 31096
rect 38151 31093 38163 31127
rect 38105 31087 38163 31093
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 24946 30880 24952 30932
rect 25004 30920 25010 30932
rect 27890 30920 27896 30932
rect 25004 30892 27896 30920
rect 25004 30880 25010 30892
rect 25038 30812 25044 30864
rect 25096 30852 25102 30864
rect 25406 30852 25412 30864
rect 25096 30824 25412 30852
rect 25096 30812 25102 30824
rect 25406 30812 25412 30824
rect 25464 30812 25470 30864
rect 25584 30855 25642 30861
rect 25584 30821 25596 30855
rect 25630 30852 25642 30855
rect 26602 30852 26608 30864
rect 25630 30824 26608 30852
rect 25630 30821 25642 30824
rect 25584 30815 25642 30821
rect 26602 30812 26608 30824
rect 26660 30812 26666 30864
rect 25866 30784 25872 30796
rect 25332 30756 25872 30784
rect 25038 30676 25044 30728
rect 25096 30716 25102 30728
rect 25332 30725 25360 30756
rect 25866 30744 25872 30756
rect 25924 30744 25930 30796
rect 27816 30793 27844 30892
rect 27890 30880 27896 30892
rect 27948 30880 27954 30932
rect 34054 30880 34060 30932
rect 34112 30920 34118 30932
rect 36081 30923 36139 30929
rect 36081 30920 36093 30923
rect 34112 30892 36093 30920
rect 34112 30880 34118 30892
rect 36081 30889 36093 30892
rect 36127 30889 36139 30923
rect 36081 30883 36139 30889
rect 36262 30880 36268 30932
rect 36320 30920 36326 30932
rect 36541 30923 36599 30929
rect 36541 30920 36553 30923
rect 36320 30892 36553 30920
rect 36320 30880 36326 30892
rect 36541 30889 36553 30892
rect 36587 30889 36599 30923
rect 36541 30883 36599 30889
rect 37274 30880 37280 30932
rect 37332 30920 37338 30932
rect 37369 30923 37427 30929
rect 37369 30920 37381 30923
rect 37332 30892 37381 30920
rect 37332 30880 37338 30892
rect 37369 30889 37381 30892
rect 37415 30889 37427 30923
rect 37369 30883 37427 30889
rect 34514 30812 34520 30864
rect 34572 30852 34578 30864
rect 35250 30852 35256 30864
rect 34572 30824 35256 30852
rect 34572 30812 34578 30824
rect 35250 30812 35256 30824
rect 35308 30812 35314 30864
rect 27801 30787 27859 30793
rect 27801 30753 27813 30787
rect 27847 30753 27859 30787
rect 27801 30747 27859 30753
rect 35802 30744 35808 30796
rect 35860 30784 35866 30796
rect 35897 30787 35955 30793
rect 35897 30784 35909 30787
rect 35860 30756 35909 30784
rect 35860 30744 35866 30756
rect 35897 30753 35909 30756
rect 35943 30753 35955 30787
rect 36722 30784 36728 30796
rect 36683 30756 36728 30784
rect 35897 30747 35955 30753
rect 36722 30744 36728 30756
rect 36780 30744 36786 30796
rect 37185 30787 37243 30793
rect 37185 30753 37197 30787
rect 37231 30753 37243 30787
rect 37185 30747 37243 30753
rect 25317 30719 25375 30725
rect 25317 30716 25329 30719
rect 25096 30688 25329 30716
rect 25096 30676 25102 30688
rect 25317 30685 25329 30688
rect 25363 30685 25375 30719
rect 37200 30716 37228 30747
rect 25317 30679 25375 30685
rect 36372 30688 37228 30716
rect 23934 30608 23940 30660
rect 23992 30648 23998 30660
rect 24670 30648 24676 30660
rect 23992 30620 24676 30648
rect 23992 30608 23998 30620
rect 24670 30608 24676 30620
rect 24728 30608 24734 30660
rect 25332 30580 25360 30679
rect 36372 30660 36400 30688
rect 26418 30608 26424 30660
rect 26476 30648 26482 30660
rect 26602 30648 26608 30660
rect 26476 30620 26608 30648
rect 26476 30608 26482 30620
rect 26602 30608 26608 30620
rect 26660 30608 26666 30660
rect 26970 30608 26976 30660
rect 27028 30648 27034 30660
rect 27890 30648 27896 30660
rect 27028 30620 27896 30648
rect 27028 30608 27034 30620
rect 27890 30608 27896 30620
rect 27948 30608 27954 30660
rect 34054 30608 34060 30660
rect 34112 30648 34118 30660
rect 36354 30648 36360 30660
rect 34112 30620 36360 30648
rect 34112 30608 34118 30620
rect 36354 30608 36360 30620
rect 36412 30608 36418 30660
rect 26234 30580 26240 30592
rect 25332 30552 26240 30580
rect 26234 30540 26240 30552
rect 26292 30540 26298 30592
rect 26694 30580 26700 30592
rect 26655 30552 26700 30580
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 26878 30540 26884 30592
rect 26936 30580 26942 30592
rect 27985 30583 28043 30589
rect 27985 30580 27997 30583
rect 26936 30552 27997 30580
rect 26936 30540 26942 30552
rect 27985 30549 27997 30552
rect 28031 30580 28043 30583
rect 28626 30580 28632 30592
rect 28031 30552 28632 30580
rect 28031 30549 28043 30552
rect 27985 30543 28043 30549
rect 28626 30540 28632 30552
rect 28684 30540 28690 30592
rect 35434 30540 35440 30592
rect 35492 30580 35498 30592
rect 35710 30580 35716 30592
rect 35492 30552 35716 30580
rect 35492 30540 35498 30552
rect 35710 30540 35716 30552
rect 35768 30540 35774 30592
rect 35986 30540 35992 30592
rect 36044 30580 36050 30592
rect 36170 30580 36176 30592
rect 36044 30552 36176 30580
rect 36044 30540 36050 30552
rect 36170 30540 36176 30552
rect 36228 30540 36234 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 2774 30336 2780 30388
rect 2832 30376 2838 30388
rect 27338 30376 27344 30388
rect 2832 30348 27344 30376
rect 2832 30336 2838 30348
rect 27338 30336 27344 30348
rect 27396 30336 27402 30388
rect 33594 30336 33600 30388
rect 33652 30376 33658 30388
rect 34606 30376 34612 30388
rect 33652 30348 34612 30376
rect 33652 30336 33658 30348
rect 34606 30336 34612 30348
rect 34664 30336 34670 30388
rect 35897 30379 35955 30385
rect 35897 30345 35909 30379
rect 35943 30376 35955 30379
rect 36633 30379 36691 30385
rect 36633 30376 36645 30379
rect 35943 30348 36645 30376
rect 35943 30345 35955 30348
rect 35897 30339 35955 30345
rect 36633 30345 36645 30348
rect 36679 30345 36691 30379
rect 36633 30339 36691 30345
rect 1581 30311 1639 30317
rect 1581 30277 1593 30311
rect 1627 30308 1639 30311
rect 4706 30308 4712 30320
rect 1627 30280 4712 30308
rect 1627 30277 1639 30280
rect 1581 30271 1639 30277
rect 4706 30268 4712 30280
rect 4764 30268 4770 30320
rect 26418 30268 26424 30320
rect 26476 30308 26482 30320
rect 26605 30311 26663 30317
rect 26605 30308 26617 30311
rect 26476 30280 26617 30308
rect 26476 30268 26482 30280
rect 26605 30277 26617 30280
rect 26651 30277 26663 30311
rect 26605 30271 26663 30277
rect 31726 30280 37596 30308
rect 1210 30200 1216 30252
rect 1268 30240 1274 30252
rect 23382 30240 23388 30252
rect 1268 30212 23388 30240
rect 1268 30200 1274 30212
rect 23382 30200 23388 30212
rect 23440 30200 23446 30252
rect 23934 30200 23940 30252
rect 23992 30240 23998 30252
rect 24394 30240 24400 30252
rect 23992 30212 24400 30240
rect 23992 30200 23998 30212
rect 24394 30200 24400 30212
rect 24452 30200 24458 30252
rect 26234 30200 26240 30252
rect 26292 30240 26298 30252
rect 27157 30243 27215 30249
rect 27157 30240 27169 30243
rect 26292 30212 27169 30240
rect 26292 30200 26298 30212
rect 27157 30209 27169 30212
rect 27203 30209 27215 30243
rect 27157 30203 27215 30209
rect 1394 30172 1400 30184
rect 1355 30144 1400 30172
rect 1394 30132 1400 30144
rect 1452 30132 1458 30184
rect 25038 30132 25044 30184
rect 25096 30172 25102 30184
rect 25225 30175 25283 30181
rect 25225 30172 25237 30175
rect 25096 30144 25237 30172
rect 25096 30132 25102 30144
rect 25225 30141 25237 30144
rect 25271 30141 25283 30175
rect 26326 30172 26332 30184
rect 25225 30135 25283 30141
rect 25613 30144 26332 30172
rect 22370 30064 22376 30116
rect 22428 30104 22434 30116
rect 23290 30104 23296 30116
rect 22428 30076 23296 30104
rect 22428 30064 22434 30076
rect 23290 30064 23296 30076
rect 23348 30064 23354 30116
rect 23382 30064 23388 30116
rect 23440 30104 23446 30116
rect 25314 30104 25320 30116
rect 23440 30076 25320 30104
rect 23440 30064 23446 30076
rect 25314 30064 25320 30076
rect 25372 30064 25378 30116
rect 25492 30107 25550 30113
rect 25492 30073 25504 30107
rect 25538 30104 25550 30107
rect 25613 30104 25641 30144
rect 26326 30132 26332 30144
rect 26384 30132 26390 30184
rect 27424 30175 27482 30181
rect 27424 30141 27436 30175
rect 27470 30172 27482 30175
rect 28258 30172 28264 30184
rect 27470 30144 28264 30172
rect 27470 30141 27482 30144
rect 27424 30135 27482 30141
rect 28258 30132 28264 30144
rect 28316 30132 28322 30184
rect 28350 30132 28356 30184
rect 28408 30172 28414 30184
rect 31726 30172 31754 30280
rect 34698 30200 34704 30252
rect 34756 30240 34762 30252
rect 34756 30212 36497 30240
rect 34756 30200 34762 30212
rect 35986 30172 35992 30184
rect 28408 30144 31754 30172
rect 35947 30144 35992 30172
rect 28408 30132 28414 30144
rect 35986 30132 35992 30144
rect 36044 30132 36050 30184
rect 36082 30175 36140 30181
rect 36082 30141 36094 30175
rect 36128 30141 36140 30175
rect 36082 30135 36140 30141
rect 25538 30076 25641 30104
rect 25700 30076 28994 30104
rect 25538 30073 25550 30076
rect 25492 30067 25550 30073
rect 19978 29996 19984 30048
rect 20036 30036 20042 30048
rect 25700 30036 25728 30076
rect 20036 30008 25728 30036
rect 20036 29996 20042 30008
rect 28442 29996 28448 30048
rect 28500 30036 28506 30048
rect 28537 30039 28595 30045
rect 28537 30036 28549 30039
rect 28500 30008 28549 30036
rect 28500 29996 28506 30008
rect 28537 30005 28549 30008
rect 28583 30036 28595 30039
rect 28718 30036 28724 30048
rect 28583 30008 28724 30036
rect 28583 30005 28595 30008
rect 28537 29999 28595 30005
rect 28718 29996 28724 30008
rect 28776 29996 28782 30048
rect 28966 30036 28994 30076
rect 34974 30064 34980 30116
rect 35032 30104 35038 30116
rect 35897 30107 35955 30113
rect 35897 30104 35909 30107
rect 35032 30076 35909 30104
rect 35032 30064 35038 30076
rect 35897 30073 35909 30076
rect 35943 30073 35955 30107
rect 36097 30104 36125 30135
rect 36170 30132 36176 30184
rect 36228 30181 36234 30184
rect 36228 30175 36277 30181
rect 36228 30141 36231 30175
rect 36265 30141 36277 30175
rect 36354 30172 36360 30184
rect 36315 30144 36360 30172
rect 36228 30135 36277 30141
rect 36228 30132 36234 30135
rect 36354 30132 36360 30144
rect 36412 30132 36418 30184
rect 36469 30181 36497 30212
rect 37568 30181 37596 30280
rect 36454 30175 36512 30181
rect 36454 30141 36466 30175
rect 36500 30141 36512 30175
rect 36454 30135 36512 30141
rect 37553 30175 37611 30181
rect 37553 30141 37565 30175
rect 37599 30141 37611 30175
rect 37826 30172 37832 30184
rect 37787 30144 37832 30172
rect 37553 30135 37611 30141
rect 37826 30132 37832 30144
rect 37884 30132 37890 30184
rect 37921 30175 37979 30181
rect 37921 30141 37933 30175
rect 37967 30172 37979 30175
rect 38194 30172 38200 30184
rect 37967 30144 38200 30172
rect 37967 30141 37979 30144
rect 37921 30135 37979 30141
rect 38194 30132 38200 30144
rect 38252 30132 38258 30184
rect 37274 30104 37280 30116
rect 36097 30076 37280 30104
rect 35897 30067 35955 30073
rect 37274 30064 37280 30076
rect 37332 30064 37338 30116
rect 37734 30104 37740 30116
rect 37695 30076 37740 30104
rect 37734 30064 37740 30076
rect 37792 30064 37798 30116
rect 36446 30036 36452 30048
rect 28966 30008 36452 30036
rect 36446 29996 36452 30008
rect 36504 29996 36510 30048
rect 36722 29996 36728 30048
rect 36780 30036 36786 30048
rect 38105 30039 38163 30045
rect 38105 30036 38117 30039
rect 36780 30008 38117 30036
rect 36780 29996 36786 30008
rect 38105 30005 38117 30008
rect 38151 30005 38163 30039
rect 38105 29999 38163 30005
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 19242 29832 19248 29844
rect 19168 29804 19248 29832
rect 19168 29773 19196 29804
rect 19242 29792 19248 29804
rect 19300 29792 19306 29844
rect 19429 29835 19487 29841
rect 19429 29801 19441 29835
rect 19475 29832 19487 29835
rect 23934 29832 23940 29844
rect 19475 29804 23940 29832
rect 19475 29801 19487 29804
rect 19429 29795 19487 29801
rect 23934 29792 23940 29804
rect 23992 29792 23998 29844
rect 36170 29832 36176 29844
rect 24136 29804 36176 29832
rect 19153 29767 19211 29773
rect 19153 29733 19165 29767
rect 19199 29733 19211 29767
rect 24136 29764 24164 29804
rect 36170 29792 36176 29804
rect 36228 29792 36234 29844
rect 37185 29835 37243 29841
rect 36288 29804 37136 29832
rect 19153 29727 19211 29733
rect 19352 29736 24164 29764
rect 24572 29767 24630 29773
rect 17586 29656 17592 29708
rect 17644 29696 17650 29708
rect 18966 29705 18972 29708
rect 18785 29699 18843 29705
rect 18785 29696 18797 29699
rect 17644 29668 18797 29696
rect 17644 29656 17650 29668
rect 18785 29665 18797 29668
rect 18831 29665 18843 29699
rect 18785 29659 18843 29665
rect 18933 29699 18972 29705
rect 18933 29665 18945 29699
rect 18933 29659 18972 29665
rect 18966 29656 18972 29659
rect 19024 29656 19030 29708
rect 19061 29699 19119 29705
rect 19061 29665 19073 29699
rect 19107 29665 19119 29699
rect 19061 29659 19119 29665
rect 19250 29699 19308 29705
rect 19250 29665 19262 29699
rect 19296 29665 19308 29699
rect 19250 29659 19308 29665
rect 1670 29588 1676 29640
rect 1728 29628 1734 29640
rect 15286 29628 15292 29640
rect 1728 29600 15292 29628
rect 1728 29588 1734 29600
rect 15286 29588 15292 29600
rect 15344 29588 15350 29640
rect 18322 29588 18328 29640
rect 18380 29628 18386 29640
rect 19076 29628 19104 29659
rect 18380 29600 19104 29628
rect 18380 29588 18386 29600
rect 4890 29520 4896 29572
rect 4948 29560 4954 29572
rect 19260 29560 19288 29659
rect 4948 29532 19288 29560
rect 4948 29520 4954 29532
rect 18874 29452 18880 29504
rect 18932 29492 18938 29504
rect 19352 29492 19380 29736
rect 24572 29733 24584 29767
rect 24618 29764 24630 29767
rect 25222 29764 25228 29776
rect 24618 29736 25228 29764
rect 24618 29733 24630 29736
rect 24572 29727 24630 29733
rect 25222 29724 25228 29736
rect 25280 29724 25286 29776
rect 26510 29724 26516 29776
rect 26568 29764 26574 29776
rect 32950 29764 32956 29776
rect 26568 29736 32956 29764
rect 26568 29724 26574 29736
rect 32950 29724 32956 29736
rect 33008 29724 33014 29776
rect 36288 29764 36316 29804
rect 36152 29736 36316 29764
rect 20346 29656 20352 29708
rect 20404 29696 20410 29708
rect 22741 29699 22799 29705
rect 22741 29696 22753 29699
rect 20404 29668 22753 29696
rect 20404 29656 20410 29668
rect 22741 29665 22753 29668
rect 22787 29665 22799 29699
rect 22922 29696 22928 29708
rect 22883 29668 22928 29696
rect 22741 29659 22799 29665
rect 22922 29656 22928 29668
rect 22980 29656 22986 29708
rect 23201 29699 23259 29705
rect 23201 29665 23213 29699
rect 23247 29696 23259 29699
rect 24026 29696 24032 29708
rect 23247 29668 24032 29696
rect 23247 29665 23259 29668
rect 23201 29659 23259 29665
rect 24026 29656 24032 29668
rect 24084 29656 24090 29708
rect 24210 29656 24216 29708
rect 24268 29696 24274 29708
rect 24305 29699 24363 29705
rect 24305 29696 24317 29699
rect 24268 29668 24317 29696
rect 24268 29656 24274 29668
rect 24305 29665 24317 29668
rect 24351 29665 24363 29699
rect 24305 29659 24363 29665
rect 26326 29656 26332 29708
rect 26384 29696 26390 29708
rect 26421 29699 26479 29705
rect 26421 29696 26433 29699
rect 26384 29668 26433 29696
rect 26384 29656 26390 29668
rect 26421 29665 26433 29668
rect 26467 29665 26479 29699
rect 26421 29659 26479 29665
rect 26697 29699 26755 29705
rect 26697 29665 26709 29699
rect 26743 29665 26755 29699
rect 26878 29696 26884 29708
rect 26839 29668 26884 29696
rect 26697 29659 26755 29665
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 23017 29631 23075 29637
rect 23017 29628 23029 29631
rect 21508 29600 23029 29628
rect 21508 29588 21514 29600
rect 23017 29597 23029 29600
rect 23063 29597 23075 29631
rect 23017 29591 23075 29597
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 24228 29628 24256 29656
rect 26510 29628 26516 29640
rect 23624 29600 24256 29628
rect 26471 29600 26516 29628
rect 23624 29588 23630 29600
rect 26510 29588 26516 29600
rect 26568 29588 26574 29640
rect 26605 29631 26663 29637
rect 26605 29597 26617 29631
rect 26651 29628 26663 29631
rect 26712 29628 26740 29659
rect 26878 29656 26884 29668
rect 26936 29656 26942 29708
rect 27522 29656 27528 29708
rect 27580 29696 27586 29708
rect 30282 29696 30288 29708
rect 27580 29668 30288 29696
rect 27580 29656 27586 29668
rect 30282 29656 30288 29668
rect 30340 29656 30346 29708
rect 35345 29699 35403 29705
rect 35345 29665 35357 29699
rect 35391 29696 35403 29699
rect 35802 29696 35808 29708
rect 35391 29668 35808 29696
rect 35391 29665 35403 29668
rect 35345 29659 35403 29665
rect 35802 29656 35808 29668
rect 35860 29656 35866 29708
rect 36152 29705 36180 29736
rect 36354 29724 36360 29776
rect 36412 29764 36418 29776
rect 37108 29764 37136 29804
rect 37185 29801 37197 29835
rect 37231 29832 37243 29835
rect 38286 29832 38292 29844
rect 37231 29804 38292 29832
rect 37231 29801 37243 29804
rect 37185 29795 37243 29801
rect 38286 29792 38292 29804
rect 38344 29792 38350 29844
rect 37734 29764 37740 29776
rect 36412 29736 36457 29764
rect 37108 29736 37740 29764
rect 36412 29724 36418 29736
rect 37734 29724 37740 29736
rect 37792 29724 37798 29776
rect 35989 29699 36047 29705
rect 35989 29665 36001 29699
rect 36035 29665 36047 29699
rect 35989 29659 36047 29665
rect 36137 29699 36195 29705
rect 36137 29665 36149 29699
rect 36183 29665 36195 29699
rect 36137 29659 36195 29665
rect 26970 29628 26976 29640
rect 26651 29597 26676 29628
rect 26712 29600 26976 29628
rect 26605 29591 26676 29597
rect 22833 29563 22891 29569
rect 22833 29529 22845 29563
rect 22879 29560 22891 29563
rect 23106 29560 23112 29572
rect 22879 29532 23112 29560
rect 22879 29529 22891 29532
rect 22833 29523 22891 29529
rect 23106 29520 23112 29532
rect 23164 29520 23170 29572
rect 25682 29560 25688 29572
rect 25643 29532 25688 29560
rect 25682 29520 25688 29532
rect 25740 29520 25746 29572
rect 26648 29560 26676 29591
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 29270 29628 29276 29640
rect 27816 29600 29276 29628
rect 27816 29560 27844 29600
rect 29270 29588 29276 29600
rect 29328 29588 29334 29640
rect 36004 29628 36032 29659
rect 36262 29656 36268 29708
rect 36320 29696 36326 29708
rect 36320 29668 36365 29696
rect 36320 29656 36326 29668
rect 36446 29656 36452 29708
rect 36504 29705 36510 29708
rect 36504 29696 36512 29705
rect 37366 29696 37372 29708
rect 36504 29668 36549 29696
rect 37327 29668 37372 29696
rect 36504 29659 36512 29668
rect 36504 29656 36510 29659
rect 37366 29656 37372 29668
rect 37424 29656 37430 29708
rect 37182 29628 37188 29640
rect 36004 29600 37188 29628
rect 37182 29588 37188 29600
rect 37240 29588 37246 29640
rect 31110 29560 31116 29572
rect 25792 29532 26372 29560
rect 26648 29532 27844 29560
rect 28966 29532 31116 29560
rect 18932 29464 19380 29492
rect 22557 29495 22615 29501
rect 18932 29452 18938 29464
rect 22557 29461 22569 29495
rect 22603 29492 22615 29495
rect 22922 29492 22928 29504
rect 22603 29464 22928 29492
rect 22603 29461 22615 29464
rect 22557 29455 22615 29461
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 23934 29452 23940 29504
rect 23992 29492 23998 29504
rect 25792 29492 25820 29532
rect 26234 29492 26240 29504
rect 23992 29464 25820 29492
rect 26195 29464 26240 29492
rect 23992 29452 23998 29464
rect 26234 29452 26240 29464
rect 26292 29452 26298 29504
rect 26344 29492 26372 29532
rect 28966 29492 28994 29532
rect 31110 29520 31116 29532
rect 31168 29520 31174 29572
rect 34606 29520 34612 29572
rect 34664 29560 34670 29572
rect 34974 29560 34980 29572
rect 34664 29532 34980 29560
rect 34664 29520 34670 29532
rect 34974 29520 34980 29532
rect 35032 29520 35038 29572
rect 35434 29520 35440 29572
rect 35492 29560 35498 29572
rect 36633 29563 36691 29569
rect 36633 29560 36645 29563
rect 35492 29532 36645 29560
rect 35492 29520 35498 29532
rect 36633 29529 36645 29532
rect 36679 29529 36691 29563
rect 36633 29523 36691 29529
rect 26344 29464 28994 29492
rect 32306 29452 32312 29504
rect 32364 29492 32370 29504
rect 35529 29495 35587 29501
rect 35529 29492 35541 29495
rect 32364 29464 35541 29492
rect 32364 29452 32370 29464
rect 35529 29461 35541 29464
rect 35575 29461 35587 29495
rect 35529 29455 35587 29461
rect 35986 29452 35992 29504
rect 36044 29492 36050 29504
rect 38746 29492 38752 29504
rect 36044 29464 38752 29492
rect 36044 29452 36050 29464
rect 38746 29452 38752 29464
rect 38804 29452 38810 29504
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1581 29291 1639 29297
rect 1581 29257 1593 29291
rect 1627 29288 1639 29291
rect 2682 29288 2688 29300
rect 1627 29260 2688 29288
rect 1627 29257 1639 29260
rect 1581 29251 1639 29257
rect 2682 29248 2688 29260
rect 2740 29248 2746 29300
rect 18874 29288 18880 29300
rect 9646 29260 18880 29288
rect 9646 29152 9674 29260
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 20254 29248 20260 29300
rect 20312 29288 20318 29300
rect 20312 29260 24072 29288
rect 20312 29248 20318 29260
rect 23934 29220 23940 29232
rect 6886 29124 9674 29152
rect 18524 29192 23940 29220
rect 1394 29084 1400 29096
rect 1355 29056 1400 29084
rect 1394 29044 1400 29056
rect 1452 29044 1458 29096
rect 6546 28976 6552 29028
rect 6604 29016 6610 29028
rect 6886 29016 6914 29124
rect 17402 29044 17408 29096
rect 17460 29084 17466 29096
rect 18524 29093 18552 29192
rect 23934 29180 23940 29192
rect 23992 29180 23998 29232
rect 22554 29152 22560 29164
rect 22388 29124 22560 29152
rect 18424 29087 18482 29093
rect 18424 29084 18436 29087
rect 17460 29056 18436 29084
rect 17460 29044 17466 29056
rect 18424 29053 18436 29056
rect 18470 29053 18482 29087
rect 18424 29047 18482 29053
rect 18510 29087 18568 29093
rect 18510 29053 18522 29087
rect 18556 29053 18568 29087
rect 18510 29047 18568 29053
rect 18874 29044 18880 29096
rect 18932 29093 18938 29096
rect 22388 29093 22416 29124
rect 22554 29112 22560 29124
rect 22612 29112 22618 29164
rect 23290 29112 23296 29164
rect 23348 29152 23354 29164
rect 24044 29161 24072 29260
rect 26510 29248 26516 29300
rect 26568 29288 26574 29300
rect 26970 29288 26976 29300
rect 26568 29260 26976 29288
rect 26568 29248 26574 29260
rect 26970 29248 26976 29260
rect 27028 29248 27034 29300
rect 37277 29291 37335 29297
rect 27080 29260 27953 29288
rect 24302 29180 24308 29232
rect 24360 29220 24366 29232
rect 27080 29220 27108 29260
rect 24360 29192 27108 29220
rect 24360 29180 24366 29192
rect 27522 29180 27528 29232
rect 27580 29220 27586 29232
rect 27709 29223 27767 29229
rect 27709 29220 27721 29223
rect 27580 29192 27721 29220
rect 27580 29180 27586 29192
rect 27709 29189 27721 29192
rect 27755 29189 27767 29223
rect 27709 29183 27767 29189
rect 23569 29155 23627 29161
rect 23569 29152 23581 29155
rect 23348 29124 23581 29152
rect 23348 29112 23354 29124
rect 23569 29121 23581 29124
rect 23615 29121 23627 29155
rect 23569 29115 23627 29121
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29121 24087 29155
rect 24578 29152 24584 29164
rect 24029 29115 24087 29121
rect 24136 29124 24584 29152
rect 18932 29084 18940 29093
rect 22373 29087 22431 29093
rect 18932 29056 18977 29084
rect 18932 29047 18940 29056
rect 22373 29053 22385 29087
rect 22419 29053 22431 29087
rect 22373 29047 22431 29053
rect 18932 29044 18938 29047
rect 22462 29044 22468 29096
rect 22520 29084 22526 29096
rect 22649 29087 22707 29093
rect 22520 29056 22565 29084
rect 22520 29044 22526 29056
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 23474 29084 23480 29096
rect 22695 29056 23480 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 23474 29044 23480 29056
rect 23532 29044 23538 29096
rect 23753 29087 23811 29093
rect 23753 29053 23765 29087
rect 23799 29053 23811 29087
rect 23753 29047 23811 29053
rect 23845 29087 23903 29093
rect 23845 29053 23857 29087
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 23937 29087 23995 29093
rect 23937 29053 23949 29087
rect 23983 29084 23995 29087
rect 24136 29084 24164 29124
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 26970 29112 26976 29164
rect 27028 29152 27034 29164
rect 27925 29161 27953 29260
rect 36096 29260 36492 29288
rect 31846 29180 31852 29232
rect 31904 29220 31910 29232
rect 35066 29220 35072 29232
rect 31904 29192 35072 29220
rect 31904 29180 31910 29192
rect 35066 29180 35072 29192
rect 35124 29180 35130 29232
rect 35986 29220 35992 29232
rect 35268 29192 35992 29220
rect 27433 29155 27491 29161
rect 27433 29152 27445 29155
rect 27028 29124 27445 29152
rect 27028 29112 27034 29124
rect 27433 29121 27445 29124
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 27910 29155 27968 29161
rect 27910 29121 27922 29155
rect 27956 29121 27968 29155
rect 31202 29152 31208 29164
rect 27910 29115 27968 29121
rect 28000 29124 31208 29152
rect 23983 29056 24164 29084
rect 23983 29053 23995 29056
rect 23937 29047 23995 29053
rect 6604 28988 6914 29016
rect 6604 28976 6610 28988
rect 18322 28976 18328 29028
rect 18380 29016 18386 29028
rect 18693 29019 18751 29025
rect 18693 29016 18705 29019
rect 18380 28988 18705 29016
rect 18380 28976 18386 28988
rect 18693 28985 18705 28988
rect 18739 28985 18751 29019
rect 18693 28979 18751 28985
rect 18785 29019 18843 29025
rect 18785 28985 18797 29019
rect 18831 29016 18843 29019
rect 19150 29016 19156 29028
rect 18831 28988 19156 29016
rect 18831 28985 18843 28988
rect 18785 28979 18843 28985
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 20714 28976 20720 29028
rect 20772 29016 20778 29028
rect 23768 29016 23796 29047
rect 20772 28988 23796 29016
rect 23860 29016 23888 29047
rect 24210 29044 24216 29096
rect 24268 29084 24274 29096
rect 27522 29084 27528 29096
rect 24268 29056 24313 29084
rect 25148 29056 27528 29084
rect 24268 29044 24274 29056
rect 25148 29016 25176 29056
rect 27522 29044 27528 29056
rect 27580 29044 27586 29096
rect 27617 29087 27675 29093
rect 27617 29053 27629 29087
rect 27663 29084 27675 29087
rect 27801 29087 27859 29093
rect 27663 29056 27752 29084
rect 27663 29053 27675 29056
rect 27617 29047 27675 29053
rect 23860 28988 25176 29016
rect 25225 29019 25283 29025
rect 20772 28976 20778 28988
rect 25225 28985 25237 29019
rect 25271 29016 25283 29019
rect 25314 29016 25320 29028
rect 25271 28988 25320 29016
rect 25271 28985 25283 28988
rect 25225 28979 25283 28985
rect 25314 28976 25320 28988
rect 25372 28976 25378 29028
rect 26973 29019 27031 29025
rect 26973 28985 26985 29019
rect 27019 29016 27031 29019
rect 27062 29016 27068 29028
rect 27019 28988 27068 29016
rect 27019 28985 27031 28988
rect 26973 28979 27031 28985
rect 27062 28976 27068 28988
rect 27120 29016 27126 29028
rect 27338 29016 27344 29028
rect 27120 28988 27344 29016
rect 27120 28976 27126 28988
rect 27338 28976 27344 28988
rect 27396 28976 27402 29028
rect 27724 29016 27752 29056
rect 27801 29053 27813 29087
rect 27847 29084 27859 29087
rect 28000 29084 28028 29124
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 35158 29152 35164 29164
rect 34572 29124 35164 29152
rect 34572 29112 34578 29124
rect 35158 29112 35164 29124
rect 35216 29112 35222 29164
rect 27847 29056 28028 29084
rect 28089 29087 28147 29093
rect 27847 29053 27859 29056
rect 27801 29047 27859 29053
rect 28089 29053 28101 29087
rect 28135 29084 28147 29087
rect 28626 29084 28632 29096
rect 28135 29056 28632 29084
rect 28135 29053 28147 29056
rect 28089 29047 28147 29053
rect 28626 29044 28632 29056
rect 28684 29044 28690 29096
rect 28350 29016 28356 29028
rect 27724 28988 28356 29016
rect 28350 28976 28356 28988
rect 28408 28976 28414 29028
rect 19061 28951 19119 28957
rect 19061 28917 19073 28951
rect 19107 28948 19119 28951
rect 22462 28948 22468 28960
rect 19107 28920 22468 28948
rect 19107 28917 19119 28920
rect 19061 28911 19119 28917
rect 22462 28908 22468 28920
rect 22520 28908 22526 28960
rect 22830 28908 22836 28960
rect 22888 28948 22894 28960
rect 22888 28920 22933 28948
rect 22888 28908 22894 28920
rect 24026 28908 24032 28960
rect 24084 28948 24090 28960
rect 24210 28948 24216 28960
rect 24084 28920 24216 28948
rect 24084 28908 24090 28920
rect 24210 28908 24216 28920
rect 24268 28908 24274 28960
rect 27706 28908 27712 28960
rect 27764 28948 27770 28960
rect 35268 28948 35296 29192
rect 35986 29180 35992 29192
rect 36044 29180 36050 29232
rect 36096 29152 36124 29260
rect 36464 29220 36492 29260
rect 37277 29257 37289 29291
rect 37323 29288 37335 29291
rect 37550 29288 37556 29300
rect 37323 29260 37556 29288
rect 37323 29257 37335 29260
rect 37277 29251 37335 29257
rect 37550 29248 37556 29260
rect 37608 29248 37614 29300
rect 37918 29288 37924 29300
rect 37879 29260 37924 29288
rect 37918 29248 37924 29260
rect 37976 29248 37982 29300
rect 37458 29220 37464 29232
rect 36464 29192 37464 29220
rect 37458 29180 37464 29192
rect 37516 29180 37522 29232
rect 35912 29124 36124 29152
rect 35912 29093 35940 29124
rect 36170 29112 36176 29164
rect 36228 29112 36234 29164
rect 35897 29087 35955 29093
rect 35897 29053 35909 29087
rect 35943 29053 35955 29087
rect 35897 29047 35955 29053
rect 35986 29044 35992 29096
rect 36044 29084 36050 29096
rect 36188 29084 36216 29112
rect 36362 29087 36420 29093
rect 36362 29084 36374 29087
rect 36044 29056 36089 29084
rect 36188 29056 36374 29084
rect 36044 29044 36050 29056
rect 36362 29053 36374 29056
rect 36408 29053 36420 29087
rect 37458 29084 37464 29096
rect 37419 29056 37464 29084
rect 36362 29047 36420 29053
rect 37458 29044 37464 29056
rect 37516 29044 37522 29096
rect 38102 29084 38108 29096
rect 38063 29056 38108 29084
rect 38102 29044 38108 29056
rect 38160 29044 38166 29096
rect 36170 29016 36176 29028
rect 36131 28988 36176 29016
rect 36170 28976 36176 28988
rect 36228 28976 36234 29028
rect 36265 29019 36323 29025
rect 36265 28985 36277 29019
rect 36311 29016 36323 29019
rect 36446 29016 36452 29028
rect 36311 28988 36452 29016
rect 36311 28985 36323 28988
rect 36265 28979 36323 28985
rect 36446 28976 36452 28988
rect 36504 28976 36510 29028
rect 27764 28920 35296 28948
rect 27764 28908 27770 28920
rect 35802 28908 35808 28960
rect 35860 28948 35866 28960
rect 36541 28951 36599 28957
rect 36541 28948 36553 28951
rect 35860 28920 36553 28948
rect 35860 28908 35866 28920
rect 36541 28917 36553 28920
rect 36587 28917 36599 28951
rect 36541 28911 36599 28917
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 19337 28747 19395 28753
rect 9646 28716 19196 28744
rect 9646 28676 9674 28716
rect 6886 28648 9674 28676
rect 1670 28608 1676 28620
rect 1631 28580 1676 28608
rect 1670 28568 1676 28580
rect 1728 28568 1734 28620
rect 2958 28568 2964 28620
rect 3016 28608 3022 28620
rect 6886 28608 6914 28648
rect 18322 28636 18328 28688
rect 18380 28676 18386 28688
rect 18969 28679 19027 28685
rect 18969 28676 18981 28679
rect 18380 28648 18981 28676
rect 18380 28636 18386 28648
rect 18969 28645 18981 28648
rect 19015 28645 19027 28679
rect 18969 28639 19027 28645
rect 3016 28580 6914 28608
rect 3016 28568 3022 28580
rect 17218 28568 17224 28620
rect 17276 28608 17282 28620
rect 19168 28617 19196 28716
rect 19337 28713 19349 28747
rect 19383 28744 19395 28747
rect 19978 28744 19984 28756
rect 19383 28716 19984 28744
rect 19383 28713 19395 28716
rect 19337 28707 19395 28713
rect 19978 28704 19984 28716
rect 20036 28704 20042 28756
rect 20162 28704 20168 28756
rect 20220 28744 20226 28756
rect 20441 28747 20499 28753
rect 20220 28716 20392 28744
rect 20220 28704 20226 28716
rect 19242 28636 19248 28688
rect 19300 28676 19306 28688
rect 20073 28679 20131 28685
rect 20073 28676 20085 28679
rect 19300 28648 20085 28676
rect 19300 28636 19306 28648
rect 20073 28645 20085 28648
rect 20119 28645 20131 28679
rect 20364 28676 20392 28716
rect 20441 28713 20453 28747
rect 20487 28744 20499 28747
rect 22370 28744 22376 28756
rect 20487 28716 22376 28744
rect 20487 28713 20499 28716
rect 20441 28707 20499 28713
rect 22370 28704 22376 28716
rect 22428 28704 22434 28756
rect 22646 28704 22652 28756
rect 22704 28744 22710 28756
rect 23014 28744 23020 28756
rect 22704 28716 23020 28744
rect 22704 28704 22710 28716
rect 23014 28704 23020 28716
rect 23072 28704 23078 28756
rect 23382 28704 23388 28756
rect 23440 28744 23446 28756
rect 26326 28744 26332 28756
rect 23440 28716 26332 28744
rect 23440 28704 23446 28716
rect 26326 28704 26332 28716
rect 26384 28704 26390 28756
rect 27154 28704 27160 28756
rect 27212 28744 27218 28756
rect 33042 28744 33048 28756
rect 27212 28716 33048 28744
rect 27212 28704 27218 28716
rect 33042 28704 33048 28716
rect 33100 28704 33106 28756
rect 35894 28704 35900 28756
rect 35952 28744 35958 28756
rect 36722 28744 36728 28756
rect 35952 28716 36728 28744
rect 35952 28704 35958 28716
rect 36722 28704 36728 28716
rect 36780 28704 36786 28756
rect 37182 28704 37188 28756
rect 37240 28744 37246 28756
rect 37369 28747 37427 28753
rect 37240 28704 37274 28744
rect 37369 28713 37381 28747
rect 37415 28713 37427 28747
rect 37369 28707 37427 28713
rect 32306 28676 32312 28688
rect 20364 28648 32312 28676
rect 20073 28639 20131 28645
rect 32306 28636 32312 28648
rect 32364 28636 32370 28688
rect 35066 28636 35072 28688
rect 35124 28676 35130 28688
rect 36078 28676 36084 28688
rect 35124 28648 36084 28676
rect 35124 28636 35130 28648
rect 36078 28636 36084 28648
rect 36136 28636 36142 28688
rect 36262 28676 36268 28688
rect 36223 28648 36268 28676
rect 36262 28636 36268 28648
rect 36320 28636 36326 28688
rect 37246 28676 37274 28704
rect 37384 28676 37412 28707
rect 37246 28648 37412 28676
rect 18682 28611 18740 28617
rect 18682 28608 18694 28611
rect 17276 28580 18694 28608
rect 17276 28568 17282 28580
rect 18682 28577 18694 28580
rect 18728 28577 18740 28611
rect 18682 28571 18740 28577
rect 18786 28611 18844 28617
rect 18786 28577 18798 28611
rect 18832 28577 18844 28611
rect 18786 28571 18844 28577
rect 19061 28611 19119 28617
rect 19061 28577 19073 28611
rect 19107 28577 19119 28611
rect 19061 28571 19119 28577
rect 19158 28611 19216 28617
rect 19158 28577 19170 28611
rect 19204 28577 19216 28611
rect 19794 28608 19800 28620
rect 19755 28580 19800 28608
rect 19158 28571 19216 28577
rect 1394 28540 1400 28552
rect 1355 28512 1400 28540
rect 1394 28500 1400 28512
rect 1452 28500 1458 28552
rect 18598 28432 18604 28484
rect 18656 28472 18662 28484
rect 18800 28472 18828 28571
rect 19076 28540 19104 28571
rect 19794 28568 19800 28580
rect 19852 28568 19858 28620
rect 19978 28617 19984 28620
rect 19945 28611 19984 28617
rect 19945 28577 19957 28611
rect 19945 28571 19984 28577
rect 19978 28568 19984 28571
rect 20036 28568 20042 28620
rect 20165 28611 20223 28617
rect 20165 28577 20177 28611
rect 20211 28577 20223 28611
rect 20165 28571 20223 28577
rect 20262 28611 20320 28617
rect 20262 28577 20274 28611
rect 20308 28577 20320 28611
rect 22554 28608 22560 28620
rect 22515 28580 22560 28608
rect 20262 28571 20320 28577
rect 20180 28540 20208 28571
rect 19076 28512 20208 28540
rect 18656 28444 18828 28472
rect 18656 28432 18662 28444
rect 19212 28416 19240 28512
rect 19610 28432 19616 28484
rect 19668 28472 19674 28484
rect 20272 28472 20300 28571
rect 22554 28568 22560 28580
rect 22612 28568 22618 28620
rect 22813 28611 22871 28617
rect 22813 28608 22825 28611
rect 22664 28580 22825 28608
rect 22462 28500 22468 28552
rect 22520 28540 22526 28552
rect 22664 28540 22692 28580
rect 22813 28577 22825 28580
rect 22859 28577 22871 28611
rect 22813 28571 22871 28577
rect 23106 28568 23112 28620
rect 23164 28608 23170 28620
rect 23164 28580 23612 28608
rect 23164 28568 23170 28580
rect 22520 28512 22692 28540
rect 23584 28540 23612 28580
rect 25038 28568 25044 28620
rect 25096 28608 25102 28620
rect 25225 28611 25283 28617
rect 25225 28608 25237 28611
rect 25096 28580 25237 28608
rect 25096 28568 25102 28580
rect 25225 28577 25237 28580
rect 25271 28577 25283 28611
rect 25225 28571 25283 28577
rect 25492 28611 25550 28617
rect 25492 28577 25504 28611
rect 25538 28608 25550 28611
rect 35897 28611 35955 28617
rect 25538 28580 27614 28608
rect 25538 28577 25550 28580
rect 25492 28571 25550 28577
rect 27586 28540 27614 28580
rect 35897 28577 35909 28611
rect 35943 28577 35955 28611
rect 35897 28571 35955 28577
rect 35990 28611 36048 28617
rect 35990 28577 36002 28611
rect 36036 28577 36048 28611
rect 36170 28608 36176 28620
rect 36131 28580 36176 28608
rect 35990 28571 36048 28577
rect 23584 28512 25084 28540
rect 27586 28512 27660 28540
rect 22520 28500 22526 28512
rect 25056 28484 25084 28512
rect 19668 28444 20300 28472
rect 19668 28432 19674 28444
rect 25038 28432 25044 28484
rect 25096 28432 25102 28484
rect 27522 28472 27528 28484
rect 26160 28444 27528 28472
rect 19150 28364 19156 28416
rect 19208 28376 19240 28416
rect 19208 28364 19214 28376
rect 20806 28364 20812 28416
rect 20864 28404 20870 28416
rect 23937 28407 23995 28413
rect 23937 28404 23949 28407
rect 20864 28376 23949 28404
rect 20864 28364 20870 28376
rect 23937 28373 23949 28376
rect 23983 28373 23995 28407
rect 23937 28367 23995 28373
rect 24210 28364 24216 28416
rect 24268 28404 24274 28416
rect 26160 28404 26188 28444
rect 27522 28432 27528 28444
rect 27580 28432 27586 28484
rect 27632 28472 27660 28512
rect 28258 28472 28264 28484
rect 27632 28444 28264 28472
rect 28258 28432 28264 28444
rect 28316 28432 28322 28484
rect 31938 28432 31944 28484
rect 31996 28472 32002 28484
rect 35158 28472 35164 28484
rect 31996 28444 35164 28472
rect 31996 28432 32002 28444
rect 35158 28432 35164 28444
rect 35216 28432 35222 28484
rect 35912 28472 35940 28571
rect 36004 28540 36032 28571
rect 36170 28568 36176 28580
rect 36228 28568 36234 28620
rect 36403 28611 36461 28617
rect 36403 28577 36415 28611
rect 36449 28608 36461 28611
rect 37182 28608 37188 28620
rect 36449 28580 36860 28608
rect 37143 28580 37188 28608
rect 36449 28577 36461 28580
rect 36403 28571 36461 28577
rect 36630 28540 36636 28552
rect 36004 28512 36636 28540
rect 36630 28500 36636 28512
rect 36688 28500 36694 28552
rect 36832 28540 36860 28580
rect 37182 28568 37188 28580
rect 37240 28568 37246 28620
rect 37366 28540 37372 28552
rect 36832 28512 37372 28540
rect 37366 28500 37372 28512
rect 37424 28500 37430 28552
rect 36998 28472 37004 28484
rect 35912 28444 37004 28472
rect 36998 28432 37004 28444
rect 37056 28432 37062 28484
rect 26602 28404 26608 28416
rect 24268 28376 26188 28404
rect 26515 28376 26608 28404
rect 24268 28364 24274 28376
rect 26602 28364 26608 28376
rect 26660 28404 26666 28416
rect 28994 28404 29000 28416
rect 26660 28376 29000 28404
rect 26660 28364 26666 28376
rect 28994 28364 29000 28376
rect 29052 28364 29058 28416
rect 35250 28364 35256 28416
rect 35308 28404 35314 28416
rect 36541 28407 36599 28413
rect 36541 28404 36553 28407
rect 35308 28376 36553 28404
rect 35308 28364 35314 28376
rect 36541 28373 36553 28376
rect 36587 28373 36599 28407
rect 36541 28367 36599 28373
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 2314 28160 2320 28212
rect 2372 28200 2378 28212
rect 6362 28200 6368 28212
rect 2372 28172 6368 28200
rect 2372 28160 2378 28172
rect 6362 28160 6368 28172
rect 6420 28160 6426 28212
rect 19061 28203 19119 28209
rect 19061 28169 19073 28203
rect 19107 28200 19119 28203
rect 21634 28200 21640 28212
rect 19107 28172 21640 28200
rect 19107 28169 19119 28172
rect 19061 28163 19119 28169
rect 21634 28160 21640 28172
rect 21692 28160 21698 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22152 28172 36405 28200
rect 22152 28160 22158 28172
rect 18046 28092 18052 28144
rect 18104 28132 18110 28144
rect 18104 28104 18920 28132
rect 18104 28092 18110 28104
rect 18782 28024 18788 28076
rect 18840 28024 18846 28076
rect 18892 28064 18920 28104
rect 24394 28092 24400 28144
rect 24452 28132 24458 28144
rect 27154 28132 27160 28144
rect 24452 28104 26280 28132
rect 27115 28104 27160 28132
rect 24452 28092 24458 28104
rect 26142 28064 26148 28076
rect 18892 28036 21128 28064
rect 16022 27956 16028 28008
rect 16080 27996 16086 28008
rect 18417 27999 18475 28005
rect 18417 27996 18429 27999
rect 16080 27968 18429 27996
rect 16080 27956 16086 27968
rect 18417 27965 18429 27968
rect 18463 27965 18475 27999
rect 18417 27959 18475 27965
rect 18565 27999 18623 28005
rect 18565 27965 18577 27999
rect 18611 27996 18623 27999
rect 18800 27996 18828 28024
rect 18611 27968 18828 27996
rect 18923 27999 18981 28005
rect 18611 27965 18623 27968
rect 18565 27959 18623 27965
rect 18923 27965 18935 27999
rect 18969 27996 18981 27999
rect 20993 27999 21051 28005
rect 18969 27968 19288 27996
rect 18969 27965 18981 27968
rect 18923 27959 18981 27965
rect 18322 27888 18328 27940
rect 18380 27928 18386 27940
rect 18693 27931 18751 27937
rect 18693 27928 18705 27931
rect 18380 27900 18705 27928
rect 18380 27888 18386 27900
rect 18693 27897 18705 27900
rect 18739 27897 18751 27931
rect 18693 27891 18751 27897
rect 18785 27931 18843 27937
rect 18785 27897 18797 27931
rect 18831 27928 18843 27931
rect 19150 27928 19156 27940
rect 18831 27900 19156 27928
rect 18831 27897 18843 27900
rect 18785 27891 18843 27897
rect 19150 27888 19156 27900
rect 19208 27888 19214 27940
rect 5810 27820 5816 27872
rect 5868 27860 5874 27872
rect 19260 27860 19288 27968
rect 20993 27965 21005 27999
rect 21039 27965 21051 27999
rect 21100 27996 21128 28036
rect 22066 28036 22968 28064
rect 26103 28036 26148 28064
rect 22066 27996 22094 28036
rect 21100 27968 22094 27996
rect 20993 27959 21051 27965
rect 19978 27888 19984 27940
rect 20036 27928 20042 27940
rect 20530 27928 20536 27940
rect 20036 27900 20536 27928
rect 20036 27888 20042 27900
rect 20530 27888 20536 27900
rect 20588 27888 20594 27940
rect 5868 27832 19288 27860
rect 5868 27820 5874 27832
rect 20254 27820 20260 27872
rect 20312 27860 20318 27872
rect 21008 27860 21036 27959
rect 22554 27956 22560 28008
rect 22612 27996 22618 28008
rect 22833 27999 22891 28005
rect 22833 27996 22845 27999
rect 22612 27968 22845 27996
rect 22612 27956 22618 27968
rect 22833 27965 22845 27968
rect 22879 27965 22891 27999
rect 22940 27996 22968 28036
rect 26142 28024 26148 28036
rect 26200 28024 26206 28076
rect 26252 28073 26280 28104
rect 27154 28092 27160 28104
rect 27212 28092 27218 28144
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28033 26295 28067
rect 28258 28064 28264 28076
rect 26237 28027 26295 28033
rect 27080 28036 28264 28064
rect 25961 27999 26019 28005
rect 25961 27996 25973 27999
rect 22940 27968 25973 27996
rect 22833 27959 22891 27965
rect 25961 27965 25973 27968
rect 26007 27965 26019 27999
rect 25961 27959 26019 27965
rect 26053 27999 26111 28005
rect 26053 27965 26065 27999
rect 26099 27965 26111 27999
rect 26053 27959 26111 27965
rect 21266 27937 21272 27940
rect 21260 27928 21272 27937
rect 21227 27900 21272 27928
rect 21260 27891 21272 27900
rect 21266 27888 21272 27891
rect 21324 27888 21330 27940
rect 21450 27888 21456 27940
rect 21508 27928 21514 27940
rect 22462 27928 22468 27940
rect 21508 27900 22468 27928
rect 21508 27888 21514 27900
rect 22462 27888 22468 27900
rect 22520 27928 22526 27940
rect 23106 27937 23112 27940
rect 22520 27900 23051 27928
rect 22520 27888 22526 27900
rect 21634 27860 21640 27872
rect 20312 27832 21640 27860
rect 20312 27820 20318 27832
rect 21634 27820 21640 27832
rect 21692 27820 21698 27872
rect 22370 27860 22376 27872
rect 22331 27832 22376 27860
rect 22370 27820 22376 27832
rect 22428 27820 22434 27872
rect 23023 27860 23051 27900
rect 23100 27891 23112 27937
rect 23164 27928 23170 27940
rect 23164 27900 23200 27928
rect 23106 27888 23112 27891
rect 23164 27888 23170 27900
rect 24670 27888 24676 27940
rect 24728 27928 24734 27940
rect 26068 27928 26096 27959
rect 26326 27956 26332 28008
rect 26384 27996 26390 28008
rect 26421 27999 26479 28005
rect 26421 27996 26433 27999
rect 26384 27968 26433 27996
rect 26384 27956 26390 27968
rect 26421 27965 26433 27968
rect 26467 27996 26479 27999
rect 26878 27996 26884 28008
rect 26467 27968 26884 27996
rect 26467 27965 26479 27968
rect 26421 27959 26479 27965
rect 26878 27956 26884 27968
rect 26936 27956 26942 28008
rect 27080 28005 27108 28036
rect 28258 28024 28264 28036
rect 28316 28024 28322 28076
rect 27065 27999 27123 28005
rect 27065 27965 27077 27999
rect 27111 27965 27123 27999
rect 27246 27996 27252 28008
rect 27207 27968 27252 27996
rect 27065 27959 27123 27965
rect 27246 27956 27252 27968
rect 27304 27956 27310 28008
rect 27358 27999 27416 28005
rect 27358 27996 27370 27999
rect 27356 27965 27370 27996
rect 27404 27965 27416 27999
rect 27522 27996 27528 28008
rect 27483 27968 27528 27996
rect 27356 27959 27416 27965
rect 27356 27928 27384 27959
rect 27522 27956 27528 27968
rect 27580 27956 27586 28008
rect 35894 27996 35900 28008
rect 35855 27968 35900 27996
rect 35894 27956 35900 27968
rect 35952 27956 35958 28008
rect 35990 27999 36048 28005
rect 35990 27965 36002 27999
rect 36036 27965 36048 27999
rect 36262 27996 36268 28008
rect 36223 27968 36268 27996
rect 35990 27959 36048 27965
rect 27706 27928 27712 27940
rect 24728 27900 26004 27928
rect 26068 27900 27200 27928
rect 27356 27900 27712 27928
rect 24728 27888 24734 27900
rect 24213 27863 24271 27869
rect 24213 27860 24225 27863
rect 23023 27832 24225 27860
rect 24213 27829 24225 27832
rect 24259 27829 24271 27863
rect 25774 27860 25780 27872
rect 25735 27832 25780 27860
rect 24213 27823 24271 27829
rect 25774 27820 25780 27832
rect 25832 27820 25838 27872
rect 25976 27860 26004 27900
rect 26142 27860 26148 27872
rect 25976 27832 26148 27860
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 26878 27860 26884 27872
rect 26839 27832 26884 27860
rect 26878 27820 26884 27832
rect 26936 27820 26942 27872
rect 27172 27860 27200 27900
rect 27706 27888 27712 27900
rect 27764 27888 27770 27940
rect 32674 27860 32680 27872
rect 27172 27832 32680 27860
rect 32674 27820 32680 27832
rect 32732 27820 32738 27872
rect 36004 27860 36032 27959
rect 36262 27956 36268 27968
rect 36320 27956 36326 28008
rect 36377 28005 36405 28172
rect 36722 28160 36728 28212
rect 36780 28200 36786 28212
rect 37277 28203 37335 28209
rect 37277 28200 37289 28203
rect 36780 28172 37289 28200
rect 36780 28160 36786 28172
rect 37277 28169 37289 28172
rect 37323 28169 37335 28203
rect 37277 28163 37335 28169
rect 38105 28203 38163 28209
rect 38105 28169 38117 28203
rect 38151 28200 38163 28203
rect 38470 28200 38476 28212
rect 38151 28172 38476 28200
rect 38151 28169 38163 28172
rect 38105 28163 38163 28169
rect 38470 28160 38476 28172
rect 38528 28160 38534 28212
rect 36446 28092 36452 28144
rect 36504 28132 36510 28144
rect 36541 28135 36599 28141
rect 36541 28132 36553 28135
rect 36504 28104 36553 28132
rect 36504 28092 36510 28104
rect 36541 28101 36553 28104
rect 36587 28101 36599 28135
rect 36541 28095 36599 28101
rect 36362 27999 36420 28005
rect 36362 27965 36374 27999
rect 36408 27965 36420 27999
rect 37458 27996 37464 28008
rect 37419 27968 37464 27996
rect 36362 27959 36420 27965
rect 37458 27956 37464 27968
rect 37516 27956 37522 28008
rect 37918 27996 37924 28008
rect 37879 27968 37924 27996
rect 37918 27956 37924 27968
rect 37976 27956 37982 28008
rect 36170 27928 36176 27940
rect 36131 27900 36176 27928
rect 36170 27888 36176 27900
rect 36228 27888 36234 27940
rect 36998 27860 37004 27872
rect 36004 27832 37004 27860
rect 36998 27820 37004 27832
rect 37056 27820 37062 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 2958 27656 2964 27668
rect 2792 27628 2964 27656
rect 2792 27600 2820 27628
rect 2958 27616 2964 27628
rect 3016 27616 3022 27668
rect 18322 27616 18328 27668
rect 18380 27656 18386 27668
rect 19242 27656 19248 27668
rect 18380 27628 19248 27656
rect 18380 27616 18386 27628
rect 19242 27616 19248 27628
rect 19300 27616 19306 27668
rect 19797 27659 19855 27665
rect 19797 27625 19809 27659
rect 19843 27656 19855 27659
rect 20070 27656 20076 27668
rect 19843 27628 20076 27656
rect 19843 27625 19855 27628
rect 19797 27619 19855 27625
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 20898 27656 20904 27668
rect 20539 27628 20904 27656
rect 1854 27588 1860 27600
rect 1815 27560 1860 27588
rect 1854 27548 1860 27560
rect 1912 27548 1918 27600
rect 2038 27588 2044 27600
rect 1999 27560 2044 27588
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 2774 27548 2780 27600
rect 2832 27548 2838 27600
rect 10226 27548 10232 27600
rect 10284 27588 10290 27600
rect 15286 27588 15292 27600
rect 10284 27560 15292 27588
rect 10284 27548 10290 27560
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 20539 27597 20567 27628
rect 20898 27616 20904 27628
rect 20956 27656 20962 27668
rect 22370 27656 22376 27668
rect 20956 27628 22376 27656
rect 20956 27616 20962 27628
rect 22370 27616 22376 27628
rect 22428 27616 22434 27668
rect 27062 27656 27068 27668
rect 22480 27628 27068 27656
rect 20524 27591 20582 27597
rect 20524 27557 20536 27591
rect 20570 27557 20582 27591
rect 20524 27551 20582 27557
rect 20622 27548 20628 27600
rect 20680 27588 20686 27600
rect 22480 27588 22508 27628
rect 27062 27616 27068 27628
rect 27120 27616 27126 27668
rect 27706 27616 27712 27668
rect 27764 27656 27770 27668
rect 31662 27656 31668 27668
rect 27764 27628 31668 27656
rect 27764 27616 27770 27628
rect 31662 27616 31668 27628
rect 31720 27616 31726 27668
rect 36173 27659 36231 27665
rect 36173 27625 36185 27659
rect 36219 27656 36231 27659
rect 36262 27656 36268 27668
rect 36219 27628 36268 27656
rect 36219 27625 36231 27628
rect 36173 27619 36231 27625
rect 36262 27616 36268 27628
rect 36320 27616 36326 27668
rect 20680 27560 22508 27588
rect 20680 27548 20686 27560
rect 22646 27548 22652 27600
rect 22704 27588 22710 27600
rect 22802 27591 22860 27597
rect 22802 27588 22814 27591
rect 22704 27560 22814 27588
rect 22704 27548 22710 27560
rect 22802 27557 22814 27560
rect 22848 27557 22860 27591
rect 22802 27551 22860 27557
rect 24210 27548 24216 27600
rect 24268 27588 24274 27600
rect 24397 27591 24455 27597
rect 24397 27588 24409 27591
rect 24268 27560 24409 27588
rect 24268 27548 24274 27560
rect 24397 27557 24409 27560
rect 24443 27557 24455 27591
rect 24397 27551 24455 27557
rect 24486 27548 24492 27600
rect 24544 27588 24550 27600
rect 24544 27560 26096 27588
rect 24544 27548 24550 27560
rect 2222 27480 2228 27532
rect 2280 27520 2286 27532
rect 6270 27520 6276 27532
rect 2280 27492 6276 27520
rect 2280 27480 2286 27492
rect 6270 27480 6276 27492
rect 6328 27480 6334 27532
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 14918 27520 14924 27532
rect 8168 27492 14924 27520
rect 8168 27480 8174 27492
rect 14918 27480 14924 27492
rect 14976 27480 14982 27532
rect 19429 27523 19487 27529
rect 19429 27489 19441 27523
rect 19475 27520 19487 27523
rect 20806 27520 20812 27532
rect 19475 27492 20812 27520
rect 19475 27489 19487 27492
rect 19429 27483 19487 27489
rect 20806 27480 20812 27492
rect 20864 27480 20870 27532
rect 22094 27480 22100 27532
rect 22152 27520 22158 27532
rect 24736 27523 24794 27529
rect 24736 27520 24748 27523
rect 22152 27492 24748 27520
rect 22152 27480 22158 27492
rect 24736 27489 24748 27492
rect 24782 27489 24794 27523
rect 24736 27483 24794 27489
rect 25777 27523 25835 27529
rect 25777 27489 25789 27523
rect 25823 27489 25835 27523
rect 25958 27520 25964 27532
rect 25919 27492 25964 27520
rect 25777 27483 25835 27489
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19536 27384 19564 27415
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20254 27452 20260 27464
rect 20036 27424 20260 27452
rect 20036 27412 20042 27424
rect 20254 27412 20260 27424
rect 20312 27412 20318 27464
rect 21634 27412 21640 27464
rect 21692 27452 21698 27464
rect 22557 27455 22615 27461
rect 22557 27452 22569 27455
rect 21692 27424 22569 27452
rect 21692 27412 21698 27424
rect 22557 27421 22569 27424
rect 22603 27421 22615 27455
rect 22557 27415 22615 27421
rect 24578 27412 24584 27464
rect 24636 27452 24642 27464
rect 25792 27452 25820 27483
rect 25958 27480 25964 27492
rect 26016 27480 26022 27532
rect 26068 27529 26096 27560
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 31018 27588 31024 27600
rect 26200 27560 31024 27588
rect 26200 27548 26206 27560
rect 31018 27548 31024 27560
rect 31076 27548 31082 27600
rect 26053 27523 26111 27529
rect 26053 27489 26065 27523
rect 26099 27489 26111 27523
rect 26053 27483 26111 27489
rect 26237 27523 26295 27529
rect 26237 27489 26249 27523
rect 26283 27520 26295 27523
rect 26326 27520 26332 27532
rect 26283 27492 26332 27520
rect 26283 27489 26295 27492
rect 26237 27483 26295 27489
rect 26326 27480 26332 27492
rect 26384 27480 26390 27532
rect 26697 27523 26755 27529
rect 26697 27489 26709 27523
rect 26743 27489 26755 27523
rect 26697 27483 26755 27489
rect 24636 27424 25820 27452
rect 24636 27412 24642 27424
rect 26142 27412 26148 27464
rect 26200 27452 26206 27464
rect 26712 27452 26740 27483
rect 35894 27480 35900 27532
rect 35952 27520 35958 27532
rect 35989 27523 36047 27529
rect 35989 27520 36001 27523
rect 35952 27492 36001 27520
rect 35952 27480 35958 27492
rect 35989 27489 36001 27492
rect 36035 27520 36047 27523
rect 36354 27520 36360 27532
rect 36035 27492 36360 27520
rect 36035 27489 36047 27492
rect 35989 27483 36047 27489
rect 36354 27480 36360 27492
rect 36412 27480 36418 27532
rect 26200 27424 26740 27452
rect 26200 27412 26206 27424
rect 26878 27412 26884 27464
rect 26936 27452 26942 27464
rect 27062 27452 27068 27464
rect 26936 27424 27068 27452
rect 26936 27412 26942 27424
rect 27062 27412 27068 27424
rect 27120 27412 27126 27464
rect 19536 27356 20305 27384
rect 2130 27276 2136 27328
rect 2188 27316 2194 27328
rect 2406 27316 2412 27328
rect 2188 27288 2412 27316
rect 2188 27276 2194 27288
rect 2406 27276 2412 27288
rect 2464 27276 2470 27328
rect 19610 27316 19616 27328
rect 19571 27288 19616 27316
rect 19610 27276 19616 27288
rect 19668 27276 19674 27328
rect 20277 27316 20305 27356
rect 23566 27344 23572 27396
rect 23624 27384 23630 27396
rect 25593 27387 25651 27393
rect 25593 27384 25605 27387
rect 23624 27356 25605 27384
rect 23624 27344 23630 27356
rect 25593 27353 25605 27356
rect 25639 27353 25651 27387
rect 25593 27347 25651 27353
rect 25869 27387 25927 27393
rect 25869 27353 25881 27387
rect 25915 27384 25927 27387
rect 33962 27384 33968 27396
rect 25915 27356 33968 27384
rect 25915 27353 25927 27356
rect 25869 27347 25927 27353
rect 33962 27344 33968 27356
rect 34020 27344 34026 27396
rect 21450 27316 21456 27328
rect 20277 27288 21456 27316
rect 21450 27276 21456 27288
rect 21508 27276 21514 27328
rect 21634 27316 21640 27328
rect 21595 27288 21640 27316
rect 21634 27276 21640 27288
rect 21692 27276 21698 27328
rect 22462 27276 22468 27328
rect 22520 27316 22526 27328
rect 22830 27316 22836 27328
rect 22520 27288 22836 27316
rect 22520 27276 22526 27288
rect 22830 27276 22836 27288
rect 22888 27276 22894 27328
rect 23934 27316 23940 27328
rect 23895 27288 23940 27316
rect 23934 27276 23940 27288
rect 23992 27276 23998 27328
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 24535 27319 24593 27325
rect 24535 27316 24547 27319
rect 24176 27288 24547 27316
rect 24176 27276 24182 27288
rect 24535 27285 24547 27288
rect 24581 27285 24593 27319
rect 24670 27316 24676 27328
rect 24631 27288 24676 27316
rect 24535 27279 24593 27285
rect 24670 27276 24676 27288
rect 24728 27276 24734 27328
rect 25038 27316 25044 27328
rect 24999 27288 25044 27316
rect 25038 27276 25044 27288
rect 25096 27276 25102 27328
rect 25314 27276 25320 27328
rect 25372 27316 25378 27328
rect 26142 27316 26148 27328
rect 25372 27288 26148 27316
rect 25372 27276 25378 27288
rect 26142 27276 26148 27288
rect 26200 27276 26206 27328
rect 26878 27316 26884 27328
rect 26839 27288 26884 27316
rect 26878 27276 26884 27288
rect 26936 27276 26942 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 22922 27112 22928 27124
rect 21600 27084 22928 27112
rect 21600 27072 21606 27084
rect 22922 27072 22928 27084
rect 22980 27072 22986 27124
rect 25222 27072 25228 27124
rect 25280 27112 25286 27124
rect 25866 27112 25872 27124
rect 25280 27084 25872 27112
rect 25280 27072 25286 27084
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 36078 27072 36084 27124
rect 36136 27112 36142 27124
rect 37461 27115 37519 27121
rect 37461 27112 37473 27115
rect 36136 27084 37473 27112
rect 36136 27072 36142 27084
rect 37461 27081 37473 27084
rect 37507 27081 37519 27115
rect 37461 27075 37519 27081
rect 37826 27072 37832 27124
rect 37884 27112 37890 27124
rect 38105 27115 38163 27121
rect 38105 27112 38117 27115
rect 37884 27084 38117 27112
rect 37884 27072 37890 27084
rect 38105 27081 38117 27084
rect 38151 27081 38163 27115
rect 38105 27075 38163 27081
rect 2041 27047 2099 27053
rect 2041 27013 2053 27047
rect 2087 27044 2099 27047
rect 2682 27044 2688 27056
rect 2087 27016 2688 27044
rect 2087 27013 2099 27016
rect 2041 27007 2099 27013
rect 2682 27004 2688 27016
rect 2740 27004 2746 27056
rect 21361 27047 21419 27053
rect 21361 27013 21373 27047
rect 21407 27013 21419 27047
rect 21361 27007 21419 27013
rect 19978 26976 19984 26988
rect 19939 26948 19984 26976
rect 19978 26936 19984 26948
rect 20036 26936 20042 26988
rect 21376 26976 21404 27007
rect 21450 27004 21456 27056
rect 21508 27044 21514 27056
rect 21726 27044 21732 27056
rect 21508 27016 21732 27044
rect 21508 27004 21514 27016
rect 21726 27004 21732 27016
rect 21784 27004 21790 27056
rect 23474 27004 23480 27056
rect 23532 27044 23538 27056
rect 23532 27016 25728 27044
rect 23532 27004 23538 27016
rect 25590 26976 25596 26988
rect 21376 26948 21956 26976
rect 19996 26908 20024 26936
rect 20806 26908 20812 26920
rect 19996 26880 20812 26908
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 21818 26908 21824 26920
rect 21779 26880 21824 26908
rect 21818 26868 21824 26880
rect 21876 26868 21882 26920
rect 21928 26908 21956 26948
rect 23308 26948 25452 26976
rect 25551 26948 25596 26976
rect 22094 26917 22100 26920
rect 22088 26908 22100 26917
rect 21928 26880 22100 26908
rect 22088 26871 22100 26880
rect 22152 26908 22158 26920
rect 22152 26880 22236 26908
rect 22094 26868 22100 26871
rect 22152 26868 22158 26880
rect 22370 26868 22376 26920
rect 22428 26908 22434 26920
rect 23308 26908 23336 26948
rect 24670 26908 24676 26920
rect 22428 26880 23336 26908
rect 23400 26880 24676 26908
rect 22428 26868 22434 26880
rect 1854 26840 1860 26852
rect 1815 26812 1860 26840
rect 1854 26800 1860 26812
rect 1912 26800 1918 26852
rect 20070 26800 20076 26852
rect 20128 26840 20134 26852
rect 20248 26843 20306 26849
rect 20248 26840 20260 26843
rect 20128 26812 20260 26840
rect 20128 26800 20134 26812
rect 20248 26809 20260 26812
rect 20294 26840 20306 26843
rect 23400 26840 23428 26880
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 25424 26917 25452 26948
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 25700 26985 25728 27016
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26945 25743 26979
rect 30742 26976 30748 26988
rect 25685 26939 25743 26945
rect 25792 26948 30748 26976
rect 25409 26911 25467 26917
rect 25409 26877 25421 26911
rect 25455 26877 25467 26911
rect 25409 26871 25467 26877
rect 25501 26911 25559 26917
rect 25501 26877 25513 26911
rect 25547 26908 25559 26911
rect 25792 26908 25820 26948
rect 30742 26936 30748 26948
rect 30800 26936 30806 26988
rect 34606 26936 34612 26988
rect 34664 26976 34670 26988
rect 35526 26976 35532 26988
rect 34664 26948 35532 26976
rect 34664 26936 34670 26948
rect 35526 26936 35532 26948
rect 35584 26936 35590 26988
rect 25547 26880 25820 26908
rect 25869 26911 25927 26917
rect 25547 26877 25559 26880
rect 25501 26871 25559 26877
rect 25869 26877 25881 26911
rect 25915 26908 25927 26911
rect 26878 26908 26884 26920
rect 25915 26880 26884 26908
rect 25915 26877 25927 26880
rect 25869 26871 25927 26877
rect 26878 26868 26884 26880
rect 26936 26868 26942 26920
rect 37274 26908 37280 26920
rect 37235 26880 37280 26908
rect 37274 26868 37280 26880
rect 37332 26868 37338 26920
rect 37918 26908 37924 26920
rect 37879 26880 37924 26908
rect 37918 26868 37924 26880
rect 37976 26868 37982 26920
rect 20294 26812 23428 26840
rect 24121 26843 24179 26849
rect 20294 26809 20306 26812
rect 20248 26803 20306 26809
rect 24121 26809 24133 26843
rect 24167 26840 24179 26843
rect 24946 26840 24952 26852
rect 24167 26812 24952 26840
rect 24167 26809 24179 26812
rect 24121 26803 24179 26809
rect 24946 26800 24952 26812
rect 25004 26840 25010 26852
rect 25314 26840 25320 26852
rect 25004 26812 25320 26840
rect 25004 26800 25010 26812
rect 25314 26800 25320 26812
rect 25372 26800 25378 26852
rect 25958 26800 25964 26852
rect 26016 26840 26022 26852
rect 34146 26840 34152 26852
rect 26016 26812 34152 26840
rect 26016 26800 26022 26812
rect 34146 26800 34152 26812
rect 34204 26800 34210 26852
rect 35342 26800 35348 26852
rect 35400 26840 35406 26852
rect 35526 26840 35532 26852
rect 35400 26812 35532 26840
rect 35400 26800 35406 26812
rect 35526 26800 35532 26812
rect 35584 26800 35590 26852
rect 21266 26732 21272 26784
rect 21324 26772 21330 26784
rect 23201 26775 23259 26781
rect 23201 26772 23213 26775
rect 21324 26744 23213 26772
rect 21324 26732 21330 26744
rect 23201 26741 23213 26744
rect 23247 26741 23259 26775
rect 24210 26772 24216 26784
rect 24171 26744 24216 26772
rect 23201 26735 23259 26741
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 25222 26772 25228 26784
rect 25183 26744 25228 26772
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 20070 26568 20076 26580
rect 20031 26540 20076 26568
rect 20070 26528 20076 26540
rect 20128 26528 20134 26580
rect 21269 26571 21327 26577
rect 21269 26537 21281 26571
rect 21315 26568 21327 26571
rect 24118 26568 24124 26580
rect 21315 26540 24124 26568
rect 21315 26537 21327 26540
rect 21269 26531 21327 26537
rect 24118 26528 24124 26540
rect 24176 26528 24182 26580
rect 18598 26460 18604 26512
rect 18656 26500 18662 26512
rect 20254 26500 20260 26512
rect 18656 26472 20260 26500
rect 18656 26460 18662 26472
rect 20254 26460 20260 26472
rect 20312 26460 20318 26512
rect 20625 26503 20683 26509
rect 20625 26469 20637 26503
rect 20671 26500 20683 26503
rect 21634 26500 21640 26512
rect 20671 26472 21640 26500
rect 20671 26469 20683 26472
rect 20625 26463 20683 26469
rect 21634 26460 21640 26472
rect 21692 26460 21698 26512
rect 23468 26503 23526 26509
rect 23468 26469 23480 26503
rect 23514 26500 23526 26503
rect 25774 26500 25780 26512
rect 23514 26472 25780 26500
rect 23514 26469 23526 26472
rect 23468 26463 23526 26469
rect 25774 26460 25780 26472
rect 25832 26460 25838 26512
rect 7926 26392 7932 26444
rect 7984 26432 7990 26444
rect 18509 26435 18567 26441
rect 18509 26432 18521 26435
rect 7984 26404 18521 26432
rect 7984 26392 7990 26404
rect 18509 26401 18521 26404
rect 18555 26432 18567 26435
rect 18949 26435 19007 26441
rect 18949 26432 18961 26435
rect 18555 26404 18961 26432
rect 18555 26401 18567 26404
rect 18509 26395 18567 26401
rect 18949 26401 18961 26404
rect 18995 26432 19007 26435
rect 18995 26404 21128 26432
rect 18995 26401 19007 26404
rect 18949 26395 19007 26401
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 18708 26228 18736 26327
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20956 26336 21005 26364
rect 20956 26324 20962 26336
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 21100 26364 21128 26404
rect 21818 26392 21824 26444
rect 21876 26432 21882 26444
rect 21876 26404 22600 26432
rect 21876 26392 21882 26404
rect 22572 26376 22600 26404
rect 22738 26392 22744 26444
rect 22796 26432 22802 26444
rect 24394 26432 24400 26444
rect 22796 26404 24400 26432
rect 22796 26392 22802 26404
rect 24394 26392 24400 26404
rect 24452 26432 24458 26444
rect 25400 26435 25458 26441
rect 24452 26404 24532 26432
rect 24452 26392 24458 26404
rect 22186 26364 22192 26376
rect 21100 26336 22192 26364
rect 20993 26327 21051 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 22554 26324 22560 26376
rect 22612 26364 22618 26376
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22612 26336 23213 26364
rect 22612 26324 22618 26336
rect 23201 26333 23213 26336
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 20790 26299 20848 26305
rect 20790 26265 20802 26299
rect 20836 26296 20848 26299
rect 22646 26296 22652 26308
rect 20836 26268 22652 26296
rect 20836 26265 20848 26268
rect 20790 26259 20848 26265
rect 22646 26256 22652 26268
rect 22704 26256 22710 26308
rect 18874 26228 18880 26240
rect 18708 26200 18880 26228
rect 18874 26188 18880 26200
rect 18932 26228 18938 26240
rect 19978 26228 19984 26240
rect 18932 26200 19984 26228
rect 18932 26188 18938 26200
rect 19978 26188 19984 26200
rect 20036 26188 20042 26240
rect 20901 26231 20959 26237
rect 20901 26197 20913 26231
rect 20947 26228 20959 26231
rect 21266 26228 21272 26240
rect 20947 26200 21272 26228
rect 20947 26197 20959 26200
rect 20901 26191 20959 26197
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 23216 26228 23244 26327
rect 24504 26296 24532 26404
rect 25400 26401 25412 26435
rect 25446 26432 25458 26435
rect 26234 26432 26240 26444
rect 25446 26404 26240 26432
rect 25446 26401 25458 26404
rect 25400 26395 25458 26401
rect 26234 26392 26240 26404
rect 26292 26392 26298 26444
rect 25038 26364 25044 26376
rect 24688 26336 25044 26364
rect 24581 26299 24639 26305
rect 24581 26296 24593 26299
rect 24504 26268 24593 26296
rect 24581 26265 24593 26268
rect 24627 26265 24639 26299
rect 24581 26259 24639 26265
rect 24688 26228 24716 26336
rect 25038 26324 25044 26336
rect 25096 26364 25102 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 25096 26336 25145 26364
rect 25096 26324 25102 26336
rect 25133 26333 25145 26336
rect 25179 26333 25191 26367
rect 25133 26327 25191 26333
rect 26510 26296 26516 26308
rect 26471 26268 26516 26296
rect 26510 26256 26516 26268
rect 26568 26256 26574 26308
rect 23216 26200 24716 26228
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 18693 26027 18751 26033
rect 18693 25993 18705 26027
rect 18739 26024 18751 26027
rect 22281 26027 22339 26033
rect 18739 25996 22094 26024
rect 18739 25993 18751 25996
rect 18693 25987 18751 25993
rect 2041 25959 2099 25965
rect 2041 25925 2053 25959
rect 2087 25956 2099 25959
rect 2314 25956 2320 25968
rect 2087 25928 2320 25956
rect 2087 25925 2099 25928
rect 2041 25919 2099 25925
rect 2314 25916 2320 25928
rect 2372 25916 2378 25968
rect 22066 25956 22094 25996
rect 22281 25993 22293 26027
rect 22327 26024 22339 26027
rect 22646 26024 22652 26036
rect 22327 25996 22652 26024
rect 22327 25993 22339 25996
rect 22281 25987 22339 25993
rect 22646 25984 22652 25996
rect 22704 25984 22710 26036
rect 24118 26024 24124 26036
rect 22756 25996 24124 26024
rect 22756 25956 22784 25996
rect 24118 25984 24124 25996
rect 24176 25984 24182 26036
rect 24213 26027 24271 26033
rect 24213 25993 24225 26027
rect 24259 26024 24271 26027
rect 24302 26024 24308 26036
rect 24259 25996 24308 26024
rect 24259 25993 24271 25996
rect 24213 25987 24271 25993
rect 24302 25984 24308 25996
rect 24360 25984 24366 26036
rect 26605 26027 26663 26033
rect 24412 25996 26188 26024
rect 6886 25928 12434 25956
rect 22066 25928 22784 25956
rect 1854 25820 1860 25832
rect 1815 25792 1860 25820
rect 1854 25780 1860 25792
rect 1912 25780 1918 25832
rect 4798 25644 4804 25696
rect 4856 25684 4862 25696
rect 6886 25684 6914 25928
rect 12406 25888 12434 25928
rect 12406 25860 18368 25888
rect 14734 25780 14740 25832
rect 14792 25820 14798 25832
rect 18049 25823 18107 25829
rect 18049 25820 18061 25823
rect 14792 25792 18061 25820
rect 14792 25780 14798 25792
rect 18049 25789 18061 25792
rect 18095 25789 18107 25823
rect 18049 25783 18107 25789
rect 18142 25823 18200 25829
rect 18142 25789 18154 25823
rect 18188 25789 18200 25823
rect 18340 25820 18368 25860
rect 20806 25848 20812 25900
rect 20864 25888 20870 25900
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20864 25860 20913 25888
rect 20864 25848 20870 25860
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 20901 25851 20959 25857
rect 18514 25823 18572 25829
rect 18514 25820 18526 25823
rect 18340 25792 18526 25820
rect 18142 25783 18200 25789
rect 18514 25789 18526 25792
rect 18560 25789 18572 25823
rect 18514 25783 18572 25789
rect 21168 25823 21226 25829
rect 21168 25789 21180 25823
rect 21214 25820 21226 25823
rect 21634 25820 21640 25832
rect 21214 25792 21640 25820
rect 21214 25789 21226 25792
rect 21168 25783 21226 25789
rect 4856 25656 6914 25684
rect 18156 25684 18184 25783
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22554 25780 22560 25832
rect 22612 25820 22618 25832
rect 22833 25823 22891 25829
rect 22833 25820 22845 25823
rect 22612 25792 22845 25820
rect 22612 25780 22618 25792
rect 22833 25789 22845 25792
rect 22879 25789 22891 25823
rect 24412 25820 24440 25996
rect 26160 25956 26188 25996
rect 26605 25993 26617 26027
rect 26651 26024 26663 26027
rect 26786 26024 26792 26036
rect 26651 25996 26792 26024
rect 26651 25993 26663 25996
rect 26605 25987 26663 25993
rect 26786 25984 26792 25996
rect 26844 26024 26850 26036
rect 27338 26024 27344 26036
rect 26844 25996 27344 26024
rect 26844 25984 26850 25996
rect 27338 25984 27344 25996
rect 27396 25984 27402 26036
rect 36538 25984 36544 26036
rect 36596 26024 36602 26036
rect 38105 26027 38163 26033
rect 38105 26024 38117 26027
rect 36596 25996 38117 26024
rect 36596 25984 36602 25996
rect 38105 25993 38117 25996
rect 38151 25993 38163 26027
rect 38105 25987 38163 25993
rect 27522 25956 27528 25968
rect 26160 25928 27528 25956
rect 27522 25916 27528 25928
rect 27580 25916 27586 25968
rect 33226 25916 33232 25968
rect 33284 25956 33290 25968
rect 37461 25959 37519 25965
rect 37461 25956 37473 25959
rect 33284 25928 37473 25956
rect 33284 25916 33290 25928
rect 37461 25925 37473 25928
rect 37507 25925 37519 25959
rect 37461 25919 37519 25925
rect 25038 25848 25044 25900
rect 25096 25888 25102 25900
rect 25225 25891 25283 25897
rect 25225 25888 25237 25891
rect 25096 25860 25237 25888
rect 25096 25848 25102 25860
rect 25225 25857 25237 25860
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 25498 25829 25504 25832
rect 25492 25820 25504 25829
rect 22833 25783 22891 25789
rect 22940 25792 24440 25820
rect 25459 25792 25504 25820
rect 18230 25712 18236 25764
rect 18288 25752 18294 25764
rect 18325 25755 18383 25761
rect 18325 25752 18337 25755
rect 18288 25724 18337 25752
rect 18288 25712 18294 25724
rect 18325 25721 18337 25724
rect 18371 25721 18383 25755
rect 18325 25715 18383 25721
rect 18414 25712 18420 25764
rect 18472 25752 18478 25764
rect 18472 25724 18517 25752
rect 18472 25712 18478 25724
rect 22186 25712 22192 25764
rect 22244 25752 22250 25764
rect 22940 25752 22968 25792
rect 25492 25783 25504 25792
rect 25498 25780 25504 25783
rect 25556 25780 25562 25832
rect 27522 25780 27528 25832
rect 27580 25820 27586 25832
rect 27890 25820 27896 25832
rect 27580 25792 27896 25820
rect 27580 25780 27586 25792
rect 27890 25780 27896 25792
rect 27948 25780 27954 25832
rect 37274 25820 37280 25832
rect 37235 25792 37280 25820
rect 37274 25780 37280 25792
rect 37332 25780 37338 25832
rect 37918 25820 37924 25832
rect 37879 25792 37924 25820
rect 37918 25780 37924 25792
rect 37976 25780 37982 25832
rect 22244 25724 22968 25752
rect 23100 25755 23158 25761
rect 22244 25712 22250 25724
rect 23100 25721 23112 25755
rect 23146 25752 23158 25755
rect 26970 25752 26976 25764
rect 23146 25724 26976 25752
rect 23146 25721 23158 25724
rect 23100 25715 23158 25721
rect 26970 25712 26976 25724
rect 27028 25712 27034 25764
rect 23198 25684 23204 25696
rect 18156 25656 23204 25684
rect 4856 25644 4862 25656
rect 23198 25644 23204 25656
rect 23256 25644 23262 25696
rect 24118 25644 24124 25696
rect 24176 25684 24182 25696
rect 28810 25684 28816 25696
rect 24176 25656 28816 25684
rect 24176 25644 24182 25656
rect 28810 25644 28816 25656
rect 28868 25644 28874 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 18509 25483 18567 25489
rect 18028 25452 18465 25480
rect 2038 25412 2044 25424
rect 1999 25384 2044 25412
rect 2038 25372 2044 25384
rect 2096 25372 2102 25424
rect 1854 25344 1860 25356
rect 1815 25316 1860 25344
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 17770 25304 17776 25356
rect 17828 25344 17834 25356
rect 18028 25353 18056 25452
rect 18230 25412 18236 25424
rect 18191 25384 18236 25412
rect 18230 25372 18236 25384
rect 18288 25372 18294 25424
rect 18437 25412 18465 25452
rect 18509 25449 18521 25483
rect 18555 25480 18567 25483
rect 22186 25480 22192 25492
rect 18555 25452 22192 25480
rect 18555 25449 18567 25452
rect 18509 25443 18567 25449
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 23290 25480 23296 25492
rect 22756 25452 23296 25480
rect 19236 25415 19294 25421
rect 18437 25384 19095 25412
rect 17865 25347 17923 25353
rect 17865 25344 17877 25347
rect 17828 25316 17877 25344
rect 17828 25304 17834 25316
rect 17865 25313 17877 25316
rect 17911 25313 17923 25347
rect 17865 25307 17923 25313
rect 18013 25347 18071 25353
rect 18013 25313 18025 25347
rect 18059 25313 18071 25347
rect 18138 25344 18144 25356
rect 18099 25316 18144 25344
rect 18013 25307 18071 25313
rect 18138 25304 18144 25316
rect 18196 25304 18202 25356
rect 18330 25347 18388 25353
rect 18330 25313 18342 25347
rect 18376 25313 18388 25347
rect 18330 25307 18388 25313
rect 5626 25236 5632 25288
rect 5684 25276 5690 25288
rect 18345 25276 18373 25307
rect 18874 25304 18880 25356
rect 18932 25344 18938 25356
rect 18969 25347 19027 25353
rect 18969 25344 18981 25347
rect 18932 25316 18981 25344
rect 18932 25304 18938 25316
rect 18969 25313 18981 25316
rect 19015 25313 19027 25347
rect 19067 25344 19095 25384
rect 19236 25381 19248 25415
rect 19282 25412 19294 25415
rect 22756 25412 22784 25452
rect 23290 25440 23296 25452
rect 23348 25440 23354 25492
rect 23937 25483 23995 25489
rect 23937 25449 23949 25483
rect 23983 25480 23995 25483
rect 24486 25480 24492 25492
rect 23983 25452 24492 25480
rect 23983 25449 23995 25452
rect 23937 25443 23995 25449
rect 19282 25384 22784 25412
rect 22824 25415 22882 25421
rect 19282 25381 19294 25384
rect 19236 25375 19294 25381
rect 22824 25381 22836 25415
rect 22870 25412 22882 25415
rect 23566 25412 23572 25424
rect 22870 25384 23572 25412
rect 22870 25381 22882 25384
rect 22824 25375 22882 25381
rect 23566 25372 23572 25384
rect 23624 25372 23630 25424
rect 20806 25344 20812 25356
rect 19067 25316 20812 25344
rect 18969 25307 19027 25313
rect 20806 25304 20812 25316
rect 20864 25304 20870 25356
rect 21358 25344 21364 25356
rect 21319 25316 21364 25344
rect 21358 25304 21364 25316
rect 21416 25304 21422 25356
rect 22554 25276 22560 25288
rect 5684 25248 18373 25276
rect 22515 25248 22560 25276
rect 5684 25236 5690 25248
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 20070 25168 20076 25220
rect 20128 25208 20134 25220
rect 21545 25211 21603 25217
rect 21545 25208 21557 25211
rect 20128 25180 21557 25208
rect 20128 25168 20134 25180
rect 21545 25177 21557 25180
rect 21591 25177 21603 25211
rect 21545 25171 21603 25177
rect 9398 25100 9404 25152
rect 9456 25140 9462 25152
rect 20162 25140 20168 25152
rect 9456 25112 20168 25140
rect 9456 25100 9462 25112
rect 20162 25100 20168 25112
rect 20220 25140 20226 25152
rect 20349 25143 20407 25149
rect 20349 25140 20361 25143
rect 20220 25112 20361 25140
rect 20220 25100 20226 25112
rect 20349 25109 20361 25112
rect 20395 25109 20407 25143
rect 20349 25103 20407 25109
rect 20898 25100 20904 25152
rect 20956 25140 20962 25152
rect 23952 25140 23980 25443
rect 24486 25440 24492 25452
rect 24544 25440 24550 25492
rect 25038 25440 25044 25492
rect 25096 25480 25102 25492
rect 31386 25480 31392 25492
rect 25096 25452 31392 25480
rect 25096 25440 25102 25452
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 37369 25483 37427 25489
rect 37369 25449 37381 25483
rect 37415 25480 37427 25483
rect 37642 25480 37648 25492
rect 37415 25452 37648 25480
rect 37415 25449 37427 25452
rect 37369 25443 37427 25449
rect 37642 25440 37648 25452
rect 37700 25440 37706 25492
rect 24394 25372 24400 25424
rect 24452 25412 24458 25424
rect 24452 25384 25268 25412
rect 24452 25372 24458 25384
rect 24949 25347 25007 25353
rect 24949 25313 24961 25347
rect 24995 25313 25007 25347
rect 25130 25344 25136 25356
rect 25091 25316 25136 25344
rect 24949 25307 25007 25313
rect 24964 25276 24992 25307
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 25240 25353 25268 25384
rect 25424 25384 26556 25412
rect 25424 25353 25452 25384
rect 25225 25347 25283 25353
rect 25225 25313 25237 25347
rect 25271 25313 25283 25347
rect 25225 25307 25283 25313
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25313 25467 25347
rect 26050 25344 26056 25356
rect 26011 25316 26056 25344
rect 25409 25307 25467 25313
rect 26050 25304 26056 25316
rect 26108 25304 26114 25356
rect 26528 25353 26556 25384
rect 26329 25347 26387 25353
rect 26329 25344 26341 25347
rect 26160 25316 26341 25344
rect 24964 25248 25176 25276
rect 25148 25220 25176 25248
rect 25958 25236 25964 25288
rect 26016 25276 26022 25288
rect 26160 25276 26188 25316
rect 26329 25313 26341 25316
rect 26375 25313 26387 25347
rect 26329 25307 26387 25313
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25344 26571 25347
rect 26878 25344 26884 25356
rect 26559 25316 26884 25344
rect 26559 25313 26571 25316
rect 26513 25307 26571 25313
rect 26878 25304 26884 25316
rect 26936 25304 26942 25356
rect 36814 25304 36820 25356
rect 36872 25304 36878 25356
rect 37182 25344 37188 25356
rect 37143 25316 37188 25344
rect 37182 25304 37188 25316
rect 37240 25304 37246 25356
rect 26016 25248 26188 25276
rect 26237 25279 26295 25285
rect 26016 25236 26022 25248
rect 26237 25245 26249 25279
rect 26283 25276 26295 25279
rect 27706 25276 27712 25288
rect 26283 25248 27712 25276
rect 26283 25245 26295 25248
rect 26237 25239 26295 25245
rect 27706 25236 27712 25248
rect 27764 25236 27770 25288
rect 35250 25236 35256 25288
rect 35308 25276 35314 25288
rect 35434 25276 35440 25288
rect 35308 25248 35440 25276
rect 35308 25236 35314 25248
rect 35434 25236 35440 25248
rect 35492 25236 35498 25288
rect 24486 25168 24492 25220
rect 24544 25208 24550 25220
rect 25038 25208 25044 25220
rect 24544 25180 24900 25208
rect 24999 25180 25044 25208
rect 24544 25168 24550 25180
rect 20956 25112 23980 25140
rect 20956 25100 20962 25112
rect 24118 25100 24124 25152
rect 24176 25140 24182 25152
rect 24765 25143 24823 25149
rect 24765 25140 24777 25143
rect 24176 25112 24777 25140
rect 24176 25100 24182 25112
rect 24765 25109 24777 25112
rect 24811 25109 24823 25143
rect 24872 25140 24900 25180
rect 25038 25168 25044 25180
rect 25096 25168 25102 25220
rect 25130 25168 25136 25220
rect 25188 25168 25194 25220
rect 26145 25211 26203 25217
rect 26145 25177 26157 25211
rect 26191 25208 26203 25211
rect 34606 25208 34612 25220
rect 26191 25180 34612 25208
rect 26191 25177 26203 25180
rect 26145 25171 26203 25177
rect 34606 25168 34612 25180
rect 34664 25168 34670 25220
rect 25869 25143 25927 25149
rect 25869 25140 25881 25143
rect 24872 25112 25881 25140
rect 24765 25103 24823 25109
rect 25869 25109 25881 25112
rect 25915 25109 25927 25143
rect 25869 25103 25927 25109
rect 36722 25100 36728 25152
rect 36780 25140 36786 25152
rect 36832 25140 36860 25304
rect 36780 25112 36860 25140
rect 36780 25100 36786 25112
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 16574 24896 16580 24948
rect 16632 24936 16638 24948
rect 20898 24936 20904 24948
rect 16632 24908 20904 24936
rect 16632 24896 16638 24908
rect 20898 24896 20904 24908
rect 20956 24896 20962 24948
rect 23566 24936 23572 24948
rect 21008 24908 23572 24936
rect 1578 24828 1584 24880
rect 1636 24868 1642 24880
rect 4890 24868 4896 24880
rect 1636 24840 4896 24868
rect 1636 24828 1642 24840
rect 4890 24828 4896 24840
rect 4948 24828 4954 24880
rect 17144 24840 17356 24868
rect 15838 24760 15844 24812
rect 15896 24800 15902 24812
rect 17144 24800 17172 24840
rect 15896 24772 17172 24800
rect 15896 24760 15902 24772
rect 17218 24760 17224 24812
rect 17276 24760 17282 24812
rect 17328 24800 17356 24840
rect 21008 24800 21036 24908
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 23952 24908 24256 24936
rect 21266 24868 21272 24880
rect 17328 24772 18000 24800
rect 11790 24692 11796 24744
rect 11848 24732 11854 24744
rect 16853 24735 16911 24741
rect 16853 24732 16865 24735
rect 11848 24704 16865 24732
rect 11848 24692 11854 24704
rect 16853 24701 16865 24704
rect 16899 24701 16911 24735
rect 16853 24695 16911 24701
rect 17001 24735 17059 24741
rect 17001 24701 17013 24735
rect 17047 24732 17059 24735
rect 17236 24732 17264 24760
rect 17047 24704 17264 24732
rect 17047 24701 17059 24704
rect 17001 24695 17059 24701
rect 17310 24692 17316 24744
rect 17368 24741 17374 24744
rect 17972 24741 18000 24772
rect 18340 24772 21036 24800
rect 21100 24840 21272 24868
rect 17368 24732 17376 24741
rect 17957 24735 18015 24741
rect 17368 24704 17413 24732
rect 17368 24695 17376 24704
rect 17957 24701 17969 24735
rect 18003 24701 18015 24735
rect 17957 24695 18015 24701
rect 18050 24735 18108 24741
rect 18050 24701 18062 24735
rect 18096 24732 18108 24735
rect 18340 24732 18368 24772
rect 18096 24704 18368 24732
rect 18096 24701 18108 24704
rect 18050 24695 18108 24701
rect 17368 24692 17374 24695
rect 18414 24692 18420 24744
rect 18472 24741 18478 24744
rect 18472 24732 18480 24741
rect 18472 24704 18517 24732
rect 18472 24695 18480 24704
rect 18472 24692 18478 24695
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 21100 24741 21128 24840
rect 21266 24828 21272 24840
rect 21324 24828 21330 24880
rect 23952 24877 23980 24908
rect 23937 24871 23995 24877
rect 23937 24837 23949 24871
rect 23983 24837 23995 24871
rect 23937 24831 23995 24837
rect 22186 24760 22192 24812
rect 22244 24800 22250 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 22244 24772 23673 24800
rect 22244 24760 22250 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 24026 24760 24032 24812
rect 24084 24809 24090 24812
rect 24084 24800 24096 24809
rect 24228 24800 24256 24908
rect 25501 24871 25559 24877
rect 25501 24837 25513 24871
rect 25547 24868 25559 24871
rect 25547 24840 26004 24868
rect 25547 24837 25559 24840
rect 25501 24831 25559 24837
rect 25038 24800 25044 24812
rect 24084 24772 24129 24800
rect 24228 24772 25044 24800
rect 24084 24763 24096 24772
rect 24084 24760 24090 24763
rect 25038 24760 25044 24772
rect 25096 24760 25102 24812
rect 25976 24800 26004 24840
rect 28626 24828 28632 24880
rect 28684 24868 28690 24880
rect 32030 24868 32036 24880
rect 28684 24840 32036 24868
rect 28684 24828 28690 24840
rect 32030 24828 32036 24840
rect 32088 24828 32094 24880
rect 30006 24800 30012 24812
rect 25245 24772 25912 24800
rect 25976 24772 30012 24800
rect 20257 24735 20315 24741
rect 20257 24732 20269 24735
rect 19300 24704 20269 24732
rect 19300 24692 19306 24704
rect 20257 24701 20269 24704
rect 20303 24701 20315 24735
rect 20257 24695 20315 24701
rect 21085 24735 21143 24741
rect 21085 24701 21097 24735
rect 21131 24701 21143 24735
rect 21085 24695 21143 24701
rect 21177 24735 21235 24741
rect 21177 24701 21189 24735
rect 21223 24732 21235 24735
rect 21266 24732 21272 24744
rect 21223 24704 21272 24732
rect 21223 24701 21235 24704
rect 21177 24695 21235 24701
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 21361 24735 21419 24741
rect 21361 24701 21373 24735
rect 21407 24732 21419 24735
rect 21542 24732 21548 24744
rect 21407 24704 21548 24732
rect 21407 24701 21419 24704
rect 21361 24695 21419 24701
rect 21542 24692 21548 24704
rect 21600 24692 21606 24744
rect 22002 24692 22008 24744
rect 22060 24692 22066 24744
rect 22278 24692 22284 24744
rect 22336 24732 22342 24744
rect 22336 24704 22784 24732
rect 22336 24692 22342 24704
rect 17126 24664 17132 24676
rect 17087 24636 17132 24664
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17221 24667 17279 24673
rect 17221 24633 17233 24667
rect 17267 24664 17279 24667
rect 17267 24636 17632 24664
rect 17267 24633 17279 24636
rect 17221 24627 17279 24633
rect 5718 24556 5724 24608
rect 5776 24596 5782 24608
rect 17310 24596 17316 24608
rect 5776 24568 17316 24596
rect 5776 24556 5782 24568
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17402 24556 17408 24608
rect 17460 24596 17466 24608
rect 17497 24599 17555 24605
rect 17497 24596 17509 24599
rect 17460 24568 17509 24596
rect 17460 24556 17466 24568
rect 17497 24565 17509 24568
rect 17543 24565 17555 24599
rect 17604 24596 17632 24636
rect 17678 24624 17684 24676
rect 17736 24664 17742 24676
rect 18138 24664 18144 24676
rect 17736 24636 18144 24664
rect 17736 24624 17742 24636
rect 18138 24624 18144 24636
rect 18196 24664 18202 24676
rect 18233 24667 18291 24673
rect 18233 24664 18245 24667
rect 18196 24636 18245 24664
rect 18196 24624 18202 24636
rect 18233 24633 18245 24636
rect 18279 24633 18291 24667
rect 18233 24627 18291 24633
rect 18322 24624 18328 24676
rect 18380 24664 18386 24676
rect 18380 24636 18425 24664
rect 18380 24624 18386 24636
rect 18506 24624 18512 24676
rect 18564 24664 18570 24676
rect 20070 24664 20076 24676
rect 18564 24636 19933 24664
rect 20031 24636 20076 24664
rect 18564 24624 18570 24636
rect 18340 24596 18368 24624
rect 18598 24596 18604 24608
rect 17604 24568 18368 24596
rect 18559 24568 18604 24596
rect 17497 24559 17555 24565
rect 18598 24556 18604 24568
rect 18656 24556 18662 24608
rect 19905 24596 19933 24636
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 20180 24636 21772 24664
rect 20180 24596 20208 24636
rect 19905 24568 20208 24596
rect 21744 24596 21772 24636
rect 21818 24624 21824 24676
rect 21876 24664 21882 24676
rect 21913 24667 21971 24673
rect 21913 24664 21925 24667
rect 21876 24636 21925 24664
rect 21876 24624 21882 24636
rect 21913 24633 21925 24636
rect 21959 24664 21971 24667
rect 22020 24664 22048 24692
rect 22649 24667 22707 24673
rect 22649 24664 22661 24667
rect 21959 24636 22661 24664
rect 21959 24633 21971 24636
rect 21913 24627 21971 24633
rect 22649 24633 22661 24636
rect 22695 24633 22707 24667
rect 22756 24664 22784 24704
rect 23842 24692 23848 24744
rect 23900 24732 23906 24744
rect 24121 24735 24179 24741
rect 23900 24704 23945 24732
rect 23900 24692 23906 24704
rect 24121 24701 24133 24735
rect 24167 24701 24179 24735
rect 24121 24695 24179 24701
rect 24305 24735 24363 24741
rect 24305 24701 24317 24735
rect 24351 24732 24363 24735
rect 25245 24732 25273 24772
rect 25406 24732 25412 24744
rect 24351 24704 25273 24732
rect 25367 24704 25412 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 24136 24664 24164 24695
rect 25406 24692 25412 24704
rect 25464 24692 25470 24744
rect 25593 24735 25651 24741
rect 25593 24701 25605 24735
rect 25639 24701 25651 24735
rect 25593 24695 25651 24701
rect 25685 24735 25743 24741
rect 25685 24701 25697 24735
rect 25731 24732 25743 24735
rect 25774 24732 25780 24744
rect 25731 24704 25780 24732
rect 25731 24701 25743 24704
rect 25685 24695 25743 24701
rect 22756 24636 24164 24664
rect 22649 24627 22707 24633
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21744 24568 22017 24596
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22738 24596 22744 24608
rect 22699 24568 22744 24596
rect 22005 24559 22063 24565
rect 22738 24556 22744 24568
rect 22796 24556 22802 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 25225 24599 25283 24605
rect 25225 24596 25237 24599
rect 23440 24568 25237 24596
rect 23440 24556 23446 24568
rect 25225 24565 25237 24568
rect 25271 24565 25283 24599
rect 25608 24596 25636 24695
rect 25774 24692 25780 24704
rect 25832 24692 25838 24744
rect 25884 24741 25912 24772
rect 30006 24760 30012 24772
rect 30064 24760 30070 24812
rect 25869 24735 25927 24741
rect 25869 24701 25881 24735
rect 25915 24732 25927 24735
rect 26878 24732 26884 24744
rect 25915 24704 26884 24732
rect 25915 24701 25927 24704
rect 25869 24695 25927 24701
rect 26878 24692 26884 24704
rect 26936 24692 26942 24744
rect 37918 24732 37924 24744
rect 37879 24704 37924 24732
rect 37918 24692 37924 24704
rect 37976 24692 37982 24744
rect 31294 24596 31300 24608
rect 25608 24568 31300 24596
rect 25225 24559 25283 24565
rect 31294 24556 31300 24568
rect 31352 24556 31358 24608
rect 38105 24599 38163 24605
rect 38105 24565 38117 24599
rect 38151 24596 38163 24599
rect 38562 24596 38568 24608
rect 38151 24568 38568 24596
rect 38151 24565 38163 24568
rect 38105 24559 38163 24565
rect 38562 24556 38568 24568
rect 38620 24556 38626 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 18414 24392 18420 24404
rect 5592 24364 18420 24392
rect 5592 24352 5598 24364
rect 18414 24352 18420 24364
rect 18472 24352 18478 24404
rect 19242 24352 19248 24404
rect 19300 24392 19306 24404
rect 21545 24395 21603 24401
rect 21545 24392 21557 24395
rect 19300 24364 21557 24392
rect 19300 24352 19306 24364
rect 21545 24361 21557 24364
rect 21591 24361 21603 24395
rect 21545 24355 21603 24361
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 25774 24392 25780 24404
rect 23164 24364 25780 24392
rect 23164 24352 23170 24364
rect 25774 24352 25780 24364
rect 25832 24352 25838 24404
rect 29454 24352 29460 24404
rect 29512 24392 29518 24404
rect 37369 24395 37427 24401
rect 37369 24392 37381 24395
rect 29512 24364 37381 24392
rect 29512 24352 29518 24364
rect 37369 24361 37381 24364
rect 37415 24361 37427 24395
rect 37369 24355 37427 24361
rect 1854 24324 1860 24336
rect 1815 24296 1860 24324
rect 1854 24284 1860 24296
rect 1912 24284 1918 24336
rect 2041 24327 2099 24333
rect 2041 24293 2053 24327
rect 2087 24324 2099 24327
rect 2130 24324 2136 24336
rect 2087 24296 2136 24324
rect 2087 24293 2099 24296
rect 2041 24287 2099 24293
rect 2130 24284 2136 24296
rect 2188 24284 2194 24336
rect 16666 24284 16672 24336
rect 16724 24324 16730 24336
rect 17865 24327 17923 24333
rect 16724 24296 17632 24324
rect 16724 24284 16730 24296
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17604 24265 17632 24296
rect 17865 24293 17877 24327
rect 17911 24324 17923 24327
rect 18322 24324 18328 24336
rect 17911 24296 18328 24324
rect 17911 24293 17923 24296
rect 17865 24287 17923 24293
rect 18322 24284 18328 24296
rect 18380 24284 18386 24336
rect 18868 24327 18926 24333
rect 18868 24293 18880 24327
rect 18914 24324 18926 24327
rect 21634 24324 21640 24336
rect 18914 24296 21640 24324
rect 18914 24293 18926 24296
rect 18868 24287 18926 24293
rect 21634 24284 21640 24296
rect 21692 24284 21698 24336
rect 23198 24284 23204 24336
rect 23256 24324 23262 24336
rect 23256 24296 31754 24324
rect 23256 24284 23262 24296
rect 17590 24259 17648 24265
rect 17590 24225 17602 24259
rect 17636 24225 17648 24259
rect 17590 24219 17648 24225
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 17736 24228 17785 24256
rect 17736 24216 17742 24228
rect 17773 24225 17785 24228
rect 17819 24225 17831 24259
rect 17773 24219 17831 24225
rect 17962 24259 18020 24265
rect 17962 24225 17974 24259
rect 18008 24225 18020 24259
rect 17962 24219 18020 24225
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24256 18659 24259
rect 19978 24256 19984 24268
rect 18647 24228 19984 24256
rect 18647 24225 18659 24228
rect 18601 24219 18659 24225
rect 2958 24148 2964 24200
rect 3016 24188 3022 24200
rect 17972 24188 18000 24219
rect 19978 24216 19984 24228
rect 20036 24256 20042 24268
rect 20162 24256 20168 24268
rect 20036 24228 20168 24256
rect 20036 24216 20042 24228
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 21450 24256 21456 24268
rect 21411 24228 21456 24256
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 24670 24216 24676 24268
rect 24728 24256 24734 24268
rect 27246 24256 27252 24268
rect 24728 24228 27252 24256
rect 24728 24216 24734 24228
rect 27246 24216 27252 24228
rect 27304 24216 27310 24268
rect 3016 24160 6914 24188
rect 3016 24148 3022 24160
rect 1670 24080 1676 24132
rect 1728 24120 1734 24132
rect 6546 24120 6552 24132
rect 1728 24092 6552 24120
rect 1728 24080 1734 24092
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 6886 24052 6914 24160
rect 12406 24160 18000 24188
rect 12406 24052 12434 24160
rect 21358 24148 21364 24200
rect 21416 24188 21422 24200
rect 21542 24188 21548 24200
rect 21416 24160 21548 24188
rect 21416 24148 21422 24160
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 22002 24148 22008 24200
rect 22060 24188 22066 24200
rect 22738 24188 22744 24200
rect 22060 24160 22744 24188
rect 22060 24148 22066 24160
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 24026 24148 24032 24200
rect 24084 24188 24090 24200
rect 24302 24188 24308 24200
rect 24084 24160 24308 24188
rect 24084 24148 24090 24160
rect 24302 24148 24308 24160
rect 24360 24148 24366 24200
rect 31726 24188 31754 24296
rect 37182 24256 37188 24268
rect 37143 24228 37188 24256
rect 37182 24216 37188 24228
rect 37240 24216 37246 24268
rect 37550 24188 37556 24200
rect 31726 24160 37556 24188
rect 37550 24148 37556 24160
rect 37608 24148 37614 24200
rect 17126 24080 17132 24132
rect 17184 24120 17190 24132
rect 17678 24120 17684 24132
rect 17184 24092 17684 24120
rect 17184 24080 17190 24092
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 19536 24092 20116 24120
rect 18138 24052 18144 24064
rect 6886 24024 12434 24052
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 18414 24012 18420 24064
rect 18472 24052 18478 24064
rect 19536 24052 19564 24092
rect 18472 24024 19564 24052
rect 18472 24012 18478 24024
rect 19610 24012 19616 24064
rect 19668 24052 19674 24064
rect 19981 24055 20039 24061
rect 19981 24052 19993 24055
rect 19668 24024 19993 24052
rect 19668 24012 19674 24024
rect 19981 24021 19993 24024
rect 20027 24021 20039 24055
rect 20088 24052 20116 24092
rect 22554 24080 22560 24132
rect 22612 24120 22618 24132
rect 24489 24123 24547 24129
rect 24489 24120 24501 24123
rect 22612 24092 24501 24120
rect 22612 24080 22618 24092
rect 24489 24089 24501 24092
rect 24535 24089 24547 24123
rect 24489 24083 24547 24089
rect 27430 24080 27436 24132
rect 27488 24120 27494 24132
rect 36630 24120 36636 24132
rect 27488 24092 36636 24120
rect 27488 24080 27494 24092
rect 36630 24080 36636 24092
rect 36688 24080 36694 24132
rect 22002 24052 22008 24064
rect 20088 24024 22008 24052
rect 19981 24015 20039 24021
rect 22002 24012 22008 24024
rect 22060 24012 22066 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 31202 24052 31208 24064
rect 23624 24024 31208 24052
rect 23624 24012 23630 24024
rect 31202 24012 31208 24024
rect 31260 24012 31266 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 10502 23808 10508 23860
rect 10560 23848 10566 23860
rect 18046 23848 18052 23860
rect 10560 23820 18052 23848
rect 10560 23808 10566 23820
rect 18046 23808 18052 23820
rect 18104 23808 18110 23860
rect 18138 23808 18144 23860
rect 18196 23848 18202 23860
rect 27154 23848 27160 23860
rect 18196 23820 27160 23848
rect 18196 23808 18202 23820
rect 27154 23808 27160 23820
rect 27212 23808 27218 23860
rect 37277 23851 37335 23857
rect 37277 23817 37289 23851
rect 37323 23848 37335 23851
rect 37366 23848 37372 23860
rect 37323 23820 37372 23848
rect 37323 23817 37335 23820
rect 37277 23811 37335 23817
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 37921 23851 37979 23857
rect 37921 23817 37933 23851
rect 37967 23848 37979 23851
rect 38930 23848 38936 23860
rect 37967 23820 38936 23848
rect 37967 23817 37979 23820
rect 37921 23811 37979 23817
rect 38930 23808 38936 23820
rect 38988 23808 38994 23860
rect 2041 23783 2099 23789
rect 2041 23749 2053 23783
rect 2087 23780 2099 23783
rect 2222 23780 2228 23792
rect 2087 23752 2228 23780
rect 2087 23749 2099 23752
rect 2041 23743 2099 23749
rect 2222 23740 2228 23752
rect 2280 23740 2286 23792
rect 18693 23783 18751 23789
rect 18693 23749 18705 23783
rect 18739 23780 18751 23783
rect 19150 23780 19156 23792
rect 18739 23752 19156 23780
rect 18739 23749 18751 23752
rect 18693 23743 18751 23749
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 22094 23740 22100 23792
rect 22152 23780 22158 23792
rect 25406 23780 25412 23792
rect 22152 23752 25412 23780
rect 22152 23740 22158 23752
rect 25406 23740 25412 23752
rect 25464 23740 25470 23792
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 28534 23712 28540 23724
rect 18656 23684 28540 23712
rect 18656 23672 18662 23684
rect 28534 23672 28540 23684
rect 28592 23672 28598 23724
rect 1854 23644 1860 23656
rect 1815 23616 1860 23644
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 18506 23644 18512 23656
rect 18467 23616 18512 23644
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 19794 23644 19800 23656
rect 19208 23616 19800 23644
rect 19208 23604 19214 23616
rect 19794 23604 19800 23616
rect 19852 23604 19858 23656
rect 19978 23644 19984 23656
rect 19939 23616 19984 23644
rect 19978 23604 19984 23616
rect 20036 23604 20042 23656
rect 20714 23604 20720 23656
rect 20772 23644 20778 23656
rect 20898 23644 20904 23656
rect 20772 23616 20904 23644
rect 20772 23604 20778 23616
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23644 21419 23647
rect 21450 23644 21456 23656
rect 21407 23616 21456 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21450 23604 21456 23616
rect 21508 23604 21514 23656
rect 21545 23647 21603 23653
rect 21545 23613 21557 23647
rect 21591 23644 21603 23647
rect 21726 23644 21732 23656
rect 21591 23616 21732 23644
rect 21591 23613 21603 23616
rect 21545 23607 21603 23613
rect 21726 23604 21732 23616
rect 21784 23604 21790 23656
rect 22189 23647 22247 23653
rect 22189 23613 22201 23647
rect 22235 23644 22247 23647
rect 24670 23644 24676 23656
rect 22235 23616 24676 23644
rect 22235 23613 22247 23616
rect 22189 23607 22247 23613
rect 24670 23604 24676 23616
rect 24728 23604 24734 23656
rect 37458 23644 37464 23656
rect 37419 23616 37464 23644
rect 37458 23604 37464 23616
rect 37516 23604 37522 23656
rect 38102 23644 38108 23656
rect 38063 23616 38108 23644
rect 38102 23604 38108 23616
rect 38160 23604 38166 23656
rect 17402 23536 17408 23588
rect 17460 23576 17466 23588
rect 27522 23576 27528 23588
rect 17460 23548 27528 23576
rect 17460 23536 17466 23548
rect 27522 23536 27528 23548
rect 27580 23536 27586 23588
rect 20073 23511 20131 23517
rect 20073 23477 20085 23511
rect 20119 23508 20131 23511
rect 20898 23508 20904 23520
rect 20119 23480 20904 23508
rect 20119 23477 20131 23480
rect 20073 23471 20131 23477
rect 20898 23468 20904 23480
rect 20956 23468 20962 23520
rect 21450 23468 21456 23520
rect 21508 23508 21514 23520
rect 22005 23511 22063 23517
rect 22005 23508 22017 23511
rect 21508 23480 22017 23508
rect 21508 23468 21514 23480
rect 22005 23477 22017 23480
rect 22051 23477 22063 23511
rect 22005 23471 22063 23477
rect 23842 23468 23848 23520
rect 23900 23508 23906 23520
rect 24302 23508 24308 23520
rect 23900 23480 24308 23508
rect 23900 23468 23906 23480
rect 24302 23468 24308 23480
rect 24360 23468 24366 23520
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 31938 23508 31944 23520
rect 25096 23480 31944 23508
rect 25096 23468 25102 23480
rect 31938 23468 31944 23480
rect 31996 23468 32002 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 13538 23264 13544 23316
rect 13596 23304 13602 23316
rect 16114 23304 16120 23316
rect 13596 23276 16120 23304
rect 13596 23264 13602 23276
rect 16114 23264 16120 23276
rect 16172 23264 16178 23316
rect 17678 23304 17684 23316
rect 17639 23276 17684 23304
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 18322 23304 18328 23316
rect 18283 23276 18328 23304
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 19978 23264 19984 23316
rect 20036 23304 20042 23316
rect 20165 23307 20223 23313
rect 20165 23304 20177 23307
rect 20036 23276 20177 23304
rect 20036 23264 20042 23276
rect 20165 23273 20177 23276
rect 20211 23304 20223 23307
rect 20622 23304 20628 23316
rect 20211 23276 20628 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 20806 23264 20812 23316
rect 20864 23304 20870 23316
rect 22002 23304 22008 23316
rect 20864 23276 22008 23304
rect 20864 23264 20870 23276
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23900 23276 23949 23304
rect 23900 23264 23906 23276
rect 23937 23273 23949 23276
rect 23983 23304 23995 23307
rect 24394 23304 24400 23316
rect 23983 23276 24400 23304
rect 23983 23273 23995 23276
rect 23937 23267 23995 23273
rect 24394 23264 24400 23276
rect 24452 23264 24458 23316
rect 27890 23264 27896 23316
rect 27948 23304 27954 23316
rect 28902 23304 28908 23316
rect 27948 23276 28908 23304
rect 27948 23264 27954 23276
rect 28902 23264 28908 23276
rect 28960 23264 28966 23316
rect 34146 23264 34152 23316
rect 34204 23304 34210 23316
rect 37369 23307 37427 23313
rect 37369 23304 37381 23307
rect 34204 23276 37381 23304
rect 34204 23264 34210 23276
rect 37369 23273 37381 23276
rect 37415 23273 37427 23307
rect 37369 23267 37427 23273
rect 15930 23196 15936 23248
rect 15988 23236 15994 23248
rect 16574 23236 16580 23248
rect 15988 23208 16580 23236
rect 15988 23196 15994 23208
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 19052 23239 19110 23245
rect 17512 23208 18633 23236
rect 17512 23180 17540 23208
rect 17494 23168 17500 23180
rect 17407 23140 17500 23168
rect 17494 23128 17500 23140
rect 17552 23128 17558 23180
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 18230 23168 18236 23180
rect 18187 23140 18236 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 18230 23128 18236 23140
rect 18288 23168 18294 23180
rect 18506 23168 18512 23180
rect 18288 23140 18512 23168
rect 18288 23128 18294 23140
rect 18506 23128 18512 23140
rect 18564 23128 18570 23180
rect 18605 23168 18633 23208
rect 19052 23205 19064 23239
rect 19098 23236 19110 23239
rect 22824 23239 22882 23245
rect 19098 23208 22784 23236
rect 19098 23205 19110 23208
rect 19052 23199 19110 23205
rect 20070 23168 20076 23180
rect 18605 23140 20076 23168
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 21177 23171 21235 23177
rect 21177 23168 21189 23171
rect 20864 23140 21189 23168
rect 20864 23128 20870 23140
rect 21177 23137 21189 23140
rect 21223 23168 21235 23171
rect 21818 23168 21824 23180
rect 21223 23140 21824 23168
rect 21223 23137 21235 23140
rect 21177 23131 21235 23137
rect 21818 23128 21824 23140
rect 21876 23128 21882 23180
rect 22756 23168 22784 23208
rect 22824 23205 22836 23239
rect 22870 23236 22882 23239
rect 24118 23236 24124 23248
rect 22870 23208 24124 23236
rect 22870 23205 22882 23208
rect 22824 23199 22882 23205
rect 24118 23196 24124 23208
rect 24176 23196 24182 23248
rect 25498 23196 25504 23248
rect 25556 23236 25562 23248
rect 28534 23236 28540 23248
rect 25556 23208 28540 23236
rect 25556 23196 25562 23208
rect 28534 23196 28540 23208
rect 28592 23196 28598 23248
rect 27062 23168 27068 23180
rect 22756 23140 27068 23168
rect 27062 23128 27068 23140
rect 27120 23128 27126 23180
rect 37182 23168 37188 23180
rect 37143 23140 37188 23168
rect 37182 23128 37188 23140
rect 37240 23128 37246 23180
rect 9950 23060 9956 23112
rect 10008 23100 10014 23112
rect 13170 23100 13176 23112
rect 10008 23072 13176 23100
rect 10008 23060 10014 23072
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23069 18843 23103
rect 18785 23063 18843 23069
rect 18138 22992 18144 23044
rect 18196 23032 18202 23044
rect 18506 23032 18512 23044
rect 18196 23004 18512 23032
rect 18196 22992 18202 23004
rect 18506 22992 18512 23004
rect 18564 22992 18570 23044
rect 18800 22964 18828 23063
rect 20162 23060 20168 23112
rect 20220 23100 20226 23112
rect 21450 23100 21456 23112
rect 20220 23072 21456 23100
rect 20220 23060 20226 23072
rect 21450 23060 21456 23072
rect 21508 23060 21514 23112
rect 22554 23100 22560 23112
rect 22515 23072 22560 23100
rect 22554 23060 22560 23072
rect 22612 23060 22618 23112
rect 20180 22964 20208 23060
rect 18800 22936 20208 22964
rect 20622 22924 20628 22976
rect 20680 22964 20686 22976
rect 21269 22967 21327 22973
rect 21269 22964 21281 22967
rect 20680 22936 21281 22964
rect 20680 22924 20686 22936
rect 21269 22933 21281 22936
rect 21315 22933 21327 22967
rect 21269 22927 21327 22933
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 24578 22964 24584 22976
rect 22152 22936 24584 22964
rect 22152 22924 22158 22936
rect 24578 22924 24584 22936
rect 24636 22924 24642 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 18874 22760 18880 22772
rect 18253 22732 18880 22760
rect 18046 22652 18052 22704
rect 18104 22692 18110 22704
rect 18253 22692 18281 22732
rect 18874 22720 18880 22732
rect 18932 22720 18938 22772
rect 22370 22720 22376 22772
rect 22428 22760 22434 22772
rect 22741 22763 22799 22769
rect 22741 22760 22753 22763
rect 22428 22732 22753 22760
rect 22428 22720 22434 22732
rect 22741 22729 22753 22732
rect 22787 22760 22799 22763
rect 23106 22760 23112 22772
rect 22787 22732 23112 22760
rect 22787 22729 22799 22732
rect 22741 22723 22799 22729
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 23934 22760 23940 22772
rect 23768 22732 23940 22760
rect 18598 22692 18604 22704
rect 18104 22664 18281 22692
rect 18559 22664 18604 22692
rect 18104 22652 18110 22664
rect 1394 22556 1400 22568
rect 1355 22528 1400 22556
rect 1394 22516 1400 22528
rect 1452 22516 1458 22568
rect 13262 22516 13268 22568
rect 13320 22556 13326 22568
rect 18138 22565 18144 22568
rect 17957 22559 18015 22565
rect 17957 22556 17969 22559
rect 13320 22528 17969 22556
rect 13320 22516 13326 22528
rect 17957 22525 17969 22528
rect 18003 22525 18015 22559
rect 17957 22519 18015 22525
rect 18105 22559 18144 22565
rect 18105 22525 18117 22559
rect 18105 22519 18144 22525
rect 18138 22516 18144 22519
rect 18196 22516 18202 22568
rect 18253 22565 18281 22664
rect 18598 22652 18604 22664
rect 18656 22652 18662 22704
rect 19150 22624 19156 22636
rect 18340 22596 19156 22624
rect 18340 22565 18368 22596
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 23768 22624 23796 22732
rect 23934 22720 23940 22732
rect 23992 22720 23998 22772
rect 37461 22763 37519 22769
rect 37461 22729 37473 22763
rect 37507 22760 37519 22763
rect 37734 22760 37740 22772
rect 37507 22732 37740 22760
rect 37507 22729 37519 22732
rect 37461 22723 37519 22729
rect 37734 22720 37740 22732
rect 37792 22720 37798 22772
rect 38010 22720 38016 22772
rect 38068 22760 38074 22772
rect 38105 22763 38163 22769
rect 38105 22760 38117 22763
rect 38068 22732 38117 22760
rect 38068 22720 38074 22732
rect 38105 22729 38117 22732
rect 38151 22729 38163 22763
rect 38105 22723 38163 22729
rect 23845 22695 23903 22701
rect 23845 22661 23857 22695
rect 23891 22692 23903 22695
rect 34514 22692 34520 22704
rect 23891 22664 34520 22692
rect 23891 22661 23903 22664
rect 23845 22655 23903 22661
rect 34514 22652 34520 22664
rect 34572 22652 34578 22704
rect 23946 22627 24004 22633
rect 23946 22624 23958 22627
rect 23768 22596 23958 22624
rect 23946 22593 23958 22596
rect 23992 22593 24004 22627
rect 23946 22587 24004 22593
rect 18233 22559 18291 22565
rect 18233 22525 18245 22559
rect 18279 22525 18291 22559
rect 18233 22519 18291 22525
rect 18325 22559 18383 22565
rect 18325 22525 18337 22559
rect 18371 22525 18383 22559
rect 18325 22519 18383 22525
rect 18422 22559 18480 22565
rect 18422 22525 18434 22559
rect 18468 22525 18480 22559
rect 18422 22519 18480 22525
rect 21361 22559 21419 22565
rect 21361 22525 21373 22559
rect 21407 22556 21419 22559
rect 21450 22556 21456 22568
rect 21407 22528 21456 22556
rect 21407 22525 21419 22528
rect 21361 22519 21419 22525
rect 1762 22448 1768 22500
rect 1820 22488 1826 22500
rect 5810 22488 5816 22500
rect 1820 22460 5816 22488
rect 1820 22448 1826 22460
rect 5810 22448 5816 22460
rect 5868 22448 5874 22500
rect 7558 22448 7564 22500
rect 7616 22488 7622 22500
rect 18432 22488 18460 22519
rect 21450 22516 21456 22528
rect 21508 22516 21514 22568
rect 21628 22559 21686 22565
rect 21628 22525 21640 22559
rect 21674 22556 21686 22559
rect 23382 22556 23388 22568
rect 21674 22528 23388 22556
rect 21674 22525 21686 22528
rect 21628 22519 21686 22525
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 23753 22559 23811 22565
rect 23753 22525 23765 22559
rect 23799 22556 23811 22559
rect 24046 22559 24104 22565
rect 23799 22528 23884 22556
rect 23799 22525 23811 22528
rect 23753 22519 23811 22525
rect 7616 22460 18460 22488
rect 7616 22448 7622 22460
rect 23566 22420 23572 22432
rect 23527 22392 23572 22420
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 23856 22420 23884 22528
rect 24046 22525 24058 22559
rect 24092 22525 24104 22559
rect 24210 22556 24216 22568
rect 24171 22528 24216 22556
rect 24046 22519 24104 22525
rect 24053 22488 24081 22519
rect 24210 22516 24216 22528
rect 24268 22556 24274 22568
rect 24394 22556 24400 22568
rect 24268 22528 24400 22556
rect 24268 22516 24274 22528
rect 24394 22516 24400 22528
rect 24452 22516 24458 22568
rect 37274 22556 37280 22568
rect 37235 22528 37280 22556
rect 37274 22516 37280 22528
rect 37332 22516 37338 22568
rect 37918 22556 37924 22568
rect 37879 22528 37924 22556
rect 37918 22516 37924 22528
rect 37976 22516 37982 22568
rect 24053 22460 24256 22488
rect 24228 22432 24256 22460
rect 34054 22448 34060 22500
rect 34112 22488 34118 22500
rect 34606 22488 34612 22500
rect 34112 22460 34612 22488
rect 34112 22448 34118 22460
rect 34606 22448 34612 22460
rect 34664 22448 34670 22500
rect 24026 22420 24032 22432
rect 23856 22392 24032 22420
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 24210 22380 24216 22432
rect 24268 22380 24274 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 14700 22188 17908 22216
rect 14700 22176 14706 22188
rect 17880 22148 17908 22188
rect 18598 22176 18604 22228
rect 18656 22216 18662 22228
rect 23198 22216 23204 22228
rect 18656 22188 23204 22216
rect 18656 22176 18662 22188
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 23842 22176 23848 22228
rect 23900 22216 23906 22228
rect 24486 22216 24492 22228
rect 23900 22188 24492 22216
rect 23900 22176 23906 22188
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 18874 22148 18880 22160
rect 17880 22120 18644 22148
rect 18835 22120 18880 22148
rect 1394 22080 1400 22092
rect 1355 22052 1400 22080
rect 1394 22040 1400 22052
rect 1452 22040 1458 22092
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 18616 22089 18644 22120
rect 18874 22108 18880 22120
rect 18932 22108 18938 22160
rect 18969 22151 19027 22157
rect 18969 22117 18981 22151
rect 19015 22148 19027 22151
rect 19150 22148 19156 22160
rect 19015 22120 19156 22148
rect 19015 22117 19027 22120
rect 18969 22111 19027 22117
rect 19150 22108 19156 22120
rect 19208 22108 19214 22160
rect 20714 22148 20720 22160
rect 19260 22120 20720 22148
rect 18590 22083 18648 22089
rect 17828 22052 17873 22080
rect 17828 22040 17834 22052
rect 18590 22049 18602 22083
rect 18636 22049 18648 22083
rect 18590 22043 18648 22049
rect 18721 22083 18779 22089
rect 18721 22049 18733 22083
rect 18767 22049 18779 22083
rect 19066 22083 19124 22089
rect 19066 22080 19078 22083
rect 18721 22043 18779 22049
rect 18892 22052 19078 22080
rect 3602 21972 3608 22024
rect 3660 22012 3666 22024
rect 17126 22012 17132 22024
rect 3660 21984 17132 22012
rect 3660 21972 3666 21984
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 17402 22012 17408 22024
rect 17363 21984 17408 22012
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 17954 22012 17960 22024
rect 17915 21984 17960 22012
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 1581 21947 1639 21953
rect 1581 21913 1593 21947
rect 1627 21944 1639 21947
rect 1670 21944 1676 21956
rect 1627 21916 1676 21944
rect 1627 21913 1639 21916
rect 1581 21907 1639 21913
rect 1670 21904 1676 21916
rect 1728 21904 1734 21956
rect 17954 21836 17960 21888
rect 18012 21876 18018 21888
rect 18230 21876 18236 21888
rect 18012 21848 18236 21876
rect 18012 21836 18018 21848
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18736 21876 18764 22043
rect 18892 22024 18920 22052
rect 19066 22049 19078 22052
rect 19112 22049 19124 22083
rect 19066 22043 19124 22049
rect 18874 21972 18880 22024
rect 18932 21972 18938 22024
rect 19260 21953 19288 22120
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 24394 22108 24400 22160
rect 24452 22148 24458 22160
rect 24452 22120 25176 22148
rect 24452 22108 24458 22120
rect 20162 22080 20168 22092
rect 20123 22052 20168 22080
rect 20162 22040 20168 22052
rect 20220 22040 20226 22092
rect 20432 22083 20490 22089
rect 20432 22049 20444 22083
rect 20478 22080 20490 22083
rect 21358 22080 21364 22092
rect 20478 22052 21364 22080
rect 20478 22049 20490 22052
rect 20432 22043 20490 22049
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 22554 22080 22560 22092
rect 22515 22052 22560 22080
rect 22554 22040 22560 22052
rect 22612 22040 22618 22092
rect 22824 22083 22882 22089
rect 22824 22049 22836 22083
rect 22870 22080 22882 22083
rect 24670 22080 24676 22092
rect 22870 22052 24072 22080
rect 24631 22052 24676 22080
rect 22870 22049 22882 22052
rect 22824 22043 22882 22049
rect 24044 22012 24072 22052
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 25148 22089 25176 22120
rect 24857 22083 24915 22089
rect 24857 22049 24869 22083
rect 24903 22080 24915 22083
rect 25133 22083 25191 22089
rect 24903 22052 25084 22080
rect 24903 22049 24915 22052
rect 24857 22043 24915 22049
rect 24946 22012 24952 22024
rect 24044 21984 24624 22012
rect 24907 21984 24952 22012
rect 19245 21947 19303 21953
rect 19245 21913 19257 21947
rect 19291 21913 19303 21947
rect 19245 21907 19303 21913
rect 21450 21876 21456 21888
rect 18736 21848 21456 21876
rect 21450 21836 21456 21848
rect 21508 21836 21514 21888
rect 21545 21879 21603 21885
rect 21545 21845 21557 21879
rect 21591 21876 21603 21879
rect 21726 21876 21732 21888
rect 21591 21848 21732 21876
rect 21591 21845 21603 21848
rect 21545 21839 21603 21845
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 23198 21836 23204 21888
rect 23256 21876 23262 21888
rect 23474 21876 23480 21888
rect 23256 21848 23480 21876
rect 23256 21836 23262 21848
rect 23474 21836 23480 21848
rect 23532 21876 23538 21888
rect 23937 21879 23995 21885
rect 23937 21876 23949 21879
rect 23532 21848 23949 21876
rect 23532 21836 23538 21848
rect 23937 21845 23949 21848
rect 23983 21845 23995 21879
rect 24486 21876 24492 21888
rect 24447 21848 24492 21876
rect 23937 21839 23995 21845
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 24596 21876 24624 21984
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 25056 22012 25084 22052
rect 25133 22049 25145 22083
rect 25179 22049 25191 22083
rect 37182 22080 37188 22092
rect 37143 22052 37188 22080
rect 25133 22043 25191 22049
rect 37182 22040 37188 22052
rect 37240 22040 37246 22092
rect 30466 22012 30472 22024
rect 25056 21984 30472 22012
rect 30466 21972 30472 21984
rect 30524 21972 30530 22024
rect 24765 21947 24823 21953
rect 24765 21913 24777 21947
rect 24811 21944 24823 21947
rect 35250 21944 35256 21956
rect 24811 21916 35256 21944
rect 24811 21913 24823 21916
rect 24765 21907 24823 21913
rect 35250 21904 35256 21916
rect 35308 21904 35314 21956
rect 25222 21876 25228 21888
rect 24596 21848 25228 21876
rect 25222 21836 25228 21848
rect 25280 21836 25286 21888
rect 28534 21836 28540 21888
rect 28592 21876 28598 21888
rect 37369 21879 37427 21885
rect 37369 21876 37381 21879
rect 28592 21848 37381 21876
rect 28592 21836 28598 21848
rect 37369 21845 37381 21848
rect 37415 21845 37427 21879
rect 37369 21839 37427 21845
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 16850 21632 16856 21684
rect 16908 21672 16914 21684
rect 16908 21644 17356 21672
rect 16908 21632 16914 21644
rect 10594 21564 10600 21616
rect 10652 21604 10658 21616
rect 10652 21576 17264 21604
rect 10652 21564 10658 21576
rect 1670 21428 1676 21480
rect 1728 21468 1734 21480
rect 5626 21468 5632 21480
rect 1728 21440 5632 21468
rect 1728 21428 1734 21440
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 14826 21428 14832 21480
rect 14884 21468 14890 21480
rect 16942 21477 16948 21480
rect 16761 21471 16819 21477
rect 16761 21468 16773 21471
rect 14884 21440 16773 21468
rect 14884 21428 14890 21440
rect 16761 21437 16773 21440
rect 16807 21437 16819 21471
rect 16761 21431 16819 21437
rect 16909 21471 16948 21477
rect 16909 21437 16921 21471
rect 16909 21431 16948 21437
rect 16942 21428 16948 21431
rect 17000 21428 17006 21480
rect 17126 21468 17132 21480
rect 17087 21440 17132 21468
rect 17126 21428 17132 21440
rect 17184 21428 17190 21480
rect 17236 21477 17264 21576
rect 17226 21471 17284 21477
rect 17226 21437 17238 21471
rect 17272 21437 17284 21471
rect 17328 21468 17356 21644
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 18506 21672 18512 21684
rect 17460 21644 18373 21672
rect 18467 21644 18512 21672
rect 17460 21632 17466 21644
rect 18046 21564 18052 21616
rect 18104 21564 18110 21616
rect 18345 21604 18373 21644
rect 18506 21632 18512 21644
rect 18564 21632 18570 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 20257 21675 20315 21681
rect 20257 21672 20269 21675
rect 18656 21644 20269 21672
rect 18656 21632 18662 21644
rect 20257 21641 20269 21644
rect 20303 21641 20315 21675
rect 21726 21672 21732 21684
rect 20257 21635 20315 21641
rect 20824 21644 21732 21672
rect 18874 21604 18880 21616
rect 18345 21576 18880 21604
rect 18874 21564 18880 21576
rect 18932 21604 18938 21616
rect 20824 21604 20852 21644
rect 21726 21632 21732 21644
rect 21784 21632 21790 21684
rect 22189 21675 22247 21681
rect 22189 21641 22201 21675
rect 22235 21672 22247 21675
rect 22278 21672 22284 21684
rect 22235 21644 22284 21672
rect 22235 21641 22247 21644
rect 22189 21635 22247 21641
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 35986 21632 35992 21684
rect 36044 21672 36050 21684
rect 37461 21675 37519 21681
rect 37461 21672 37473 21675
rect 36044 21644 37473 21672
rect 36044 21632 36050 21644
rect 37461 21641 37473 21644
rect 37507 21641 37519 21675
rect 37461 21635 37519 21641
rect 18932 21576 20852 21604
rect 18932 21564 18938 21576
rect 37090 21564 37096 21616
rect 37148 21604 37154 21616
rect 38105 21607 38163 21613
rect 38105 21604 38117 21607
rect 37148 21576 38117 21604
rect 37148 21564 37154 21576
rect 38105 21573 38117 21576
rect 38151 21573 38163 21607
rect 38105 21567 38163 21573
rect 18064 21536 18092 21564
rect 18064 21508 18184 21536
rect 18156 21477 18184 21508
rect 20162 21496 20168 21548
rect 20220 21536 20226 21548
rect 20622 21536 20628 21548
rect 20220 21508 20628 21536
rect 20220 21496 20226 21508
rect 20622 21496 20628 21508
rect 20680 21536 20686 21548
rect 20809 21539 20867 21545
rect 20809 21536 20821 21539
rect 20680 21508 20821 21536
rect 20680 21496 20686 21508
rect 20809 21505 20821 21508
rect 20855 21505 20867 21539
rect 20809 21499 20867 21505
rect 22554 21496 22560 21548
rect 22612 21536 22618 21548
rect 22741 21539 22799 21545
rect 22741 21536 22753 21539
rect 22612 21508 22753 21536
rect 22612 21496 22618 21508
rect 22741 21505 22753 21508
rect 22787 21505 22799 21539
rect 22741 21499 22799 21505
rect 17854 21471 17912 21477
rect 17854 21468 17866 21471
rect 17328 21440 17866 21468
rect 17226 21431 17284 21437
rect 17854 21437 17866 21440
rect 17900 21437 17912 21471
rect 17854 21431 17912 21437
rect 18013 21471 18071 21477
rect 18013 21437 18025 21471
rect 18059 21437 18071 21471
rect 18013 21431 18071 21437
rect 18141 21471 18199 21477
rect 18141 21437 18153 21471
rect 18187 21437 18199 21471
rect 18141 21431 18199 21437
rect 1578 21360 1584 21412
rect 1636 21400 1642 21412
rect 14458 21400 14464 21412
rect 1636 21372 14464 21400
rect 1636 21360 1642 21372
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 17034 21400 17040 21412
rect 16995 21372 17040 21400
rect 17034 21360 17040 21372
rect 17092 21360 17098 21412
rect 17402 21332 17408 21344
rect 17363 21304 17408 21332
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 18028 21332 18056 21431
rect 18322 21428 18328 21480
rect 18380 21477 18386 21480
rect 18380 21468 18388 21477
rect 18380 21440 18425 21468
rect 18380 21431 18388 21440
rect 18380 21428 18386 21431
rect 18782 21428 18788 21480
rect 18840 21468 18846 21480
rect 21076 21471 21134 21477
rect 18840 21440 20116 21468
rect 18840 21428 18846 21440
rect 18233 21403 18291 21409
rect 18233 21369 18245 21403
rect 18279 21400 18291 21403
rect 18506 21400 18512 21412
rect 18279 21372 18512 21400
rect 18279 21369 18291 21372
rect 18233 21363 18291 21369
rect 18506 21360 18512 21372
rect 18564 21400 18570 21412
rect 19150 21400 19156 21412
rect 18564 21372 19156 21400
rect 18564 21360 18570 21372
rect 19150 21360 19156 21372
rect 19208 21360 19214 21412
rect 19978 21332 19984 21344
rect 18028 21304 19984 21332
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20088 21332 20116 21440
rect 21076 21437 21088 21471
rect 21122 21468 21134 21471
rect 22186 21468 22192 21480
rect 21122 21440 22192 21468
rect 21122 21437 21134 21440
rect 21076 21431 21134 21437
rect 22186 21428 22192 21440
rect 22244 21428 22250 21480
rect 23008 21471 23066 21477
rect 23008 21437 23020 21471
rect 23054 21468 23066 21471
rect 23842 21468 23848 21480
rect 23054 21440 23848 21468
rect 23054 21437 23066 21440
rect 23008 21431 23066 21437
rect 23842 21428 23848 21440
rect 23900 21428 23906 21480
rect 37274 21468 37280 21480
rect 37235 21440 37280 21468
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 37918 21468 37924 21480
rect 37879 21440 37924 21468
rect 37918 21428 37924 21440
rect 37976 21428 37982 21480
rect 20165 21403 20223 21409
rect 20165 21369 20177 21403
rect 20211 21400 20223 21403
rect 21542 21400 21548 21412
rect 20211 21372 21548 21400
rect 20211 21369 20223 21372
rect 20165 21363 20223 21369
rect 21542 21360 21548 21372
rect 21600 21360 21606 21412
rect 25958 21400 25964 21412
rect 24136 21372 25964 21400
rect 24136 21341 24164 21372
rect 25958 21360 25964 21372
rect 26016 21360 26022 21412
rect 32674 21360 32680 21412
rect 32732 21400 32738 21412
rect 33410 21400 33416 21412
rect 32732 21372 33416 21400
rect 32732 21360 32738 21372
rect 33410 21360 33416 21372
rect 33468 21360 33474 21412
rect 24121 21335 24179 21341
rect 24121 21332 24133 21335
rect 20088 21304 24133 21332
rect 24121 21301 24133 21304
rect 24167 21301 24179 21335
rect 24121 21295 24179 21301
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 2682 21128 2688 21140
rect 1627 21100 2688 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 2682 21088 2688 21100
rect 2740 21088 2746 21140
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 22094 21128 22100 21140
rect 17460 21100 22100 21128
rect 17460 21088 17466 21100
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 28166 21128 28172 21140
rect 22612 21100 28172 21128
rect 22612 21088 22618 21100
rect 28166 21088 28172 21100
rect 28224 21088 28230 21140
rect 17034 21020 17040 21072
rect 17092 21060 17098 21072
rect 18046 21060 18052 21072
rect 17092 21032 18052 21060
rect 17092 21020 17098 21032
rect 18046 21020 18052 21032
rect 18104 21020 18110 21072
rect 18141 21063 18199 21069
rect 18141 21029 18153 21063
rect 18187 21060 18199 21063
rect 18506 21060 18512 21072
rect 18187 21032 18512 21060
rect 18187 21029 18199 21032
rect 18141 21023 18199 21029
rect 18506 21020 18512 21032
rect 18564 21020 18570 21072
rect 20806 21060 20812 21072
rect 20767 21032 20812 21060
rect 20806 21020 20812 21032
rect 20864 21020 20870 21072
rect 23750 21020 23756 21072
rect 23808 21020 23814 21072
rect 24118 21060 24124 21072
rect 23952 21032 24124 21060
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 17773 20995 17831 21001
rect 17773 20992 17785 20995
rect 15344 20964 17785 20992
rect 15344 20952 15350 20964
rect 17773 20961 17785 20964
rect 17819 20961 17831 20995
rect 17773 20955 17831 20961
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 17920 20964 17965 20992
rect 17920 20952 17926 20964
rect 18230 20952 18236 21004
rect 18288 21001 18294 21004
rect 18288 20992 18296 21001
rect 22554 20992 22560 21004
rect 18288 20964 18333 20992
rect 18432 20964 22560 20992
rect 18288 20955 18296 20964
rect 18288 20952 18294 20955
rect 6454 20884 6460 20936
rect 6512 20924 6518 20936
rect 18322 20924 18328 20936
rect 6512 20896 18328 20924
rect 6512 20884 6518 20896
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 18432 20865 18460 20964
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23474 20992 23480 21004
rect 23435 20964 23480 20992
rect 23474 20952 23480 20964
rect 23532 20952 23538 21004
rect 23661 20995 23719 21001
rect 23661 20961 23673 20995
rect 23707 20992 23719 20995
rect 23768 20992 23796 21020
rect 23952 21001 23980 21032
rect 24118 21020 24124 21032
rect 24176 21060 24182 21072
rect 24394 21060 24400 21072
rect 24176 21032 24400 21060
rect 24176 21020 24182 21032
rect 24394 21020 24400 21032
rect 24452 21060 24458 21072
rect 24452 21032 25084 21060
rect 24452 21020 24458 21032
rect 23707 20964 23796 20992
rect 23937 20995 23995 21001
rect 23707 20961 23719 20964
rect 23661 20955 23719 20961
rect 23937 20961 23949 20995
rect 23983 20961 23995 20995
rect 24578 20992 24584 21004
rect 24539 20964 24584 20992
rect 23937 20955 23995 20961
rect 24578 20952 24584 20964
rect 24636 20952 24642 21004
rect 24762 20992 24768 21004
rect 24723 20964 24768 20992
rect 24762 20952 24768 20964
rect 24820 20952 24826 21004
rect 25056 21001 25084 21032
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 21876 20896 23765 20924
rect 21876 20884 21882 20896
rect 23753 20893 23765 20896
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 23842 20884 23848 20936
rect 23900 20924 23906 20936
rect 24857 20927 24915 20933
rect 24857 20924 24869 20927
rect 23900 20896 24869 20924
rect 23900 20884 23906 20896
rect 24857 20893 24869 20896
rect 24903 20893 24915 20927
rect 36446 20924 36452 20936
rect 24857 20887 24915 20893
rect 25424 20896 36452 20924
rect 18417 20859 18475 20865
rect 18417 20825 18429 20859
rect 18463 20825 18475 20859
rect 18417 20819 18475 20825
rect 19978 20816 19984 20868
rect 20036 20856 20042 20868
rect 20622 20856 20628 20868
rect 20036 20828 20628 20856
rect 20036 20816 20042 20828
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 23569 20859 23627 20865
rect 23569 20825 23581 20859
rect 23615 20856 23627 20859
rect 24673 20859 24731 20865
rect 23615 20828 24624 20856
rect 23615 20825 23627 20828
rect 23569 20819 23627 20825
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 20901 20791 20959 20797
rect 20901 20788 20913 20791
rect 17184 20760 20913 20788
rect 17184 20748 17190 20760
rect 20901 20757 20913 20760
rect 20947 20757 20959 20791
rect 20901 20751 20959 20757
rect 21358 20748 21364 20800
rect 21416 20788 21422 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 21416 20760 23305 20788
rect 21416 20748 21422 20760
rect 23293 20757 23305 20760
rect 23339 20757 23351 20791
rect 24394 20788 24400 20800
rect 24355 20760 24400 20788
rect 23293 20751 23351 20757
rect 24394 20748 24400 20760
rect 24452 20748 24458 20800
rect 24596 20788 24624 20828
rect 24673 20825 24685 20859
rect 24719 20856 24731 20859
rect 25424 20856 25452 20896
rect 36446 20884 36452 20896
rect 36504 20884 36510 20936
rect 24719 20828 25452 20856
rect 24719 20825 24731 20828
rect 24673 20819 24731 20825
rect 35802 20788 35808 20800
rect 24596 20760 35808 20788
rect 35802 20748 35808 20760
rect 35860 20748 35866 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 23198 20584 23204 20596
rect 20588 20556 23204 20584
rect 20588 20544 20594 20556
rect 23198 20544 23204 20556
rect 23256 20544 23262 20596
rect 36814 20544 36820 20596
rect 36872 20584 36878 20596
rect 38105 20587 38163 20593
rect 38105 20584 38117 20587
rect 36872 20556 38117 20584
rect 36872 20544 36878 20556
rect 38105 20553 38117 20556
rect 38151 20553 38163 20587
rect 38105 20547 38163 20553
rect 18046 20476 18052 20528
rect 18104 20516 18110 20528
rect 22830 20516 22836 20528
rect 18104 20488 22836 20516
rect 18104 20476 18110 20488
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 23385 20519 23443 20525
rect 23385 20485 23397 20519
rect 23431 20516 23443 20519
rect 35434 20516 35440 20528
rect 23431 20488 35440 20516
rect 23431 20485 23443 20488
rect 23385 20479 23443 20485
rect 35434 20476 35440 20488
rect 35492 20476 35498 20528
rect 13446 20408 13452 20460
rect 13504 20448 13510 20460
rect 16850 20448 16856 20460
rect 13504 20420 16856 20448
rect 13504 20408 13510 20420
rect 16850 20408 16856 20420
rect 16908 20408 16914 20460
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20448 23535 20451
rect 29638 20448 29644 20460
rect 23523 20420 29644 20448
rect 23523 20417 23535 20420
rect 23477 20411 23535 20417
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 22554 20340 22560 20392
rect 22612 20380 22618 20392
rect 23293 20383 23351 20389
rect 23293 20380 23305 20383
rect 22612 20352 23305 20380
rect 22612 20340 22618 20352
rect 23293 20349 23305 20352
rect 23339 20349 23351 20383
rect 23293 20343 23351 20349
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 23753 20383 23811 20389
rect 23753 20349 23765 20383
rect 23799 20380 23811 20383
rect 24118 20380 24124 20392
rect 23799 20352 24124 20380
rect 23799 20349 23811 20352
rect 23753 20343 23811 20349
rect 21542 20272 21548 20324
rect 21600 20312 21606 20324
rect 23584 20312 23612 20343
rect 24118 20340 24124 20352
rect 24176 20340 24182 20392
rect 37274 20380 37280 20392
rect 37235 20352 37280 20380
rect 37274 20340 37280 20352
rect 37332 20340 37338 20392
rect 37918 20380 37924 20392
rect 37879 20352 37924 20380
rect 37918 20340 37924 20352
rect 37976 20340 37982 20392
rect 21600 20284 23612 20312
rect 21600 20272 21606 20284
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 18230 20244 18236 20256
rect 16816 20216 18236 20244
rect 16816 20204 16822 20216
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 23109 20247 23167 20253
rect 23109 20244 23121 20247
rect 20772 20216 23121 20244
rect 20772 20204 20778 20216
rect 23109 20213 23121 20216
rect 23155 20213 23167 20247
rect 23109 20207 23167 20213
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 37461 20247 37519 20253
rect 37461 20244 37473 20247
rect 26292 20216 37473 20244
rect 26292 20204 26298 20216
rect 37461 20213 37473 20216
rect 37507 20213 37519 20247
rect 37461 20207 37519 20213
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 16574 20040 16580 20052
rect 7800 20012 16580 20040
rect 7800 20000 7806 20012
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17420 20012 19472 20040
rect 1854 19932 1860 19984
rect 1912 19972 1918 19984
rect 16758 19972 16764 19984
rect 1912 19944 16764 19972
rect 1912 19932 1918 19944
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 6886 19876 12434 19904
rect 6270 19796 6276 19848
rect 6328 19836 6334 19848
rect 6886 19836 6914 19876
rect 6328 19808 6914 19836
rect 12406 19836 12434 19876
rect 13170 19864 13176 19916
rect 13228 19904 13234 19916
rect 17420 19913 17448 20012
rect 17494 19932 17500 19984
rect 17552 19972 17558 19984
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 17552 19944 17601 19972
rect 17552 19932 17558 19944
rect 17589 19941 17601 19944
rect 17635 19941 17647 19975
rect 17589 19935 17647 19941
rect 17681 19975 17739 19981
rect 17681 19941 17693 19975
rect 17727 19972 17739 19975
rect 17954 19972 17960 19984
rect 17727 19944 17960 19972
rect 17727 19941 17739 19944
rect 17681 19935 17739 19941
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 13228 19876 17325 19904
rect 13228 19864 13234 19876
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17313 19867 17371 19873
rect 17406 19907 17464 19913
rect 17406 19873 17418 19907
rect 17452 19873 17464 19907
rect 17406 19867 17464 19873
rect 17778 19907 17836 19913
rect 17778 19873 17790 19907
rect 17824 19873 17836 19907
rect 17778 19867 17836 19873
rect 17788 19836 17816 19867
rect 12406 19808 17816 19836
rect 6328 19796 6334 19808
rect 16482 19728 16488 19780
rect 16540 19768 16546 19780
rect 17880 19768 17908 19944
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 19444 19836 19472 20012
rect 19518 19932 19524 19984
rect 19576 19972 19582 19984
rect 20346 19972 20352 19984
rect 19576 19944 20352 19972
rect 19576 19932 19582 19944
rect 20346 19932 20352 19944
rect 20404 19932 20410 19984
rect 27798 19932 27804 19984
rect 27856 19972 27862 19984
rect 36538 19972 36544 19984
rect 27856 19944 36544 19972
rect 27856 19932 27862 19944
rect 36538 19932 36544 19944
rect 36596 19932 36602 19984
rect 20346 19836 20352 19848
rect 19444 19808 20352 19836
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 16540 19740 17908 19768
rect 16540 19728 16546 19740
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 20530 19768 20536 19780
rect 19392 19740 20536 19768
rect 19392 19728 19398 19740
rect 20530 19728 20536 19740
rect 20588 19728 20594 19780
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17494 19700 17500 19712
rect 16816 19672 17500 19700
rect 16816 19660 16822 19672
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 28258 19700 28264 19712
rect 18003 19672 28264 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 28258 19660 28264 19672
rect 28316 19660 28322 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 16758 19496 16764 19508
rect 16408 19468 16764 19496
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 5534 19360 5540 19372
rect 1636 19332 5540 19360
rect 1636 19320 1642 19332
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 1486 19252 1492 19304
rect 1544 19292 1550 19304
rect 2958 19292 2964 19304
rect 1544 19264 2964 19292
rect 1544 19252 1550 19264
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16117 19295 16175 19301
rect 16117 19292 16129 19295
rect 16071 19264 16129 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16117 19261 16129 19264
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 16206 19252 16212 19304
rect 16264 19301 16270 19304
rect 16408 19301 16436 19468
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 18598 19456 18604 19508
rect 18656 19496 18662 19508
rect 21726 19496 21732 19508
rect 18656 19468 21732 19496
rect 18656 19456 18662 19468
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 16482 19388 16488 19440
rect 16540 19388 16546 19440
rect 17310 19428 17316 19440
rect 17057 19400 17316 19428
rect 16500 19301 16528 19388
rect 17057 19360 17085 19400
rect 17310 19388 17316 19400
rect 17368 19388 17374 19440
rect 17586 19428 17592 19440
rect 17499 19400 17592 19428
rect 16960 19332 17085 19360
rect 16264 19295 16295 19301
rect 16283 19261 16295 19295
rect 16264 19255 16295 19261
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19261 16451 19295
rect 16393 19255 16451 19261
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 16582 19295 16640 19301
rect 16582 19261 16594 19295
rect 16628 19261 16640 19295
rect 16582 19255 16640 19261
rect 16264 19252 16270 19255
rect 8938 19184 8944 19236
rect 8996 19224 9002 19236
rect 8996 19196 16160 19224
rect 8996 19184 9002 19196
rect 1581 19159 1639 19165
rect 1581 19125 1593 19159
rect 1627 19156 1639 19159
rect 1762 19156 1768 19168
rect 1627 19128 1768 19156
rect 1627 19125 1639 19128
rect 1581 19119 1639 19125
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 13446 19156 13452 19168
rect 8720 19128 13452 19156
rect 8720 19116 8726 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 16022 19156 16028 19168
rect 15983 19128 16028 19156
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16132 19156 16160 19196
rect 16592 19156 16620 19255
rect 16132 19128 16620 19156
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 16960 19156 16988 19332
rect 17512 19301 17540 19400
rect 17586 19388 17592 19400
rect 17644 19428 17650 19440
rect 18616 19428 18644 19456
rect 17644 19400 18644 19428
rect 17644 19388 17650 19400
rect 17696 19332 17908 19360
rect 17696 19301 17724 19332
rect 17880 19304 17908 19332
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 16807 19128 16988 19156
rect 17144 19264 17233 19292
rect 17144 19156 17172 19264
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17314 19295 17372 19301
rect 17314 19261 17326 19295
rect 17360 19261 17372 19295
rect 17314 19255 17372 19261
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 17686 19295 17744 19301
rect 17686 19261 17698 19295
rect 17732 19261 17744 19295
rect 17686 19255 17744 19261
rect 17218 19156 17224 19168
rect 17144 19128 17224 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 17329 19156 17357 19255
rect 17862 19252 17868 19304
rect 17920 19252 17926 19304
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 19978 19292 19984 19304
rect 19484 19264 19984 19292
rect 19484 19252 19490 19264
rect 19978 19252 19984 19264
rect 20036 19292 20042 19304
rect 21913 19295 21971 19301
rect 21913 19292 21925 19295
rect 20036 19264 21925 19292
rect 20036 19252 20042 19264
rect 21913 19261 21925 19264
rect 21959 19261 21971 19295
rect 21913 19255 21971 19261
rect 22180 19295 22238 19301
rect 22180 19261 22192 19295
rect 22226 19292 22238 19295
rect 23566 19292 23572 19304
rect 22226 19264 23572 19292
rect 22226 19261 22238 19264
rect 22180 19255 22238 19261
rect 23566 19252 23572 19264
rect 23624 19252 23630 19304
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 32766 19292 32772 19304
rect 26936 19264 32772 19292
rect 26936 19252 26942 19264
rect 32766 19252 32772 19264
rect 32824 19252 32830 19304
rect 37274 19292 37280 19304
rect 37235 19264 37280 19292
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 37918 19292 37924 19304
rect 37879 19264 37924 19292
rect 37918 19252 37924 19264
rect 37976 19252 37982 19304
rect 17589 19227 17647 19233
rect 17589 19193 17601 19227
rect 17635 19224 17647 19227
rect 18230 19224 18236 19236
rect 17635 19196 18236 19224
rect 17635 19193 17647 19196
rect 17589 19187 17647 19193
rect 18230 19184 18236 19196
rect 18288 19224 18294 19236
rect 19242 19224 19248 19236
rect 18288 19196 19248 19224
rect 18288 19184 18294 19196
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 20248 19227 20306 19233
rect 20248 19193 20260 19227
rect 20294 19224 20306 19227
rect 24486 19224 24492 19236
rect 20294 19196 24492 19224
rect 20294 19193 20306 19196
rect 20248 19187 20306 19193
rect 24486 19184 24492 19196
rect 24544 19184 24550 19236
rect 36906 19184 36912 19236
rect 36964 19224 36970 19236
rect 36964 19196 38148 19224
rect 36964 19184 36970 19196
rect 17494 19156 17500 19168
rect 17329 19128 17500 19156
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 17865 19159 17923 19165
rect 17865 19125 17877 19159
rect 17911 19156 17923 19159
rect 19978 19156 19984 19168
rect 17911 19128 19984 19156
rect 17911 19125 17923 19128
rect 17865 19119 17923 19125
rect 19978 19116 19984 19128
rect 20036 19116 20042 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21361 19159 21419 19165
rect 21361 19156 21373 19159
rect 20864 19128 21373 19156
rect 20864 19116 20870 19128
rect 21361 19125 21373 19128
rect 21407 19125 21419 19159
rect 23290 19156 23296 19168
rect 23251 19128 23296 19156
rect 21361 19119 21419 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 31386 19116 31392 19168
rect 31444 19156 31450 19168
rect 38120 19165 38148 19196
rect 37461 19159 37519 19165
rect 37461 19156 37473 19159
rect 31444 19128 37473 19156
rect 31444 19116 31450 19128
rect 37461 19125 37473 19128
rect 37507 19125 37519 19159
rect 37461 19119 37519 19125
rect 38105 19159 38163 19165
rect 38105 19125 38117 19159
rect 38151 19125 38163 19159
rect 38105 19119 38163 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 4798 18952 4804 18964
rect 1627 18924 4804 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 17862 18952 17868 18964
rect 16264 18924 17868 18952
rect 16264 18912 16270 18924
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 19061 18955 19119 18961
rect 19061 18952 19073 18955
rect 18472 18924 19073 18952
rect 18472 18912 18478 18924
rect 19061 18921 19073 18924
rect 19107 18921 19119 18955
rect 19242 18952 19248 18964
rect 19155 18924 19248 18952
rect 19061 18915 19119 18921
rect 14458 18844 14464 18896
rect 14516 18884 14522 18896
rect 16117 18887 16175 18893
rect 16117 18884 16129 18887
rect 14516 18856 16129 18884
rect 14516 18844 14522 18856
rect 16117 18853 16129 18856
rect 16163 18853 16175 18887
rect 18230 18884 18236 18896
rect 16117 18847 16175 18853
rect 17696 18856 18236 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 15746 18816 15752 18828
rect 15707 18788 15752 18816
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 15897 18819 15955 18825
rect 15897 18785 15909 18819
rect 15943 18785 15955 18819
rect 15897 18779 15955 18785
rect 15912 18748 15940 18779
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16255 18819 16313 18825
rect 16080 18788 16125 18816
rect 16080 18776 16086 18788
rect 16255 18785 16267 18819
rect 16301 18816 16313 18819
rect 16482 18816 16488 18828
rect 16301 18788 16488 18816
rect 16301 18785 16313 18788
rect 16255 18779 16313 18785
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 16908 18788 17325 18816
rect 16908 18776 16914 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17406 18819 17464 18825
rect 17406 18785 17418 18819
rect 17452 18785 17464 18819
rect 17586 18816 17592 18828
rect 17547 18788 17592 18816
rect 17406 18779 17464 18785
rect 16758 18748 16764 18760
rect 15912 18720 16764 18748
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17420 18748 17448 18779
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 17696 18825 17724 18856
rect 18230 18844 18236 18856
rect 18288 18844 18294 18896
rect 18598 18844 18604 18896
rect 18656 18884 18662 18896
rect 18693 18887 18751 18893
rect 18693 18884 18705 18887
rect 18656 18856 18705 18884
rect 18656 18844 18662 18856
rect 18693 18853 18705 18856
rect 18739 18853 18751 18887
rect 18693 18847 18751 18853
rect 18785 18887 18843 18893
rect 18785 18853 18797 18887
rect 18831 18884 18843 18887
rect 19168 18884 19196 18924
rect 19242 18912 19248 18924
rect 19300 18952 19306 18964
rect 20622 18952 20628 18964
rect 19300 18924 20628 18952
rect 19300 18912 19306 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 24946 18952 24952 18964
rect 20864 18924 24952 18952
rect 20864 18912 20870 18924
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 36998 18912 37004 18964
rect 37056 18952 37062 18964
rect 37369 18955 37427 18961
rect 37369 18952 37381 18955
rect 37056 18924 37381 18952
rect 37056 18912 37062 18924
rect 37369 18921 37381 18924
rect 37415 18921 37427 18955
rect 37369 18915 37427 18921
rect 18831 18856 19196 18884
rect 18831 18853 18843 18856
rect 18785 18847 18843 18853
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 25130 18884 25136 18896
rect 20036 18856 25136 18884
rect 20036 18844 20042 18856
rect 25130 18844 25136 18856
rect 25188 18844 25194 18896
rect 28166 18844 28172 18896
rect 28224 18884 28230 18896
rect 29178 18884 29184 18896
rect 28224 18856 29184 18884
rect 28224 18844 28230 18856
rect 29178 18844 29184 18856
rect 29236 18844 29242 18896
rect 17689 18819 17747 18825
rect 17689 18785 17701 18819
rect 17735 18785 17747 18819
rect 17689 18779 17747 18785
rect 17819 18819 17877 18825
rect 17819 18785 17831 18819
rect 17865 18816 17877 18819
rect 18414 18816 18420 18828
rect 17865 18785 17897 18816
rect 18375 18788 18420 18816
rect 17819 18779 17897 18785
rect 17276 18720 17448 18748
rect 17869 18748 17897 18779
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 18510 18819 18568 18825
rect 18510 18785 18522 18819
rect 18556 18785 18568 18819
rect 18510 18779 18568 18785
rect 18882 18819 18940 18825
rect 18882 18785 18894 18819
rect 18928 18785 18940 18819
rect 18882 18779 18940 18785
rect 17954 18748 17960 18760
rect 17869 18720 17960 18748
rect 17276 18708 17282 18720
rect 17954 18708 17960 18720
rect 18012 18708 18018 18760
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18524 18748 18552 18779
rect 18380 18720 18552 18748
rect 18380 18708 18386 18720
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 18892 18748 18920 18779
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19484 18788 19533 18816
rect 19484 18776 19490 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 19788 18819 19846 18825
rect 19788 18785 19800 18819
rect 19834 18816 19846 18819
rect 20714 18816 20720 18828
rect 19834 18788 20720 18816
rect 19834 18785 19846 18788
rect 19788 18779 19846 18785
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 37182 18816 37188 18828
rect 37143 18788 37188 18816
rect 37182 18776 37188 18788
rect 37240 18776 37246 18828
rect 21634 18748 21640 18760
rect 18656 18720 18920 18748
rect 20548 18720 21640 18748
rect 18656 18708 18662 18720
rect 19518 18680 19524 18692
rect 17880 18652 19524 18680
rect 16393 18615 16451 18621
rect 16393 18581 16405 18615
rect 16439 18612 16451 18615
rect 17880 18612 17908 18652
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 16439 18584 17908 18612
rect 17957 18615 18015 18621
rect 16439 18581 16451 18584
rect 16393 18575 16451 18581
rect 17957 18581 17969 18615
rect 18003 18612 18015 18615
rect 20548 18612 20576 18720
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 27982 18708 27988 18760
rect 28040 18748 28046 18760
rect 36998 18748 37004 18760
rect 28040 18720 37004 18748
rect 28040 18708 28046 18720
rect 36998 18708 37004 18720
rect 37056 18708 37062 18760
rect 21450 18640 21456 18692
rect 21508 18680 21514 18692
rect 37642 18680 37648 18692
rect 21508 18652 37648 18680
rect 21508 18640 21514 18652
rect 37642 18640 37648 18652
rect 37700 18640 37706 18692
rect 18003 18584 20576 18612
rect 20901 18615 20959 18621
rect 18003 18581 18015 18584
rect 17957 18575 18015 18581
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21542 18612 21548 18624
rect 20947 18584 21548 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21542 18572 21548 18584
rect 21600 18572 21606 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 13262 18368 13268 18420
rect 13320 18408 13326 18420
rect 17954 18408 17960 18420
rect 13320 18380 17960 18408
rect 13320 18368 13326 18380
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 18785 18411 18843 18417
rect 18785 18377 18797 18411
rect 18831 18408 18843 18411
rect 19334 18408 19340 18420
rect 18831 18380 19340 18408
rect 18831 18377 18843 18380
rect 18785 18371 18843 18377
rect 19334 18368 19340 18380
rect 19392 18408 19398 18420
rect 20714 18408 20720 18420
rect 19392 18380 20720 18408
rect 19392 18368 19398 18380
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 21542 18368 21548 18420
rect 21600 18408 21606 18420
rect 23842 18408 23848 18420
rect 21600 18380 23848 18408
rect 21600 18368 21606 18380
rect 23842 18368 23848 18380
rect 23900 18368 23906 18420
rect 38105 18411 38163 18417
rect 38105 18377 38117 18411
rect 38151 18408 38163 18411
rect 38194 18408 38200 18420
rect 38151 18380 38200 18408
rect 38151 18377 38163 18380
rect 38105 18371 38163 18377
rect 38194 18368 38200 18380
rect 38252 18368 38258 18420
rect 17586 18340 17592 18352
rect 16868 18312 17592 18340
rect 4798 18232 4804 18284
rect 4856 18272 4862 18284
rect 4856 18244 9674 18272
rect 4856 18232 4862 18244
rect 9646 18068 9674 18244
rect 16574 18204 16580 18216
rect 16535 18176 16580 18204
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 16758 18213 16764 18216
rect 16725 18207 16764 18213
rect 16725 18173 16737 18207
rect 16725 18167 16764 18173
rect 16758 18164 16764 18167
rect 16816 18164 16822 18216
rect 16868 18213 16896 18312
rect 17586 18300 17592 18312
rect 17644 18300 17650 18352
rect 18230 18272 18236 18284
rect 16960 18244 18236 18272
rect 16960 18213 16988 18244
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19484 18244 19993 18272
rect 19484 18232 19490 18244
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 17042 18207 17100 18213
rect 17042 18173 17054 18207
rect 17088 18173 17100 18207
rect 17042 18167 17100 18173
rect 17057 18068 17085 18167
rect 17770 18164 17776 18216
rect 17828 18204 17834 18216
rect 17957 18207 18015 18213
rect 17957 18204 17969 18207
rect 17828 18176 17969 18204
rect 17828 18164 17834 18176
rect 17957 18173 17969 18176
rect 18003 18173 18015 18207
rect 18874 18204 18880 18216
rect 18835 18176 18880 18204
rect 17957 18167 18015 18173
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 20248 18207 20306 18213
rect 20248 18173 20260 18207
rect 20294 18204 20306 18207
rect 24394 18204 24400 18216
rect 20294 18176 24400 18204
rect 20294 18173 20306 18176
rect 20248 18167 20306 18173
rect 24394 18164 24400 18176
rect 24452 18164 24458 18216
rect 26050 18204 26056 18216
rect 24504 18176 26056 18204
rect 17236 18108 22094 18136
rect 17236 18077 17264 18108
rect 9646 18040 17085 18068
rect 17221 18071 17279 18077
rect 17221 18037 17233 18071
rect 17267 18037 17279 18071
rect 17221 18031 17279 18037
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21542 18068 21548 18080
rect 21407 18040 21548 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 22066 18068 22094 18108
rect 24504 18068 24532 18176
rect 26050 18164 26056 18176
rect 26108 18164 26114 18216
rect 37918 18204 37924 18216
rect 37879 18176 37924 18204
rect 37918 18164 37924 18176
rect 37976 18164 37982 18216
rect 25406 18096 25412 18148
rect 25464 18136 25470 18148
rect 28074 18136 28080 18148
rect 25464 18108 28080 18136
rect 25464 18096 25470 18108
rect 28074 18096 28080 18108
rect 28132 18096 28138 18148
rect 22066 18040 24532 18068
rect 25314 18028 25320 18080
rect 25372 18068 25378 18080
rect 27706 18068 27712 18080
rect 25372 18040 27712 18068
rect 25372 18028 25378 18040
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 34422 18028 34428 18080
rect 34480 18068 34486 18080
rect 36078 18068 36084 18080
rect 34480 18040 36084 18068
rect 34480 18028 34486 18040
rect 36078 18028 36084 18040
rect 36136 18028 36142 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1670 17864 1676 17876
rect 1627 17836 1676 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 8386 17864 8392 17876
rect 7524 17836 8392 17864
rect 7524 17824 7530 17836
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 17957 17867 18015 17873
rect 17957 17833 17969 17867
rect 18003 17833 18015 17867
rect 17957 17827 18015 17833
rect 17586 17796 17592 17808
rect 17547 17768 17592 17796
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 17681 17799 17739 17805
rect 17681 17765 17693 17799
rect 17727 17796 17739 17799
rect 17972 17796 18000 17827
rect 18322 17824 18328 17876
rect 18380 17864 18386 17876
rect 18380 17836 26234 17864
rect 18380 17824 18386 17836
rect 17727 17768 17909 17796
rect 17972 17768 22094 17796
rect 17727 17765 17739 17768
rect 17681 17759 17739 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1670 17688 1676 17740
rect 1728 17728 1734 17740
rect 5718 17728 5724 17740
rect 1728 17700 5724 17728
rect 1728 17688 1734 17700
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 11756 17700 17325 17728
rect 11756 17688 11762 17700
rect 17313 17697 17325 17700
rect 17359 17697 17371 17731
rect 17313 17691 17371 17697
rect 17461 17731 17519 17737
rect 17461 17697 17473 17731
rect 17507 17697 17519 17731
rect 17778 17731 17836 17737
rect 17778 17728 17790 17731
rect 17461 17691 17519 17697
rect 17604 17700 17790 17728
rect 17476 17592 17504 17691
rect 17604 17672 17632 17700
rect 17778 17697 17790 17700
rect 17824 17697 17836 17731
rect 17881 17728 17909 17768
rect 18230 17728 18236 17740
rect 17881 17700 18236 17728
rect 17778 17691 17836 17697
rect 18230 17688 18236 17700
rect 18288 17688 18294 17740
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19797 17731 19855 17737
rect 19797 17728 19809 17731
rect 19484 17700 19809 17728
rect 19484 17688 19490 17700
rect 19797 17697 19809 17700
rect 19843 17697 19855 17731
rect 19797 17691 19855 17697
rect 20064 17731 20122 17737
rect 20064 17697 20076 17731
rect 20110 17728 20122 17731
rect 21358 17728 21364 17740
rect 20110 17700 21364 17728
rect 20110 17697 20122 17700
rect 20064 17691 20122 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 22066 17728 22094 17768
rect 22922 17756 22928 17808
rect 22980 17796 22986 17808
rect 25958 17796 25964 17808
rect 22980 17768 25964 17796
rect 22980 17756 22986 17768
rect 25958 17756 25964 17768
rect 26016 17756 26022 17808
rect 26206 17796 26234 17836
rect 28258 17824 28264 17876
rect 28316 17864 28322 17876
rect 29086 17864 29092 17876
rect 28316 17836 29092 17864
rect 28316 17824 28322 17836
rect 29086 17824 29092 17836
rect 29144 17824 29150 17876
rect 32858 17824 32864 17876
rect 32916 17864 32922 17876
rect 37369 17867 37427 17873
rect 37369 17864 37381 17867
rect 32916 17836 37381 17864
rect 32916 17824 32922 17836
rect 37369 17833 37381 17836
rect 37415 17833 37427 17867
rect 37369 17827 37427 17833
rect 37458 17796 37464 17808
rect 26206 17768 37464 17796
rect 37458 17756 37464 17768
rect 37516 17756 37522 17808
rect 24302 17728 24308 17740
rect 22066 17700 24308 17728
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 29638 17688 29644 17740
rect 29696 17728 29702 17740
rect 33686 17728 33692 17740
rect 29696 17700 33692 17728
rect 29696 17688 29702 17700
rect 33686 17688 33692 17700
rect 33744 17688 33750 17740
rect 37182 17728 37188 17740
rect 37143 17700 37188 17728
rect 37182 17688 37188 17700
rect 37240 17688 37246 17740
rect 17586 17620 17592 17672
rect 17644 17620 17650 17672
rect 18414 17592 18420 17604
rect 17476 17564 18420 17592
rect 18414 17552 18420 17564
rect 18472 17552 18478 17604
rect 21726 17592 21732 17604
rect 21100 17564 21732 17592
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 17310 17524 17316 17536
rect 9180 17496 17316 17524
rect 9180 17484 9186 17496
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 18874 17484 18880 17536
rect 18932 17524 18938 17536
rect 21100 17524 21128 17564
rect 21726 17552 21732 17564
rect 21784 17552 21790 17604
rect 18932 17496 21128 17524
rect 21177 17527 21235 17533
rect 18932 17484 18938 17496
rect 21177 17493 21189 17527
rect 21223 17524 21235 17527
rect 21358 17524 21364 17536
rect 21223 17496 21364 17524
rect 21223 17493 21235 17496
rect 21177 17487 21235 17493
rect 21358 17484 21364 17496
rect 21416 17524 21422 17536
rect 21818 17524 21824 17536
rect 21416 17496 21824 17524
rect 21416 17484 21422 17496
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 17586 17320 17592 17332
rect 14424 17292 17592 17320
rect 14424 17280 14430 17292
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 21266 17320 21272 17332
rect 21227 17292 21272 17320
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 21376 17292 31064 17320
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 16574 17252 16580 17264
rect 8352 17224 16580 17252
rect 8352 17212 8358 17224
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 16758 17212 16764 17264
rect 16816 17252 16822 17264
rect 21376 17252 21404 17292
rect 16816 17224 21404 17252
rect 21468 17224 26234 17252
rect 16816 17212 16822 17224
rect 2038 17144 2044 17196
rect 2096 17184 2102 17196
rect 4798 17184 4804 17196
rect 2096 17156 4804 17184
rect 2096 17144 2102 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 21468 17184 21496 17224
rect 23382 17184 23388 17196
rect 17552 17156 21496 17184
rect 21560 17156 23388 17184
rect 17552 17144 17558 17156
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 21560 17125 21588 17156
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20956 17088 21465 17116
rect 20956 17076 20962 17088
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 21545 17119 21603 17125
rect 21545 17085 21557 17119
rect 21591 17085 21603 17119
rect 21545 17079 21603 17085
rect 21726 17076 21732 17128
rect 21784 17125 21790 17128
rect 21784 17119 21813 17125
rect 21801 17085 21813 17119
rect 21784 17079 21813 17085
rect 21913 17119 21971 17125
rect 21913 17085 21925 17119
rect 21959 17116 21971 17119
rect 21959 17088 22094 17116
rect 21959 17085 21971 17088
rect 21913 17079 21971 17085
rect 21784 17076 21790 17079
rect 19334 17008 19340 17060
rect 19392 17048 19398 17060
rect 21637 17051 21695 17057
rect 21637 17048 21649 17051
rect 19392 17020 21649 17048
rect 19392 17008 19398 17020
rect 21637 17017 21649 17020
rect 21683 17017 21695 17051
rect 22066 17048 22094 17088
rect 22462 17048 22468 17060
rect 22066 17020 22468 17048
rect 21637 17011 21695 17017
rect 22462 17008 22468 17020
rect 22520 17048 22526 17060
rect 23014 17048 23020 17060
rect 22520 17020 23020 17048
rect 22520 17008 22526 17020
rect 23014 17008 23020 17020
rect 23072 17008 23078 17060
rect 26206 17048 26234 17224
rect 31036 17184 31064 17292
rect 36722 17280 36728 17332
rect 36780 17320 36786 17332
rect 37461 17323 37519 17329
rect 37461 17320 37473 17323
rect 36780 17292 37473 17320
rect 36780 17280 36786 17292
rect 37461 17289 37473 17292
rect 37507 17289 37519 17323
rect 37461 17283 37519 17289
rect 34330 17212 34336 17264
rect 34388 17252 34394 17264
rect 38105 17255 38163 17261
rect 38105 17252 38117 17255
rect 34388 17224 38117 17252
rect 34388 17212 34394 17224
rect 38105 17221 38117 17224
rect 38151 17221 38163 17255
rect 38105 17215 38163 17221
rect 37090 17184 37096 17196
rect 31036 17156 37096 17184
rect 37090 17144 37096 17156
rect 37148 17144 37154 17196
rect 37274 17116 37280 17128
rect 37235 17088 37280 17116
rect 37274 17076 37280 17088
rect 37332 17076 37338 17128
rect 37918 17116 37924 17128
rect 37879 17088 37924 17116
rect 37918 17076 37924 17088
rect 37976 17076 37982 17128
rect 37366 17048 37372 17060
rect 26206 17020 37372 17048
rect 37366 17008 37372 17020
rect 37424 17008 37430 17060
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21450 16980 21456 16992
rect 20956 16952 21456 16980
rect 20956 16940 20962 16952
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 13446 16736 13452 16788
rect 13504 16776 13510 16788
rect 18598 16776 18604 16788
rect 13504 16748 18604 16776
rect 13504 16736 13510 16748
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 21358 16776 21364 16788
rect 20128 16748 21364 16776
rect 20128 16736 20134 16748
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 22922 16736 22928 16788
rect 22980 16776 22986 16788
rect 28350 16776 28356 16788
rect 22980 16748 28356 16776
rect 22980 16736 22986 16748
rect 28350 16736 28356 16748
rect 28408 16736 28414 16788
rect 36998 16736 37004 16788
rect 37056 16776 37062 16788
rect 37277 16779 37335 16785
rect 37277 16776 37289 16779
rect 37056 16748 37289 16776
rect 37056 16736 37062 16748
rect 37277 16745 37289 16748
rect 37323 16745 37335 16779
rect 37277 16739 37335 16745
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 9398 16708 9404 16720
rect 5868 16680 9404 16708
rect 5868 16668 5874 16680
rect 9398 16668 9404 16680
rect 9456 16668 9462 16720
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 28442 16640 28448 16652
rect 24360 16612 28448 16640
rect 24360 16600 24366 16612
rect 28442 16600 28448 16612
rect 28500 16600 28506 16652
rect 37182 16640 37188 16652
rect 37143 16612 37188 16640
rect 37182 16600 37188 16612
rect 37240 16600 37246 16652
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1544 16204 1593 16232
rect 1544 16192 1550 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 22002 16192 22008 16244
rect 22060 16232 22066 16244
rect 22060 16204 26234 16232
rect 22060 16192 22066 16204
rect 17221 16167 17279 16173
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 24026 16164 24032 16176
rect 17267 16136 24032 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 24026 16124 24032 16136
rect 24084 16124 24090 16176
rect 26206 16096 26234 16204
rect 35526 16192 35532 16244
rect 35584 16232 35590 16244
rect 37461 16235 37519 16241
rect 37461 16232 37473 16235
rect 35584 16204 37473 16232
rect 35584 16192 35590 16204
rect 37461 16201 37473 16204
rect 37507 16201 37519 16235
rect 37461 16195 37519 16201
rect 32214 16124 32220 16176
rect 32272 16164 32278 16176
rect 38105 16167 38163 16173
rect 38105 16164 38117 16167
rect 32272 16136 38117 16164
rect 32272 16124 32278 16136
rect 38105 16133 38117 16136
rect 38151 16133 38163 16167
rect 38105 16127 38163 16133
rect 37826 16096 37832 16108
rect 16960 16068 22094 16096
rect 26206 16068 37832 16096
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 16574 16028 16580 16040
rect 16535 16000 16580 16028
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16725 16031 16783 16037
rect 16725 15997 16737 16031
rect 16771 16028 16783 16031
rect 16960 16028 16988 16068
rect 16771 16000 16988 16028
rect 17042 16031 17100 16037
rect 16771 15997 16783 16000
rect 16725 15991 16783 15997
rect 17042 15997 17054 16031
rect 17088 16028 17100 16031
rect 22066 16028 22094 16068
rect 37826 16056 37832 16068
rect 37884 16056 37890 16108
rect 35250 16028 35256 16040
rect 17088 16000 17264 16028
rect 22066 16000 35256 16028
rect 17088 15997 17100 16000
rect 17042 15991 17100 15997
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 16850 15960 16856 15972
rect 1820 15932 6914 15960
rect 16811 15932 16856 15960
rect 1820 15920 1826 15932
rect 6886 15892 6914 15932
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 16945 15963 17003 15969
rect 16945 15929 16957 15963
rect 16991 15960 17003 15963
rect 17126 15960 17132 15972
rect 16991 15932 17132 15960
rect 16991 15929 17003 15932
rect 16945 15923 17003 15929
rect 17126 15920 17132 15932
rect 17184 15920 17190 15972
rect 17236 15892 17264 16000
rect 35250 15988 35256 16000
rect 35308 15988 35314 16040
rect 37274 16028 37280 16040
rect 37235 16000 37280 16028
rect 37274 15988 37280 16000
rect 37332 15988 37338 16040
rect 37918 16028 37924 16040
rect 37879 16000 37924 16028
rect 37918 15988 37924 16000
rect 37976 15988 37982 16040
rect 18414 15920 18420 15972
rect 18472 15960 18478 15972
rect 36170 15960 36176 15972
rect 18472 15932 36176 15960
rect 18472 15920 18478 15932
rect 36170 15920 36176 15932
rect 36228 15920 36234 15972
rect 6886 15864 17264 15892
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 1670 15688 1676 15700
rect 1627 15660 1676 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 17957 15691 18015 15697
rect 8260 15660 17816 15688
rect 8260 15648 8266 15660
rect 12342 15580 12348 15632
rect 12400 15620 12406 15632
rect 17126 15620 17132 15632
rect 12400 15592 16252 15620
rect 12400 15580 12406 15592
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 14918 15512 14924 15564
rect 14976 15552 14982 15564
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 14976 15524 15761 15552
rect 14976 15512 14982 15524
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 15838 15512 15844 15564
rect 15896 15552 15902 15564
rect 16224 15561 16252 15592
rect 16316 15592 17132 15620
rect 16025 15555 16083 15561
rect 15896 15524 15941 15552
rect 15896 15512 15902 15524
rect 16025 15521 16037 15555
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 16214 15555 16272 15561
rect 16214 15521 16226 15555
rect 16260 15521 16272 15555
rect 16214 15515 16272 15521
rect 16040 15416 16068 15515
rect 16132 15484 16160 15515
rect 16316 15484 16344 15592
rect 17126 15580 17132 15592
rect 17184 15620 17190 15632
rect 17681 15623 17739 15629
rect 17681 15620 17693 15623
rect 17184 15592 17693 15620
rect 17184 15580 17190 15592
rect 17681 15589 17693 15592
rect 17727 15589 17739 15623
rect 17681 15583 17739 15589
rect 17310 15552 17316 15564
rect 17271 15524 17316 15552
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 17494 15561 17500 15564
rect 17461 15555 17500 15561
rect 17461 15521 17473 15555
rect 17461 15515 17500 15521
rect 17494 15512 17500 15515
rect 17552 15512 17558 15564
rect 17586 15512 17592 15564
rect 17644 15552 17650 15564
rect 17788 15561 17816 15660
rect 17957 15657 17969 15691
rect 18003 15688 18015 15691
rect 24670 15688 24676 15700
rect 18003 15660 24676 15688
rect 18003 15657 18015 15660
rect 17957 15651 18015 15657
rect 24670 15648 24676 15660
rect 24728 15648 24734 15700
rect 36538 15648 36544 15700
rect 36596 15688 36602 15700
rect 37277 15691 37335 15697
rect 37277 15688 37289 15691
rect 36596 15660 37289 15688
rect 36596 15648 36602 15660
rect 37277 15657 37289 15660
rect 37323 15657 37335 15691
rect 37277 15651 37335 15657
rect 17778 15555 17836 15561
rect 17644 15524 17689 15552
rect 17644 15512 17650 15524
rect 17778 15521 17790 15555
rect 17824 15521 17836 15555
rect 37182 15552 37188 15564
rect 37143 15524 37188 15552
rect 17778 15515 17836 15521
rect 37182 15512 37188 15524
rect 37240 15512 37246 15564
rect 16132 15456 16344 15484
rect 16850 15444 16856 15496
rect 16908 15484 16914 15496
rect 17604 15484 17632 15512
rect 16908 15456 17632 15484
rect 16908 15444 16914 15456
rect 16393 15419 16451 15425
rect 16040 15388 16160 15416
rect 16132 15348 16160 15388
rect 16393 15385 16405 15419
rect 16439 15416 16451 15419
rect 24578 15416 24584 15428
rect 16439 15388 24584 15416
rect 16439 15385 16451 15388
rect 16393 15379 16451 15385
rect 24578 15376 24584 15388
rect 24636 15376 24642 15428
rect 16850 15348 16856 15360
rect 16132 15320 16856 15348
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 17129 15147 17187 15153
rect 12406 15116 16988 15144
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 12406 15008 12434 15116
rect 8444 14980 12434 15008
rect 16960 15008 16988 15116
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 18233 15147 18291 15153
rect 17175 15116 18184 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 17678 15036 17684 15088
rect 17736 15036 17742 15088
rect 18156 15076 18184 15116
rect 18233 15113 18245 15147
rect 18279 15144 18291 15147
rect 22554 15144 22560 15156
rect 18279 15116 22560 15144
rect 18279 15113 18291 15116
rect 18233 15107 18291 15113
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 35618 15104 35624 15156
rect 35676 15144 35682 15156
rect 37461 15147 37519 15153
rect 37461 15144 37473 15147
rect 35676 15116 37473 15144
rect 35676 15104 35682 15116
rect 37461 15113 37473 15116
rect 37507 15113 37519 15147
rect 37461 15107 37519 15113
rect 23474 15076 23480 15088
rect 18156 15048 23480 15076
rect 23474 15036 23480 15048
rect 23532 15036 23538 15088
rect 35710 15036 35716 15088
rect 35768 15076 35774 15088
rect 38105 15079 38163 15085
rect 38105 15076 38117 15079
rect 35768 15048 38117 15076
rect 35768 15036 35774 15048
rect 38105 15045 38117 15048
rect 38151 15045 38163 15079
rect 38105 15039 38163 15045
rect 17696 15008 17724 15036
rect 16960 14980 17632 15008
rect 17696 14980 17908 15008
rect 8444 14968 8450 14980
rect 14550 14900 14556 14952
rect 14608 14940 14614 14952
rect 16485 14943 16543 14949
rect 16485 14940 16497 14943
rect 14608 14912 16497 14940
rect 14608 14900 14614 14912
rect 16485 14909 16497 14912
rect 16531 14909 16543 14943
rect 16485 14903 16543 14909
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16758 14940 16764 14952
rect 16632 14912 16677 14940
rect 16719 14912 16764 14940
rect 16632 14900 16638 14912
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 17034 14949 17040 14952
rect 16991 14943 17040 14949
rect 16991 14909 17003 14943
rect 17037 14909 17040 14943
rect 16991 14903 17040 14909
rect 17034 14900 17040 14903
rect 17092 14900 17098 14952
rect 17604 14949 17632 14980
rect 17589 14943 17647 14949
rect 17589 14909 17601 14943
rect 17635 14909 17647 14943
rect 17589 14903 17647 14909
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 17880 14949 17908 14980
rect 19150 14968 19156 15020
rect 19208 15008 19214 15020
rect 24946 15008 24952 15020
rect 19208 14980 24952 15008
rect 19208 14968 19214 14980
rect 24946 14968 24952 14980
rect 25004 14968 25010 15020
rect 17865 14943 17923 14949
rect 17736 14912 17781 14940
rect 17736 14900 17742 14912
rect 17865 14909 17877 14943
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 18046 14900 18052 14952
rect 18104 14949 18110 14952
rect 18104 14940 18112 14949
rect 37274 14940 37280 14952
rect 18104 14912 18149 14940
rect 37235 14912 37280 14940
rect 18104 14903 18112 14912
rect 18104 14900 18110 14903
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 37918 14940 37924 14952
rect 37879 14912 37924 14940
rect 37918 14900 37924 14912
rect 37976 14900 37982 14952
rect 16853 14875 16911 14881
rect 6886 14844 9674 14872
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 6886 14804 6914 14844
rect 3568 14776 6914 14804
rect 9646 14804 9674 14844
rect 16853 14841 16865 14875
rect 16899 14872 16911 14875
rect 17126 14872 17132 14884
rect 16899 14844 17132 14872
rect 16899 14841 16911 14844
rect 16853 14835 16911 14841
rect 17126 14832 17132 14844
rect 17184 14872 17190 14884
rect 17957 14875 18015 14881
rect 17957 14872 17969 14875
rect 17184 14844 17969 14872
rect 17184 14832 17190 14844
rect 17957 14841 17969 14844
rect 18003 14841 18015 14875
rect 17957 14835 18015 14841
rect 17034 14804 17040 14816
rect 9646 14776 17040 14804
rect 3568 14764 3574 14776
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 7558 14600 7564 14612
rect 1627 14572 7564 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 37274 14600 37280 14612
rect 20036 14572 37280 14600
rect 20036 14560 20042 14572
rect 37274 14560 37280 14572
rect 37332 14560 37338 14612
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 38010 14532 38016 14544
rect 16080 14504 38016 14532
rect 16080 14492 16086 14504
rect 38010 14492 38016 14504
rect 38068 14492 38074 14544
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 24854 14464 24860 14476
rect 16632 14436 24860 14464
rect 16632 14424 16638 14436
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 25866 14424 25872 14476
rect 25924 14464 25930 14476
rect 28997 14467 29055 14473
rect 28997 14464 29009 14467
rect 25924 14436 29009 14464
rect 25924 14424 25930 14436
rect 28997 14433 29009 14436
rect 29043 14433 29055 14467
rect 28997 14427 29055 14433
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 18046 14396 18052 14408
rect 6420 14368 18052 14396
rect 6420 14356 6426 14368
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 29181 14263 29239 14269
rect 29181 14229 29193 14263
rect 29227 14260 29239 14263
rect 34514 14260 34520 14272
rect 29227 14232 34520 14260
rect 29227 14229 29239 14232
rect 29181 14223 29239 14229
rect 34514 14220 34520 14232
rect 34572 14220 34578 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 3602 14056 3608 14068
rect 1627 14028 3608 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 32490 14016 32496 14068
rect 32548 14056 32554 14068
rect 37277 14059 37335 14065
rect 37277 14056 37289 14059
rect 32548 14028 37289 14056
rect 32548 14016 32554 14028
rect 37277 14025 37289 14028
rect 37323 14025 37335 14059
rect 37277 14019 37335 14025
rect 25958 13948 25964 14000
rect 26016 13988 26022 14000
rect 38105 13991 38163 13997
rect 38105 13988 38117 13991
rect 26016 13960 38117 13988
rect 26016 13948 26022 13960
rect 38105 13957 38117 13960
rect 38151 13957 38163 13991
rect 38105 13951 38163 13957
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 37182 13852 37188 13864
rect 37143 13824 37188 13852
rect 37182 13812 37188 13824
rect 37240 13812 37246 13864
rect 37918 13852 37924 13864
rect 37879 13824 37924 13852
rect 37918 13812 37924 13824
rect 37976 13812 37982 13864
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 16390 13784 16396 13796
rect 15344 13756 16396 13784
rect 15344 13744 15350 13756
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 21818 13472 21824 13524
rect 21876 13512 21882 13524
rect 26326 13512 26332 13524
rect 21876 13484 26332 13512
rect 21876 13472 21882 13484
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 37182 13376 37188 13388
rect 37143 13348 37188 13376
rect 37182 13336 37188 13348
rect 37240 13336 37246 13388
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 19334 13308 19340 13320
rect 10468 13280 19340 13308
rect 10468 13268 10474 13280
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 17862 13200 17868 13252
rect 17920 13240 17926 13252
rect 36906 13240 36912 13252
rect 17920 13212 36912 13240
rect 17920 13200 17926 13212
rect 36906 13200 36912 13212
rect 36964 13200 36970 13252
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 14366 13172 14372 13184
rect 1820 13144 14372 13172
rect 1820 13132 1826 13144
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 37277 13175 37335 13181
rect 37277 13172 37289 13175
rect 21968 13144 37289 13172
rect 21968 13132 21974 13144
rect 37277 13141 37289 13144
rect 37323 13141 37335 13175
rect 37277 13135 37335 13141
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 6454 12968 6460 12980
rect 1627 12940 6460 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 38013 12971 38071 12977
rect 38013 12968 38025 12971
rect 29788 12940 38025 12968
rect 29788 12928 29794 12940
rect 38013 12937 38025 12940
rect 38059 12937 38071 12971
rect 38013 12931 38071 12937
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20772 12804 21005 12832
rect 20772 12792 20778 12804
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 21361 12767 21419 12773
rect 21361 12764 21373 12767
rect 20680 12736 21373 12764
rect 20680 12724 20686 12736
rect 21361 12733 21373 12736
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 21453 12699 21511 12705
rect 21453 12696 21465 12699
rect 16448 12668 21465 12696
rect 16448 12656 16454 12668
rect 21453 12665 21465 12668
rect 21499 12665 21511 12699
rect 21726 12696 21732 12708
rect 21687 12668 21732 12696
rect 21453 12659 21511 12665
rect 21726 12656 21732 12668
rect 21784 12656 21790 12708
rect 37918 12696 37924 12708
rect 37879 12668 37924 12696
rect 37918 12656 37924 12668
rect 37976 12656 37982 12708
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20588 12600 21281 12628
rect 20588 12588 20594 12600
rect 21269 12597 21281 12600
rect 21315 12597 21327 12631
rect 21269 12591 21327 12597
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1854 12424 1860 12436
rect 1627 12396 1860 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 36630 12384 36636 12436
rect 36688 12424 36694 12436
rect 37277 12427 37335 12433
rect 37277 12424 37289 12427
rect 36688 12396 37289 12424
rect 36688 12384 36694 12396
rect 37277 12393 37289 12396
rect 37323 12393 37335 12427
rect 37277 12387 37335 12393
rect 19886 12316 19892 12368
rect 19944 12356 19950 12368
rect 20530 12356 20536 12368
rect 19944 12328 20536 12356
rect 19944 12316 19950 12328
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 37182 12288 37188 12300
rect 37143 12260 37188 12288
rect 37182 12248 37188 12260
rect 37240 12248 37246 12300
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 20806 11880 20812 11892
rect 10284 11852 20812 11880
rect 10284 11840 10290 11852
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 31110 11840 31116 11892
rect 31168 11880 31174 11892
rect 38013 11883 38071 11889
rect 38013 11880 38025 11883
rect 31168 11852 38025 11880
rect 31168 11840 31174 11852
rect 38013 11849 38025 11852
rect 38059 11849 38071 11883
rect 38013 11843 38071 11849
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 36262 11812 36268 11824
rect 17552 11784 36268 11812
rect 17552 11772 17558 11784
rect 36262 11772 36268 11784
rect 36320 11772 36326 11824
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 10502 11744 10508 11756
rect 4120 11716 10508 11744
rect 4120 11704 4126 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 36722 11744 36728 11756
rect 16172 11716 36728 11744
rect 16172 11704 16178 11716
rect 36722 11704 36728 11716
rect 36780 11704 36786 11756
rect 37182 11676 37188 11688
rect 37143 11648 37188 11676
rect 37182 11636 37188 11648
rect 37240 11636 37246 11688
rect 37918 11608 37924 11620
rect 37879 11580 37924 11608
rect 37918 11568 37924 11580
rect 37976 11568 37982 11620
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 37277 11543 37335 11549
rect 37277 11540 37289 11543
rect 19024 11512 37289 11540
rect 19024 11500 19030 11512
rect 37277 11509 37289 11512
rect 37323 11509 37335 11543
rect 37277 11503 37335 11509
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 37182 11200 37188 11212
rect 37143 11172 37188 11200
rect 37182 11160 37188 11172
rect 37240 11160 37246 11212
rect 17126 11092 17132 11144
rect 17184 11132 17190 11144
rect 19886 11132 19892 11144
rect 17184 11104 19892 11132
rect 17184 11092 17190 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 20312 11104 31754 11132
rect 20312 11092 20318 11104
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 10594 11064 10600 11076
rect 1627 11036 10600 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 18782 11064 18788 11076
rect 12952 11036 18788 11064
rect 12952 11024 12958 11036
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 21726 11024 21732 11076
rect 21784 11064 21790 11076
rect 25958 11064 25964 11076
rect 21784 11036 25964 11064
rect 21784 11024 21790 11036
rect 25958 11024 25964 11036
rect 26016 11024 26022 11076
rect 31726 11064 31754 11104
rect 37369 11067 37427 11073
rect 37369 11064 37381 11067
rect 31726 11036 37381 11064
rect 37369 11033 37381 11036
rect 37415 11033 37427 11067
rect 37369 11027 37427 11033
rect 2222 10956 2228 11008
rect 2280 10996 2286 11008
rect 8202 10996 8208 11008
rect 2280 10968 8208 10996
rect 2280 10956 2286 10968
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 24762 10996 24768 11008
rect 16724 10968 24768 10996
rect 16724 10956 16730 10968
rect 24762 10956 24768 10968
rect 24820 10956 24826 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 23106 10588 23112 10600
rect 14884 10560 23112 10588
rect 14884 10548 14890 10560
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 17218 10480 17224 10532
rect 17276 10520 17282 10532
rect 37734 10520 37740 10532
rect 17276 10492 37740 10520
rect 17276 10480 17282 10492
rect 37734 10480 37740 10492
rect 37792 10480 37798 10532
rect 37918 10520 37924 10532
rect 37879 10492 37924 10520
rect 37918 10480 37924 10492
rect 37976 10480 37982 10532
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 20070 10452 20076 10464
rect 9456 10424 20076 10452
rect 9456 10412 9462 10424
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 23198 10412 23204 10464
rect 23256 10452 23262 10464
rect 38013 10455 38071 10461
rect 38013 10452 38025 10455
rect 23256 10424 38025 10452
rect 23256 10412 23262 10424
rect 38013 10421 38025 10424
rect 38059 10421 38071 10455
rect 38013 10415 38071 10421
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 37182 10112 37188 10124
rect 37143 10084 37188 10112
rect 37182 10072 37188 10084
rect 37240 10072 37246 10124
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 16206 9908 16212 9920
rect 1627 9880 16212 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 37277 9911 37335 9917
rect 37277 9908 37289 9911
rect 25004 9880 37289 9908
rect 25004 9868 25010 9880
rect 37277 9877 37289 9880
rect 37323 9877 37335 9911
rect 37277 9871 37335 9877
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 22922 9664 22928 9716
rect 22980 9704 22986 9716
rect 26694 9704 26700 9716
rect 22980 9676 26700 9704
rect 22980 9664 22986 9676
rect 26694 9664 26700 9676
rect 26752 9664 26758 9716
rect 18230 9596 18236 9648
rect 18288 9636 18294 9648
rect 23290 9636 23296 9648
rect 18288 9608 23296 9636
rect 18288 9596 18294 9608
rect 23290 9596 23296 9608
rect 23348 9596 23354 9648
rect 37369 9639 37427 9645
rect 37369 9605 37381 9639
rect 37415 9636 37427 9639
rect 37550 9636 37556 9648
rect 37415 9608 37556 9636
rect 37415 9605 37427 9608
rect 37369 9599 37427 9605
rect 37550 9596 37556 9608
rect 37608 9596 37614 9648
rect 37826 9596 37832 9648
rect 37884 9636 37890 9648
rect 38105 9639 38163 9645
rect 38105 9636 38117 9639
rect 37884 9608 38117 9636
rect 37884 9596 37890 9608
rect 38105 9605 38117 9608
rect 38151 9605 38163 9639
rect 38105 9599 38163 9605
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 23106 9568 23112 9580
rect 17000 9540 23112 9568
rect 17000 9528 17006 9540
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 37182 9500 37188 9512
rect 37143 9472 37188 9500
rect 37182 9460 37188 9472
rect 37240 9460 37246 9512
rect 37918 9432 37924 9444
rect 37879 9404 37924 9432
rect 37918 9392 37924 9404
rect 37976 9392 37982 9444
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 13262 9364 13268 9376
rect 1627 9336 13268 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 17678 9324 17684 9376
rect 17736 9364 17742 9376
rect 26878 9364 26884 9376
rect 17736 9336 26884 9364
rect 17736 9324 17742 9336
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 15838 9120 15844 9172
rect 15896 9160 15902 9172
rect 25866 9160 25872 9172
rect 15896 9132 22094 9160
rect 15896 9120 15902 9132
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 21542 8956 21548 8968
rect 6972 8928 21548 8956
rect 6972 8916 6978 8928
rect 21542 8916 21548 8928
rect 21600 8916 21606 8968
rect 22066 8956 22094 9132
rect 22664 9132 25872 9160
rect 22664 9033 22692 9132
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 31202 9120 31208 9172
rect 31260 9160 31266 9172
rect 37277 9163 37335 9169
rect 37277 9160 37289 9163
rect 31260 9132 37289 9160
rect 31260 9120 31266 9132
rect 37277 9129 37289 9132
rect 37323 9129 37335 9163
rect 37277 9123 37335 9129
rect 23382 9092 23388 9104
rect 23343 9064 23388 9092
rect 23382 9052 23388 9064
rect 23440 9052 23446 9104
rect 26878 9052 26884 9104
rect 26936 9092 26942 9104
rect 37550 9092 37556 9104
rect 26936 9064 37556 9092
rect 26936 9052 26942 9064
rect 37550 9052 37556 9064
rect 37608 9052 37614 9104
rect 22649 9027 22707 9033
rect 22649 8993 22661 9027
rect 22695 8993 22707 9027
rect 22830 9024 22836 9036
rect 22791 8996 22836 9024
rect 22649 8987 22707 8993
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 23014 9024 23020 9036
rect 22975 8996 23020 9024
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 23293 9027 23351 9033
rect 23293 8993 23305 9027
rect 23339 9024 23351 9027
rect 25590 9024 25596 9036
rect 23339 8996 25596 9024
rect 23339 8993 23351 8996
rect 23293 8987 23351 8993
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 37182 9024 37188 9036
rect 37143 8996 37188 9024
rect 37182 8984 37188 8996
rect 37240 8984 37246 9036
rect 37826 8956 37832 8968
rect 22066 8928 37832 8956
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 19150 8412 19156 8424
rect 10836 8384 19156 8412
rect 10836 8372 10842 8384
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 24762 8372 24768 8424
rect 24820 8412 24826 8424
rect 38105 8415 38163 8421
rect 38105 8412 38117 8415
rect 24820 8384 38117 8412
rect 24820 8372 24826 8384
rect 38105 8381 38117 8384
rect 38151 8381 38163 8415
rect 38105 8375 38163 8381
rect 13446 8344 13452 8356
rect 1596 8316 13452 8344
rect 1596 8285 1624 8316
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 37918 8344 37924 8356
rect 37879 8316 37924 8344
rect 37918 8304 37924 8316
rect 37976 8304 37982 8356
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8245 1639 8279
rect 1581 8239 1639 8245
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2038 8072 2044 8084
rect 1627 8044 2044 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 6270 8072 6276 8084
rect 2372 8044 6276 8072
rect 2372 8032 2378 8044
rect 6270 8032 6276 8044
rect 6328 8032 6334 8084
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 37182 7936 37188 7948
rect 37143 7908 37188 7936
rect 37182 7896 37188 7908
rect 37240 7896 37246 7948
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 12342 7868 12348 7880
rect 1636 7840 12348 7868
rect 1636 7828 1642 7840
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 23934 7868 23940 7880
rect 15068 7840 23940 7868
rect 15068 7828 15074 7840
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 23198 7800 23204 7812
rect 11020 7772 23204 7800
rect 11020 7760 11026 7772
rect 23198 7760 23204 7772
rect 23256 7760 23262 7812
rect 24854 7760 24860 7812
rect 24912 7800 24918 7812
rect 36446 7800 36452 7812
rect 24912 7772 36452 7800
rect 24912 7760 24918 7772
rect 36446 7760 36452 7772
rect 36504 7760 36510 7812
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 37277 7735 37335 7741
rect 37277 7732 37289 7735
rect 17460 7704 37289 7732
rect 17460 7692 17466 7704
rect 37277 7701 37289 7704
rect 37323 7701 37335 7735
rect 37277 7695 37335 7701
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 20622 7528 20628 7540
rect 17175 7500 20628 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22462 7488 22468 7540
rect 22520 7528 22526 7540
rect 26602 7528 26608 7540
rect 22520 7500 26608 7528
rect 22520 7488 22526 7500
rect 26602 7488 26608 7500
rect 26660 7488 26666 7540
rect 37642 7488 37648 7540
rect 37700 7528 37706 7540
rect 38013 7531 38071 7537
rect 38013 7528 38025 7531
rect 37700 7500 38025 7528
rect 37700 7488 37706 7500
rect 38013 7497 38025 7500
rect 38059 7497 38071 7531
rect 38013 7491 38071 7497
rect 16850 7324 16856 7336
rect 16811 7296 16856 7324
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 37182 7324 37188 7336
rect 37143 7296 37188 7324
rect 37182 7284 37188 7296
rect 37240 7284 37246 7336
rect 37918 7256 37924 7268
rect 37879 7228 37924 7256
rect 37918 7216 37924 7228
rect 37976 7216 37982 7268
rect 23290 7148 23296 7200
rect 23348 7188 23354 7200
rect 37277 7191 37335 7197
rect 37277 7188 37289 7191
rect 23348 7160 37289 7188
rect 23348 7148 23354 7160
rect 37277 7157 37289 7160
rect 37323 7157 37335 7191
rect 37277 7151 37335 7157
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 20070 6944 20076 6996
rect 20128 6984 20134 6996
rect 26510 6984 26516 6996
rect 20128 6956 26516 6984
rect 20128 6944 20134 6956
rect 26510 6944 26516 6956
rect 26568 6944 26574 6996
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 17310 6848 17316 6860
rect 13136 6820 17316 6848
rect 13136 6808 13142 6820
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 35250 6808 35256 6860
rect 35308 6848 35314 6860
rect 36538 6848 36544 6860
rect 35308 6820 36544 6848
rect 35308 6808 35314 6820
rect 36538 6808 36544 6820
rect 36596 6808 36602 6860
rect 37182 6848 37188 6860
rect 37143 6820 37188 6848
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 37274 6808 37280 6860
rect 37332 6848 37338 6860
rect 37369 6851 37427 6857
rect 37369 6848 37381 6851
rect 37332 6820 37381 6848
rect 37332 6808 37338 6820
rect 37369 6817 37381 6820
rect 37415 6817 37427 6851
rect 37369 6811 37427 6817
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 21266 6780 21272 6792
rect 15252 6752 21272 6780
rect 15252 6740 15258 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 1762 6712 1768 6724
rect 1627 6684 1768 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 1670 6440 1676 6452
rect 1627 6412 1676 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 37090 6400 37096 6452
rect 37148 6440 37154 6452
rect 37277 6443 37335 6449
rect 37277 6440 37289 6443
rect 37148 6412 37289 6440
rect 37148 6400 37154 6412
rect 37277 6409 37289 6412
rect 37323 6409 37335 6443
rect 37277 6403 37335 6409
rect 18874 6332 18880 6384
rect 18932 6372 18938 6384
rect 27338 6372 27344 6384
rect 18932 6344 27344 6372
rect 18932 6332 18938 6344
rect 27338 6332 27344 6344
rect 27396 6332 27402 6384
rect 36906 6332 36912 6384
rect 36964 6372 36970 6384
rect 38105 6375 38163 6381
rect 38105 6372 38117 6375
rect 36964 6344 38117 6372
rect 36964 6332 36970 6344
rect 38105 6341 38117 6344
rect 38151 6341 38163 6375
rect 38105 6335 38163 6341
rect 2498 6264 2504 6316
rect 2556 6304 2562 6316
rect 14458 6304 14464 6316
rect 2556 6276 14464 6304
rect 2556 6264 2562 6276
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 22278 6304 22284 6316
rect 14976 6276 22284 6304
rect 14976 6264 14982 6276
rect 22278 6264 22284 6276
rect 22336 6264 22342 6316
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20404 6208 22094 6236
rect 20404 6196 20410 6208
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 20162 6168 20168 6180
rect 5132 6140 20168 6168
rect 5132 6128 5138 6140
rect 20162 6128 20168 6140
rect 20220 6128 20226 6180
rect 22066 6100 22094 6208
rect 36354 6128 36360 6180
rect 36412 6168 36418 6180
rect 36449 6171 36507 6177
rect 36449 6168 36461 6171
rect 36412 6140 36461 6168
rect 36412 6128 36418 6140
rect 36449 6137 36461 6140
rect 36495 6137 36507 6171
rect 36449 6131 36507 6137
rect 36633 6171 36691 6177
rect 36633 6137 36645 6171
rect 36679 6168 36691 6171
rect 36998 6168 37004 6180
rect 36679 6140 37004 6168
rect 36679 6137 36691 6140
rect 36633 6131 36691 6137
rect 36998 6128 37004 6140
rect 37056 6128 37062 6180
rect 37090 6128 37096 6180
rect 37148 6168 37154 6180
rect 37185 6171 37243 6177
rect 37185 6168 37197 6171
rect 37148 6140 37197 6168
rect 37148 6128 37154 6140
rect 37185 6137 37197 6140
rect 37231 6137 37243 6171
rect 37918 6168 37924 6180
rect 37879 6140 37924 6168
rect 37185 6131 37243 6137
rect 37918 6128 37924 6140
rect 37976 6128 37982 6180
rect 37274 6100 37280 6112
rect 22066 6072 37280 6100
rect 37274 6060 37280 6072
rect 37332 6060 37338 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 3510 5896 3516 5908
rect 1627 5868 3516 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 28350 5788 28356 5840
rect 28408 5828 28414 5840
rect 35345 5831 35403 5837
rect 35345 5828 35357 5831
rect 28408 5800 35357 5828
rect 28408 5788 28414 5800
rect 35345 5797 35357 5800
rect 35391 5797 35403 5831
rect 35345 5791 35403 5797
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 2130 5720 2136 5772
rect 2188 5760 2194 5772
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2188 5732 2881 5760
rect 2188 5720 2194 5732
rect 2869 5729 2881 5732
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 30558 5720 30564 5772
rect 30616 5760 30622 5772
rect 36081 5763 36139 5769
rect 36081 5760 36093 5763
rect 30616 5732 36093 5760
rect 30616 5720 30622 5732
rect 36081 5729 36093 5732
rect 36127 5729 36139 5763
rect 37182 5760 37188 5772
rect 37143 5732 37188 5760
rect 36081 5723 36139 5729
rect 37182 5720 37188 5732
rect 37240 5720 37246 5772
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5534 5692 5540 5704
rect 5040 5664 5540 5692
rect 5040 5652 5046 5664
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 23106 5584 23112 5636
rect 23164 5624 23170 5636
rect 37369 5627 37427 5633
rect 37369 5624 37381 5627
rect 23164 5596 37381 5624
rect 23164 5584 23170 5596
rect 37369 5593 37381 5596
rect 37415 5593 37427 5627
rect 37369 5587 37427 5593
rect 2685 5559 2743 5565
rect 2685 5525 2697 5559
rect 2731 5556 2743 5559
rect 4890 5556 4896 5568
rect 2731 5528 4896 5556
rect 2731 5525 2743 5528
rect 2685 5519 2743 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 13354 5516 13360 5568
rect 13412 5556 13418 5568
rect 15746 5556 15752 5568
rect 13412 5528 15752 5556
rect 13412 5516 13418 5528
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 17402 5516 17408 5568
rect 17460 5556 17466 5568
rect 24210 5556 24216 5568
rect 17460 5528 24216 5556
rect 17460 5516 17466 5528
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 35437 5559 35495 5565
rect 35437 5525 35449 5559
rect 35483 5556 35495 5559
rect 35618 5556 35624 5568
rect 35483 5528 35624 5556
rect 35483 5525 35495 5528
rect 35437 5519 35495 5525
rect 35618 5516 35624 5528
rect 35676 5516 35682 5568
rect 36078 5516 36084 5568
rect 36136 5556 36142 5568
rect 36173 5559 36231 5565
rect 36173 5556 36185 5559
rect 36136 5528 36185 5556
rect 36136 5516 36142 5528
rect 36173 5525 36185 5528
rect 36219 5525 36231 5559
rect 36173 5519 36231 5525
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 6362 5352 6368 5364
rect 3007 5324 6368 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 28902 5312 28908 5364
rect 28960 5352 28966 5364
rect 29546 5352 29552 5364
rect 28960 5324 29552 5352
rect 28960 5312 28966 5324
rect 29546 5312 29552 5324
rect 29604 5312 29610 5364
rect 36538 5352 36544 5364
rect 36499 5324 36544 5352
rect 36538 5312 36544 5324
rect 36596 5312 36602 5364
rect 37734 5312 37740 5364
rect 37792 5352 37798 5364
rect 38013 5355 38071 5361
rect 38013 5352 38025 5355
rect 37792 5324 38025 5352
rect 37792 5312 37798 5324
rect 38013 5321 38025 5324
rect 38059 5321 38071 5355
rect 38013 5315 38071 5321
rect 37366 5284 37372 5296
rect 37327 5256 37372 5284
rect 37366 5244 37372 5256
rect 37424 5244 37430 5296
rect 34606 5176 34612 5228
rect 34664 5216 34670 5228
rect 35526 5216 35532 5228
rect 34664 5188 35532 5216
rect 34664 5176 34670 5188
rect 35526 5176 35532 5188
rect 35584 5176 35590 5228
rect 1302 5108 1308 5160
rect 1360 5148 1366 5160
rect 1397 5151 1455 5157
rect 1397 5148 1409 5151
rect 1360 5120 1409 5148
rect 1360 5108 1366 5120
rect 1397 5117 1409 5120
rect 1443 5117 1455 5151
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 1397 5111 1455 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 31294 5108 31300 5160
rect 31352 5148 31358 5160
rect 31481 5151 31539 5157
rect 31481 5148 31493 5151
rect 31352 5120 31493 5148
rect 31352 5108 31358 5120
rect 31481 5117 31493 5120
rect 31527 5117 31539 5151
rect 31481 5111 31539 5117
rect 34057 5151 34115 5157
rect 34057 5117 34069 5151
rect 34103 5148 34115 5151
rect 36906 5148 36912 5160
rect 34103 5120 36912 5148
rect 34103 5117 34115 5120
rect 34057 5111 34115 5117
rect 36906 5108 36912 5120
rect 36964 5108 36970 5160
rect 37182 5148 37188 5160
rect 37143 5120 37188 5148
rect 37182 5108 37188 5120
rect 37240 5108 37246 5160
rect 6178 5040 6184 5092
rect 6236 5080 6242 5092
rect 12434 5080 12440 5092
rect 6236 5052 12440 5080
rect 6236 5040 6242 5052
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 31754 5040 31760 5092
rect 31812 5080 31818 5092
rect 33873 5083 33931 5089
rect 33873 5080 33885 5083
rect 31812 5052 33885 5080
rect 31812 5040 31818 5052
rect 33873 5049 33885 5052
rect 33919 5049 33931 5083
rect 34606 5080 34612 5092
rect 34567 5052 34612 5080
rect 33873 5043 33931 5049
rect 34606 5040 34612 5052
rect 34664 5040 34670 5092
rect 36449 5083 36507 5089
rect 36449 5049 36461 5083
rect 36495 5080 36507 5083
rect 36630 5080 36636 5092
rect 36495 5052 36636 5080
rect 36495 5049 36507 5052
rect 36449 5043 36507 5049
rect 36630 5040 36636 5052
rect 36688 5040 36694 5092
rect 37918 5080 37924 5092
rect 37879 5052 37924 5080
rect 37918 5040 37924 5052
rect 37976 5040 37982 5092
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 22186 5012 22192 5024
rect 11756 4984 22192 5012
rect 11756 4972 11762 4984
rect 22186 4972 22192 4984
rect 22244 4972 22250 5024
rect 31297 5015 31355 5021
rect 31297 4981 31309 5015
rect 31343 5012 31355 5015
rect 33594 5012 33600 5024
rect 31343 4984 33600 5012
rect 31343 4981 31355 4984
rect 31297 4975 31355 4981
rect 33594 4972 33600 4984
rect 33652 4972 33658 5024
rect 34701 5015 34759 5021
rect 34701 4981 34713 5015
rect 34747 5012 34759 5015
rect 38930 5012 38936 5024
rect 34747 4984 38936 5012
rect 34747 4981 34759 4984
rect 34701 4975 34759 4981
rect 38930 4972 38936 4984
rect 38988 4972 38994 5024
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 20898 4808 20904 4820
rect 9640 4780 20904 4808
rect 9640 4768 9646 4780
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 36262 4768 36268 4820
rect 36320 4808 36326 4820
rect 36541 4811 36599 4817
rect 36541 4808 36553 4811
rect 36320 4780 36553 4808
rect 36320 4768 36326 4780
rect 36541 4777 36553 4780
rect 36587 4777 36599 4811
rect 36541 4771 36599 4777
rect 25958 4700 25964 4752
rect 26016 4740 26022 4752
rect 34241 4743 34299 4749
rect 34241 4740 34253 4743
rect 26016 4712 34253 4740
rect 26016 4700 26022 4712
rect 34241 4709 34253 4712
rect 34287 4709 34299 4743
rect 34241 4703 34299 4709
rect 34514 4700 34520 4752
rect 34572 4740 34578 4752
rect 34977 4743 35035 4749
rect 34977 4740 34989 4743
rect 34572 4712 34989 4740
rect 34572 4700 34578 4712
rect 34977 4709 34989 4712
rect 35023 4709 35035 4743
rect 34977 4703 35035 4709
rect 35897 4743 35955 4749
rect 35897 4709 35909 4743
rect 35943 4740 35955 4743
rect 36170 4740 36176 4752
rect 35943 4712 36176 4740
rect 35943 4709 35955 4712
rect 35897 4703 35955 4709
rect 36170 4700 36176 4712
rect 36228 4700 36234 4752
rect 37369 4743 37427 4749
rect 37369 4709 37381 4743
rect 37415 4740 37427 4743
rect 37458 4740 37464 4752
rect 37415 4712 37464 4740
rect 37415 4709 37427 4712
rect 37369 4703 37427 4709
rect 37458 4700 37464 4712
rect 37516 4700 37522 4752
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 3329 4675 3387 4681
rect 3329 4672 3341 4675
rect 1903 4644 3341 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 3329 4641 3341 4644
rect 3375 4641 3387 4675
rect 14642 4672 14648 4684
rect 14603 4644 14648 4672
rect 3329 4635 3387 4641
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 22278 4632 22284 4684
rect 22336 4672 22342 4684
rect 22741 4675 22799 4681
rect 22741 4672 22753 4675
rect 22336 4644 22753 4672
rect 22336 4632 22342 4644
rect 22741 4641 22753 4644
rect 22787 4641 22799 4675
rect 23385 4675 23443 4681
rect 23385 4672 23397 4675
rect 22741 4635 22799 4641
rect 22848 4644 23397 4672
rect 22646 4564 22652 4616
rect 22704 4604 22710 4616
rect 22848 4604 22876 4644
rect 23385 4641 23397 4644
rect 23431 4641 23443 4675
rect 23385 4635 23443 4641
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25409 4675 25467 4681
rect 25409 4672 25421 4675
rect 25188 4644 25421 4672
rect 25188 4632 25194 4644
rect 25409 4641 25421 4644
rect 25455 4641 25467 4675
rect 25409 4635 25467 4641
rect 26602 4632 26608 4684
rect 26660 4672 26666 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 26660 4644 26801 4672
rect 26660 4632 26666 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 30190 4632 30196 4684
rect 30248 4672 30254 4684
rect 30285 4675 30343 4681
rect 30285 4672 30297 4675
rect 30248 4644 30297 4672
rect 30248 4632 30254 4644
rect 30285 4641 30297 4644
rect 30331 4641 30343 4675
rect 30285 4635 30343 4641
rect 30745 4675 30803 4681
rect 30745 4641 30757 4675
rect 30791 4641 30803 4675
rect 30745 4635 30803 4641
rect 30760 4604 30788 4635
rect 31018 4632 31024 4684
rect 31076 4672 31082 4684
rect 31573 4675 31631 4681
rect 31573 4672 31585 4675
rect 31076 4644 31585 4672
rect 31076 4632 31082 4644
rect 31573 4641 31585 4644
rect 31619 4641 31631 4675
rect 31573 4635 31631 4641
rect 33226 4632 33232 4684
rect 33284 4672 33290 4684
rect 33505 4675 33563 4681
rect 33505 4672 33517 4675
rect 33284 4644 33517 4672
rect 33284 4632 33290 4644
rect 33505 4641 33517 4644
rect 33551 4641 33563 4675
rect 33505 4635 33563 4641
rect 35713 4675 35771 4681
rect 35713 4641 35725 4675
rect 35759 4672 35771 4675
rect 35802 4672 35808 4684
rect 35759 4644 35808 4672
rect 35759 4641 35771 4644
rect 35713 4635 35771 4641
rect 35802 4632 35808 4644
rect 35860 4632 35866 4684
rect 36449 4675 36507 4681
rect 36449 4641 36461 4675
rect 36495 4672 36507 4675
rect 36538 4672 36544 4684
rect 36495 4644 36544 4672
rect 36495 4641 36507 4644
rect 36449 4635 36507 4641
rect 36538 4632 36544 4644
rect 36596 4632 36602 4684
rect 37182 4672 37188 4684
rect 37143 4644 37188 4672
rect 37182 4632 37188 4644
rect 37240 4632 37246 4684
rect 22704 4576 22876 4604
rect 23216 4576 30788 4604
rect 33689 4607 33747 4613
rect 22704 4564 22710 4576
rect 23216 4545 23244 4576
rect 33689 4573 33701 4607
rect 33735 4604 33747 4607
rect 36262 4604 36268 4616
rect 33735 4576 36268 4604
rect 33735 4573 33747 4576
rect 33689 4567 33747 4573
rect 36262 4564 36268 4576
rect 36320 4564 36326 4616
rect 23201 4539 23259 4545
rect 23201 4505 23213 4539
rect 23247 4505 23259 4539
rect 23201 4499 23259 4505
rect 30929 4539 30987 4545
rect 30929 4505 30941 4539
rect 30975 4536 30987 4539
rect 33318 4536 33324 4548
rect 30975 4508 33324 4536
rect 30975 4505 30987 4508
rect 30929 4499 30987 4505
rect 33318 4496 33324 4508
rect 33376 4496 33382 4548
rect 34425 4539 34483 4545
rect 34425 4505 34437 4539
rect 34471 4536 34483 4539
rect 34471 4508 35894 4536
rect 34471 4505 34483 4508
rect 34425 4499 34483 4505
rect 1118 4428 1124 4480
rect 1176 4468 1182 4480
rect 1949 4471 2007 4477
rect 1949 4468 1961 4471
rect 1176 4440 1961 4468
rect 1176 4428 1182 4440
rect 1949 4437 1961 4440
rect 1995 4437 2007 4471
rect 1949 4431 2007 4437
rect 2038 4428 2044 4480
rect 2096 4468 2102 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 2096 4440 2697 4468
rect 2096 4428 2102 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 2685 4431 2743 4437
rect 2958 4428 2964 4480
rect 3016 4468 3022 4480
rect 8938 4468 8944 4480
rect 3016 4440 8944 4468
rect 3016 4428 3022 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 20714 4468 20720 4480
rect 14875 4440 20720 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 20714 4428 20720 4440
rect 20772 4428 20778 4480
rect 22554 4468 22560 4480
rect 22515 4440 22560 4468
rect 22554 4428 22560 4440
rect 22612 4428 22618 4480
rect 25222 4468 25228 4480
rect 25183 4440 25228 4468
rect 25222 4428 25228 4440
rect 25280 4428 25286 4480
rect 26234 4428 26240 4480
rect 26292 4468 26298 4480
rect 26605 4471 26663 4477
rect 26605 4468 26617 4471
rect 26292 4440 26617 4468
rect 26292 4428 26298 4440
rect 26605 4437 26617 4440
rect 26651 4437 26663 4471
rect 26605 4431 26663 4437
rect 29730 4428 29736 4480
rect 29788 4468 29794 4480
rect 30101 4471 30159 4477
rect 30101 4468 30113 4471
rect 29788 4440 30113 4468
rect 29788 4428 29794 4440
rect 30101 4437 30113 4440
rect 30147 4437 30159 4471
rect 31386 4468 31392 4480
rect 31347 4440 31392 4468
rect 30101 4431 30159 4437
rect 31386 4428 31392 4440
rect 31444 4428 31450 4480
rect 35069 4471 35127 4477
rect 35069 4437 35081 4471
rect 35115 4468 35127 4471
rect 35434 4468 35440 4480
rect 35115 4440 35440 4468
rect 35115 4437 35127 4440
rect 35069 4431 35127 4437
rect 35434 4428 35440 4440
rect 35492 4428 35498 4480
rect 35866 4468 35894 4508
rect 36170 4468 36176 4480
rect 35866 4440 36176 4468
rect 36170 4428 36176 4440
rect 36228 4428 36234 4480
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 10229 4267 10287 4273
rect 10229 4264 10241 4267
rect 6886 4236 10241 4264
rect 4249 4199 4307 4205
rect 4249 4165 4261 4199
rect 4295 4165 4307 4199
rect 4249 4159 4307 4165
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 4264 4128 4292 4159
rect 6886 4128 6914 4236
rect 10229 4233 10241 4236
rect 10275 4233 10287 4267
rect 10229 4227 10287 4233
rect 21174 4224 21180 4276
rect 21232 4264 21238 4276
rect 22370 4264 22376 4276
rect 21232 4236 22376 4264
rect 21232 4224 21238 4236
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 25222 4224 25228 4276
rect 25280 4264 25286 4276
rect 32490 4264 32496 4276
rect 25280 4236 32496 4264
rect 25280 4224 25286 4236
rect 32490 4224 32496 4236
rect 32548 4224 32554 4276
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 23934 4196 23940 4208
rect 20772 4168 22784 4196
rect 23895 4168 23940 4196
rect 20772 4156 20778 4168
rect 2004 4100 2728 4128
rect 4264 4100 6914 4128
rect 9861 4131 9919 4137
rect 2004 4088 2010 4100
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2038 4060 2044 4072
rect 1903 4032 2044 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2038 4020 2044 4032
rect 2096 4020 2102 4072
rect 2590 4060 2596 4072
rect 2551 4032 2596 4060
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 2700 4060 2728 4100
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 14734 4128 14740 4140
rect 9907 4100 14740 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 22756 4128 22784 4168
rect 23934 4156 23940 4168
rect 23992 4156 23998 4208
rect 26789 4199 26847 4205
rect 26789 4165 26801 4199
rect 26835 4165 26847 4199
rect 28534 4196 28540 4208
rect 26789 4159 26847 4165
rect 28184 4168 28396 4196
rect 28495 4168 28540 4196
rect 26804 4128 26832 4159
rect 28184 4128 28212 4168
rect 14936 4100 22692 4128
rect 22756 4100 26648 4128
rect 26804 4100 28212 4128
rect 28368 4128 28396 4168
rect 28534 4156 28540 4168
rect 28592 4156 28598 4208
rect 33042 4156 33048 4208
rect 33100 4196 33106 4208
rect 33100 4168 34008 4196
rect 33100 4156 33106 4168
rect 30282 4128 30288 4140
rect 28368 4100 30288 4128
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 2700 4032 4445 4060
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 4433 4023 4491 4029
rect 4540 4032 4905 4060
rect 1486 3952 1492 4004
rect 1544 3992 1550 4004
rect 2777 3995 2835 4001
rect 2777 3992 2789 3995
rect 1544 3964 2789 3992
rect 1544 3952 1550 3964
rect 2777 3961 2789 3964
rect 2823 3961 2835 3995
rect 2777 3955 2835 3961
rect 3602 3952 3608 4004
rect 3660 3992 3666 4004
rect 4540 3992 4568 4032
rect 4893 4029 4905 4032
rect 4939 4029 4951 4063
rect 4893 4023 4951 4029
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 3660 3964 4568 3992
rect 3660 3952 3666 3964
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5552 3992 5580 4023
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5960 4032 6193 4060
rect 5960 4020 5966 4032
rect 6181 4029 6193 4032
rect 6227 4029 6239 4063
rect 7098 4060 7104 4072
rect 7059 4032 7104 4060
rect 6181 4023 6239 4029
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 10962 4060 10968 4072
rect 10923 4032 10968 4060
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 4856 3964 5580 3992
rect 4856 3952 4862 3964
rect 8938 3952 8944 4004
rect 8996 3992 9002 4004
rect 8996 3964 11928 3992
rect 8996 3952 9002 3964
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 1949 3927 2007 3933
rect 1949 3924 1961 3927
rect 992 3896 1961 3924
rect 992 3884 998 3896
rect 1949 3893 1961 3896
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 4948 3896 10241 3924
rect 4948 3884 4954 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10229 3887 10287 3893
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10652 3896 11069 3924
rect 10652 3884 10658 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11480 3896 11805 3924
rect 11480 3884 11486 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11900 3924 11928 3964
rect 14936 3924 14964 4100
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15930 4060 15936 4072
rect 15068 4032 15113 4060
rect 15891 4032 15936 4060
rect 15068 4020 15074 4032
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 17862 4020 17868 4072
rect 17920 4060 17926 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17920 4032 18061 4060
rect 17920 4020 17926 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20165 4063 20223 4069
rect 20165 4060 20177 4063
rect 19484 4032 20177 4060
rect 19484 4020 19490 4032
rect 20165 4029 20177 4032
rect 20211 4029 20223 4063
rect 20165 4023 20223 4029
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20809 4063 20867 4069
rect 20809 4060 20821 4063
rect 20588 4032 20821 4060
rect 20588 4020 20594 4032
rect 20809 4029 20821 4032
rect 20855 4029 20867 4063
rect 20809 4023 20867 4029
rect 21358 4020 21364 4072
rect 21416 4060 21422 4072
rect 22664 4069 22692 4100
rect 21545 4063 21603 4069
rect 21545 4060 21557 4063
rect 21416 4032 21557 4060
rect 21416 4020 21422 4032
rect 21545 4029 21557 4032
rect 21591 4029 21603 4063
rect 21545 4023 21603 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4029 22063 4063
rect 22005 4023 22063 4029
rect 22649 4063 22707 4069
rect 22649 4029 22661 4063
rect 22695 4029 22707 4063
rect 23290 4060 23296 4072
rect 23251 4032 23296 4060
rect 22649 4023 22707 4029
rect 15378 3952 15384 4004
rect 15436 3992 15442 4004
rect 22020 3992 22048 4023
rect 23290 4020 23296 4032
rect 23348 4020 23354 4072
rect 24121 4063 24179 4069
rect 24121 4029 24133 4063
rect 24167 4029 24179 4063
rect 24121 4023 24179 4029
rect 15436 3964 22048 3992
rect 15436 3952 15442 3964
rect 23106 3952 23112 4004
rect 23164 3992 23170 4004
rect 24136 3992 24164 4023
rect 24854 4020 24860 4072
rect 24912 4060 24918 4072
rect 25409 4063 25467 4069
rect 25409 4060 25421 4063
rect 24912 4032 25421 4060
rect 24912 4020 24918 4032
rect 25409 4029 25421 4032
rect 25455 4029 25467 4063
rect 25409 4023 25467 4029
rect 25774 4020 25780 4072
rect 25832 4060 25838 4072
rect 26620 4069 26648 4100
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 30374 4088 30380 4140
rect 30432 4128 30438 4140
rect 33980 4128 34008 4168
rect 34330 4156 34336 4208
rect 34388 4196 34394 4208
rect 34701 4199 34759 4205
rect 34701 4196 34713 4199
rect 34388 4168 34713 4196
rect 34388 4156 34394 4168
rect 34701 4165 34713 4168
rect 34747 4165 34759 4199
rect 34701 4159 34759 4165
rect 36354 4128 36360 4140
rect 30432 4100 33916 4128
rect 33980 4100 36360 4128
rect 30432 4088 30438 4100
rect 26053 4063 26111 4069
rect 26053 4060 26065 4063
rect 25832 4032 26065 4060
rect 25832 4020 25838 4032
rect 26053 4029 26065 4032
rect 26099 4029 26111 4063
rect 26053 4023 26111 4029
rect 26605 4063 26663 4069
rect 26605 4029 26617 4063
rect 26651 4029 26663 4063
rect 26605 4023 26663 4029
rect 27249 4063 27307 4069
rect 27249 4029 27261 4063
rect 27295 4029 27307 4063
rect 27249 4023 27307 4029
rect 27154 3992 27160 4004
rect 23164 3964 24164 3992
rect 25056 3964 27160 3992
rect 23164 3952 23170 3964
rect 15102 3924 15108 3936
rect 11900 3896 14964 3924
rect 15063 3896 15108 3924
rect 11793 3887 11851 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15896 3896 16037 3924
rect 15896 3884 15902 3896
rect 16025 3893 16037 3896
rect 16071 3893 16083 3927
rect 16025 3887 16083 3893
rect 17586 3884 17592 3936
rect 17644 3924 17650 3936
rect 17865 3927 17923 3933
rect 17865 3924 17877 3927
rect 17644 3896 17877 3924
rect 17644 3884 17650 3896
rect 17865 3893 17877 3896
rect 17911 3893 17923 3927
rect 17865 3887 17923 3893
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 18012 3896 19993 3924
rect 18012 3884 18018 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 20622 3924 20628 3936
rect 20583 3896 20628 3924
rect 19981 3887 20039 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3924 21419 3927
rect 22094 3924 22100 3936
rect 21407 3896 22100 3924
rect 21407 3893 21419 3896
rect 21361 3887 21419 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22833 3927 22891 3933
rect 22244 3896 22289 3924
rect 22244 3884 22250 3896
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 23382 3924 23388 3936
rect 22879 3896 23388 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23477 3927 23535 3933
rect 23477 3893 23489 3927
rect 23523 3924 23535 3927
rect 25056 3924 25084 3964
rect 27154 3952 27160 3964
rect 27212 3952 27218 4004
rect 27264 3992 27292 4023
rect 27430 4020 27436 4072
rect 27488 4060 27494 4072
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 27488 4032 28089 4060
rect 27488 4020 27494 4032
rect 28077 4029 28089 4032
rect 28123 4029 28135 4063
rect 28077 4023 28135 4029
rect 28350 4020 28356 4072
rect 28408 4060 28414 4072
rect 28721 4063 28779 4069
rect 28721 4060 28733 4063
rect 28408 4032 28733 4060
rect 28408 4020 28414 4032
rect 28721 4029 28733 4032
rect 28767 4029 28779 4063
rect 28721 4023 28779 4029
rect 29270 4020 29276 4072
rect 29328 4060 29334 4072
rect 29457 4063 29515 4069
rect 29457 4060 29469 4063
rect 29328 4032 29469 4060
rect 29328 4020 29334 4032
rect 29457 4029 29469 4032
rect 29503 4029 29515 4063
rect 30558 4060 30564 4072
rect 29457 4023 29515 4029
rect 29564 4032 30564 4060
rect 28534 3992 28540 4004
rect 27264 3964 28540 3992
rect 28534 3952 28540 3964
rect 28592 3952 28598 4004
rect 29564 3992 29592 4032
rect 30558 4020 30564 4032
rect 30616 4020 30622 4072
rect 30834 4060 30840 4072
rect 30795 4032 30840 4060
rect 30834 4020 30840 4032
rect 30892 4020 30898 4072
rect 32490 4060 32496 4072
rect 32451 4032 32496 4060
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 33226 4060 33232 4072
rect 32876 4032 33232 4060
rect 28644 3964 29592 3992
rect 25222 3924 25228 3936
rect 23523 3896 25084 3924
rect 25183 3896 25228 3924
rect 23523 3893 23535 3896
rect 23477 3887 23535 3893
rect 25222 3884 25228 3896
rect 25280 3884 25286 3936
rect 25869 3927 25927 3933
rect 25869 3893 25881 3927
rect 25915 3924 25927 3927
rect 26510 3924 26516 3936
rect 25915 3896 26516 3924
rect 25915 3893 25927 3896
rect 25869 3887 25927 3893
rect 26510 3884 26516 3896
rect 26568 3884 26574 3936
rect 27338 3924 27344 3936
rect 27299 3896 27344 3924
rect 27338 3884 27344 3896
rect 27396 3884 27402 3936
rect 27890 3924 27896 3936
rect 27851 3896 27896 3924
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 27982 3884 27988 3936
rect 28040 3924 28046 3936
rect 28644 3924 28672 3964
rect 30466 3952 30472 4004
rect 30524 3992 30530 4004
rect 31665 3995 31723 4001
rect 31665 3992 31677 3995
rect 30524 3964 31677 3992
rect 30524 3952 30530 3964
rect 31665 3961 31677 3964
rect 31711 3961 31723 3995
rect 31665 3955 31723 3961
rect 28040 3896 28672 3924
rect 29273 3927 29331 3933
rect 28040 3884 28046 3896
rect 29273 3893 29285 3927
rect 29319 3924 29331 3927
rect 29546 3924 29552 3936
rect 29319 3896 29552 3924
rect 29319 3893 29331 3896
rect 29273 3887 29331 3893
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 30742 3884 30748 3936
rect 30800 3924 30806 3936
rect 30929 3927 30987 3933
rect 30929 3924 30941 3927
rect 30800 3896 30941 3924
rect 30800 3884 30806 3896
rect 30929 3893 30941 3896
rect 30975 3893 30987 3927
rect 30929 3887 30987 3893
rect 31570 3884 31576 3936
rect 31628 3924 31634 3936
rect 31757 3927 31815 3933
rect 31757 3924 31769 3927
rect 31628 3896 31769 3924
rect 31628 3884 31634 3896
rect 31757 3893 31769 3896
rect 31803 3893 31815 3927
rect 31757 3887 31815 3893
rect 32309 3927 32367 3933
rect 32309 3893 32321 3927
rect 32355 3924 32367 3927
rect 32876 3924 32904 4032
rect 33226 4020 33232 4032
rect 33284 4020 33290 4072
rect 33888 4069 33916 4100
rect 36354 4088 36360 4100
rect 36412 4088 36418 4140
rect 36446 4088 36452 4140
rect 36504 4128 36510 4140
rect 36633 4131 36691 4137
rect 36633 4128 36645 4131
rect 36504 4100 36645 4128
rect 36504 4088 36510 4100
rect 36633 4097 36645 4100
rect 36679 4097 36691 4131
rect 36633 4091 36691 4097
rect 37369 4131 37427 4137
rect 37369 4097 37381 4131
rect 37415 4128 37427 4131
rect 37550 4128 37556 4140
rect 37415 4100 37556 4128
rect 37415 4097 37427 4100
rect 37369 4091 37427 4097
rect 37550 4088 37556 4100
rect 37608 4088 37614 4140
rect 37826 4088 37832 4140
rect 37884 4128 37890 4140
rect 38105 4131 38163 4137
rect 38105 4128 38117 4131
rect 37884 4100 38117 4128
rect 37884 4088 37890 4100
rect 38105 4097 38117 4100
rect 38151 4097 38163 4131
rect 38105 4091 38163 4097
rect 33873 4063 33931 4069
rect 33873 4029 33885 4063
rect 33919 4029 33931 4063
rect 34514 4060 34520 4072
rect 34475 4032 34520 4060
rect 33873 4023 33931 4029
rect 34514 4020 34520 4032
rect 34572 4020 34578 4072
rect 35897 4063 35955 4069
rect 35897 4029 35909 4063
rect 35943 4029 35955 4063
rect 35897 4023 35955 4029
rect 33137 3995 33195 4001
rect 33137 3961 33149 3995
rect 33183 3992 33195 3995
rect 33318 3992 33324 4004
rect 33183 3964 33324 3992
rect 33183 3961 33195 3964
rect 33137 3955 33195 3961
rect 33318 3952 33324 3964
rect 33376 3952 33382 4004
rect 33594 3952 33600 4004
rect 33652 3992 33658 4004
rect 35912 3992 35940 4023
rect 36262 4020 36268 4072
rect 36320 4060 36326 4072
rect 39482 4060 39488 4072
rect 36320 4032 39488 4060
rect 36320 4020 36326 4032
rect 39482 4020 39488 4032
rect 39540 4020 39546 4072
rect 36446 3992 36452 4004
rect 33652 3964 35940 3992
rect 36407 3964 36452 3992
rect 33652 3952 33658 3964
rect 36446 3952 36452 3964
rect 36504 3952 36510 4004
rect 36814 3952 36820 4004
rect 36872 3992 36878 4004
rect 37185 3995 37243 4001
rect 37185 3992 37197 3995
rect 36872 3964 37197 3992
rect 36872 3952 36878 3964
rect 37185 3961 37197 3964
rect 37231 3961 37243 3995
rect 37185 3955 37243 3961
rect 37921 3995 37979 4001
rect 37921 3961 37933 3995
rect 37967 3992 37979 3995
rect 38102 3992 38108 4004
rect 37967 3964 38108 3992
rect 37967 3961 37979 3964
rect 37921 3955 37979 3961
rect 38102 3952 38108 3964
rect 38160 3952 38166 4004
rect 33226 3924 33232 3936
rect 32355 3896 32904 3924
rect 33187 3896 33232 3924
rect 32355 3893 32367 3896
rect 32309 3887 32367 3893
rect 33226 3884 33232 3896
rect 33284 3884 33290 3936
rect 33965 3927 34023 3933
rect 33965 3893 33977 3927
rect 34011 3924 34023 3927
rect 34606 3924 34612 3936
rect 34011 3896 34612 3924
rect 34011 3893 34023 3896
rect 33965 3887 34023 3893
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 35713 3927 35771 3933
rect 35713 3924 35725 3927
rect 35400 3896 35725 3924
rect 35400 3884 35406 3896
rect 35713 3893 35725 3896
rect 35759 3893 35771 3927
rect 35713 3887 35771 3893
rect 36906 3884 36912 3936
rect 36964 3924 36970 3936
rect 37458 3924 37464 3936
rect 36964 3896 37464 3924
rect 36964 3884 36970 3896
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2314 3720 2320 3732
rect 1995 3692 2320 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 3418 3720 3424 3732
rect 2464 3692 3280 3720
rect 3379 3692 3424 3720
rect 2464 3680 2470 3692
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 3050 3652 3056 3664
rect 1903 3624 3056 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3252 3593 3280 3692
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3689 7803 3723
rect 8754 3720 8760 3732
rect 8715 3692 8760 3720
rect 7745 3683 7803 3689
rect 4062 3652 4068 3664
rect 4023 3624 4068 3652
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 6972 3624 7017 3652
rect 6972 3612 6978 3624
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3584 2651 3587
rect 3237 3587 3295 3593
rect 2639 3556 3188 3584
rect 2639 3553 2651 3556
rect 2593 3547 2651 3553
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3516 2835 3519
rect 2958 3516 2964 3528
rect 2823 3488 2964 3516
rect 2823 3485 2835 3488
rect 2777 3479 2835 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3160 3516 3188 3556
rect 3237 3553 3249 3587
rect 3283 3553 3295 3587
rect 4982 3584 4988 3596
rect 4943 3556 4988 3584
rect 3237 3547 3295 3553
rect 4982 3544 4988 3556
rect 5040 3544 5046 3596
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 5408 3556 5641 3584
rect 5408 3544 5414 3556
rect 5629 3553 5641 3556
rect 5675 3553 5687 3587
rect 5629 3547 5687 3553
rect 7374 3544 7380 3596
rect 7432 3584 7438 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7432 3556 7573 3584
rect 7432 3544 7438 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 3326 3516 3332 3528
rect 3160 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 7760 3516 7788 3683
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 11054 3720 11060 3732
rect 11015 3692 11060 3720
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 12250 3720 12256 3732
rect 12211 3692 12256 3720
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 16298 3720 16304 3732
rect 16259 3692 16304 3720
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 19978 3720 19984 3732
rect 16408 3692 19984 3720
rect 9398 3652 9404 3664
rect 9359 3624 9404 3652
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3652 10195 3655
rect 10226 3652 10232 3664
rect 10183 3624 10232 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 12894 3652 12900 3664
rect 12855 3624 12900 3652
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 14056 3624 14105 3652
rect 14056 3612 14062 3624
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 14550 3612 14556 3664
rect 14608 3652 14614 3664
rect 16408 3652 16436 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20438 3680 20444 3732
rect 20496 3720 20502 3732
rect 22005 3723 22063 3729
rect 20496 3692 21128 3720
rect 20496 3680 20502 3692
rect 17402 3652 17408 3664
rect 14608 3624 16436 3652
rect 17363 3624 17408 3652
rect 14608 3612 14614 3624
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 18138 3652 18144 3664
rect 18099 3624 18144 3652
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18248 3624 21036 3652
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11054 3584 11060 3596
rect 10919 3556 11060 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 12066 3584 12072 3596
rect 12027 3556 12072 3584
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 13814 3584 13820 3596
rect 13775 3556 13820 3584
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 14826 3584 14832 3596
rect 14787 3556 14832 3584
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 15473 3587 15531 3593
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 16022 3584 16028 3596
rect 15519 3556 16028 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 16117 3587 16175 3593
rect 16117 3553 16129 3587
rect 16163 3584 16175 3587
rect 16390 3584 16396 3596
rect 16163 3556 16396 3584
rect 16163 3553 16175 3556
rect 16117 3547 16175 3553
rect 16390 3544 16396 3556
rect 16448 3544 16454 3596
rect 15378 3516 15384 3528
rect 7760 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 18248 3516 18276 3624
rect 18874 3584 18880 3596
rect 18835 3556 18880 3584
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 21008 3593 21036 3624
rect 19705 3587 19763 3593
rect 19705 3553 19717 3587
rect 19751 3553 19763 3587
rect 19705 3547 19763 3553
rect 20349 3587 20407 3593
rect 20349 3553 20361 3587
rect 20395 3553 20407 3587
rect 20349 3547 20407 3553
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3553 21051 3587
rect 21100 3584 21128 3692
rect 22005 3689 22017 3723
rect 22051 3720 22063 3723
rect 23290 3720 23296 3732
rect 22051 3692 23296 3720
rect 22051 3689 22063 3692
rect 22005 3683 22063 3689
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 26142 3720 26148 3732
rect 23768 3692 26148 3720
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 23768 3652 23796 3692
rect 26142 3680 26148 3692
rect 26200 3680 26206 3732
rect 26237 3723 26295 3729
rect 26237 3689 26249 3723
rect 26283 3720 26295 3723
rect 26786 3720 26792 3732
rect 26283 3692 26792 3720
rect 26283 3689 26295 3692
rect 26237 3683 26295 3689
rect 26786 3680 26792 3692
rect 26844 3680 26850 3732
rect 27157 3723 27215 3729
rect 27157 3689 27169 3723
rect 27203 3720 27215 3723
rect 33502 3720 33508 3732
rect 27203 3692 31340 3720
rect 33463 3692 33508 3720
rect 27203 3689 27215 3692
rect 27157 3683 27215 3689
rect 22244 3624 23796 3652
rect 23845 3655 23903 3661
rect 22244 3612 22250 3624
rect 23845 3621 23857 3655
rect 23891 3652 23903 3655
rect 24302 3652 24308 3664
rect 23891 3624 24308 3652
rect 23891 3621 23903 3624
rect 23845 3615 23903 3621
rect 24302 3612 24308 3624
rect 24360 3612 24366 3664
rect 24394 3612 24400 3664
rect 24452 3652 24458 3664
rect 25406 3652 25412 3664
rect 24452 3624 24808 3652
rect 25367 3624 25412 3652
rect 24452 3612 24458 3624
rect 22922 3584 22928 3596
rect 21100 3556 22784 3584
rect 22883 3556 22928 3584
rect 20993 3547 21051 3553
rect 15580 3488 18276 3516
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 15580 3448 15608 3488
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19720 3516 19748 3547
rect 18840 3488 19748 3516
rect 18840 3476 18846 3488
rect 5859 3420 15608 3448
rect 15657 3451 15715 3457
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 16850 3448 16856 3460
rect 15703 3420 16856 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 16942 3408 16948 3460
rect 17000 3448 17006 3460
rect 20364 3448 20392 3547
rect 22186 3516 22192 3528
rect 20548 3488 22192 3516
rect 20548 3457 20576 3488
rect 22186 3476 22192 3488
rect 22244 3476 22250 3528
rect 22756 3516 22784 3556
rect 22922 3544 22928 3556
rect 22980 3544 22986 3596
rect 23750 3584 23756 3596
rect 23032 3556 23756 3584
rect 23032 3516 23060 3556
rect 23750 3544 23756 3556
rect 23808 3544 23814 3596
rect 24026 3544 24032 3596
rect 24084 3584 24090 3596
rect 24673 3587 24731 3593
rect 24673 3584 24685 3587
rect 24084 3556 24685 3584
rect 24084 3544 24090 3556
rect 24673 3553 24685 3556
rect 24719 3553 24731 3587
rect 24780 3584 24808 3624
rect 25406 3612 25412 3624
rect 25464 3612 25470 3664
rect 27982 3652 27988 3664
rect 25516 3624 27988 3652
rect 25516 3584 25544 3624
rect 27982 3612 27988 3624
rect 28040 3612 28046 3664
rect 28169 3655 28227 3661
rect 28169 3621 28181 3655
rect 28215 3652 28227 3655
rect 28258 3652 28264 3664
rect 28215 3624 28264 3652
rect 28215 3621 28227 3624
rect 28169 3615 28227 3621
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 28902 3652 28908 3664
rect 28863 3624 28908 3652
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 30374 3652 30380 3664
rect 29380 3624 30380 3652
rect 26050 3584 26056 3596
rect 24780 3556 25544 3584
rect 26011 3556 26056 3584
rect 24673 3547 24731 3553
rect 26050 3544 26056 3556
rect 26108 3544 26114 3596
rect 26142 3544 26148 3596
rect 26200 3584 26206 3596
rect 29380 3584 29408 3624
rect 30374 3612 30380 3624
rect 30432 3612 30438 3664
rect 30466 3612 30472 3664
rect 30524 3652 30530 3664
rect 30524 3624 30569 3652
rect 30524 3612 30530 3624
rect 30650 3612 30656 3664
rect 30708 3652 30714 3664
rect 31021 3655 31079 3661
rect 31021 3652 31033 3655
rect 30708 3624 31033 3652
rect 30708 3612 30714 3624
rect 31021 3621 31033 3624
rect 31067 3621 31079 3655
rect 31021 3615 31079 3621
rect 29546 3584 29552 3596
rect 26200 3556 29408 3584
rect 29507 3556 29552 3584
rect 26200 3544 26206 3556
rect 29546 3544 29552 3556
rect 29604 3544 29610 3596
rect 29730 3544 29736 3596
rect 29788 3584 29794 3596
rect 30071 3587 30129 3593
rect 30071 3584 30083 3587
rect 29788 3556 30083 3584
rect 29788 3544 29794 3556
rect 30071 3553 30083 3556
rect 30117 3553 30129 3587
rect 30071 3547 30129 3553
rect 30558 3544 30564 3596
rect 30616 3584 30622 3596
rect 31205 3587 31263 3593
rect 31205 3584 31217 3587
rect 30616 3556 31217 3584
rect 30616 3544 30622 3556
rect 31205 3553 31217 3556
rect 31251 3553 31263 3587
rect 31312 3584 31340 3692
rect 33502 3680 33508 3692
rect 33560 3680 33566 3732
rect 34238 3720 34244 3732
rect 34199 3692 34244 3720
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 34790 3680 34796 3732
rect 34848 3720 34854 3732
rect 34977 3723 35035 3729
rect 34977 3720 34989 3723
rect 34848 3692 34989 3720
rect 34848 3680 34854 3692
rect 34977 3689 34989 3692
rect 35023 3689 35035 3723
rect 34977 3683 35035 3689
rect 35894 3680 35900 3732
rect 35952 3720 35958 3732
rect 35952 3692 35997 3720
rect 35952 3680 35958 3692
rect 36722 3680 36728 3732
rect 36780 3720 36786 3732
rect 37277 3723 37335 3729
rect 37277 3720 37289 3723
rect 36780 3692 37289 3720
rect 36780 3680 36786 3692
rect 37277 3689 37289 3692
rect 37323 3689 37335 3723
rect 37277 3683 37335 3689
rect 31478 3612 31484 3664
rect 31536 3652 31542 3664
rect 34330 3652 34336 3664
rect 31536 3624 34336 3652
rect 31536 3612 31542 3624
rect 34330 3612 34336 3624
rect 34388 3612 34394 3664
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 36906 3652 36912 3664
rect 34664 3624 36912 3652
rect 34664 3612 34670 3624
rect 36906 3612 36912 3624
rect 36964 3612 36970 3664
rect 31941 3587 31999 3593
rect 31941 3584 31953 3587
rect 31312 3556 31953 3584
rect 31205 3547 31263 3553
rect 31941 3553 31953 3556
rect 31987 3553 31999 3587
rect 33318 3584 33324 3596
rect 33279 3556 33324 3584
rect 31941 3547 31999 3553
rect 33318 3544 33324 3556
rect 33376 3544 33382 3596
rect 33962 3544 33968 3596
rect 34020 3584 34026 3596
rect 34057 3587 34115 3593
rect 34057 3584 34069 3587
rect 34020 3556 34069 3584
rect 34020 3544 34026 3556
rect 34057 3553 34069 3556
rect 34103 3553 34115 3587
rect 34057 3547 34115 3553
rect 34238 3544 34244 3596
rect 34296 3584 34302 3596
rect 34793 3587 34851 3593
rect 34793 3584 34805 3587
rect 34296 3556 34805 3584
rect 34296 3544 34302 3556
rect 34793 3553 34805 3556
rect 34839 3553 34851 3587
rect 35710 3584 35716 3596
rect 35671 3556 35716 3584
rect 34793 3547 34851 3553
rect 35710 3544 35716 3556
rect 35768 3544 35774 3596
rect 37182 3584 37188 3596
rect 37143 3556 37188 3584
rect 37182 3544 37188 3556
rect 37240 3544 37246 3596
rect 22756 3488 23060 3516
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 33042 3516 33048 3528
rect 23440 3488 33048 3516
rect 23440 3476 23446 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 39206 3516 39212 3528
rect 33284 3488 39212 3516
rect 33284 3476 33290 3488
rect 39206 3476 39212 3488
rect 39264 3476 39270 3528
rect 17000 3420 20392 3448
rect 20533 3451 20591 3457
rect 17000 3408 17006 3420
rect 20533 3417 20545 3451
rect 20579 3417 20591 3451
rect 20533 3411 20591 3417
rect 21177 3451 21235 3457
rect 21177 3417 21189 3451
rect 21223 3448 21235 3451
rect 27157 3451 27215 3457
rect 27157 3448 27169 3451
rect 21223 3420 22600 3448
rect 21223 3417 21235 3420
rect 21177 3411 21235 3417
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 4157 3383 4215 3389
rect 4157 3380 4169 3383
rect 3292 3352 4169 3380
rect 3292 3340 3298 3352
rect 4157 3349 4169 3352
rect 4203 3349 4215 3383
rect 5166 3380 5172 3392
rect 5127 3352 5172 3380
rect 4157 3343 4215 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6880 3352 7021 3380
rect 6880 3340 6886 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 9493 3383 9551 3389
rect 9493 3380 9505 3383
rect 8904 3352 9505 3380
rect 8904 3340 8910 3352
rect 9493 3349 9505 3352
rect 9539 3349 9551 3383
rect 9493 3343 9551 3349
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 9732 3352 10241 3380
rect 9732 3340 9738 3352
rect 10229 3349 10241 3352
rect 10275 3349 10287 3383
rect 10229 3343 10287 3349
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 12989 3383 13047 3389
rect 12989 3380 13001 3383
rect 12400 3352 13001 3380
rect 12400 3340 12406 3352
rect 12989 3349 13001 3352
rect 13035 3349 13047 3383
rect 12989 3343 13047 3349
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14148 3352 14933 3380
rect 14148 3340 14154 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 16724 3352 17509 3380
rect 16724 3340 16730 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 17678 3340 17684 3392
rect 17736 3380 17742 3392
rect 18233 3383 18291 3389
rect 18233 3380 18245 3383
rect 17736 3352 18245 3380
rect 17736 3340 17742 3352
rect 18233 3349 18245 3352
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 18969 3383 19027 3389
rect 18969 3380 18981 3383
rect 18564 3352 18981 3380
rect 18564 3340 18570 3352
rect 18969 3349 18981 3352
rect 19015 3349 19027 3383
rect 19518 3380 19524 3392
rect 19479 3352 19524 3380
rect 18969 3343 19027 3349
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 22005 3383 22063 3389
rect 22005 3380 22017 3383
rect 20036 3352 22017 3380
rect 20036 3340 20042 3352
rect 22005 3349 22017 3352
rect 22051 3349 22063 3383
rect 22572 3380 22600 3420
rect 22756 3420 27169 3448
rect 22756 3380 22784 3420
rect 27157 3417 27169 3420
rect 27203 3417 27215 3451
rect 27157 3411 27215 3417
rect 27338 3408 27344 3460
rect 27396 3448 27402 3460
rect 30009 3451 30067 3457
rect 30009 3448 30021 3451
rect 27396 3420 30021 3448
rect 27396 3408 27402 3420
rect 30009 3417 30021 3420
rect 30055 3417 30067 3451
rect 31386 3448 31392 3460
rect 30009 3411 30067 3417
rect 30116 3420 31392 3448
rect 22572 3352 22784 3380
rect 22005 3343 22063 3349
rect 22830 3340 22836 3392
rect 22888 3380 22894 3392
rect 23017 3383 23075 3389
rect 23017 3380 23029 3383
rect 22888 3352 23029 3380
rect 22888 3340 22894 3352
rect 23017 3349 23029 3352
rect 23063 3349 23075 3383
rect 23017 3343 23075 3349
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 23937 3383 23995 3389
rect 23937 3380 23949 3383
rect 23808 3352 23949 3380
rect 23808 3340 23814 3352
rect 23937 3349 23949 3352
rect 23983 3349 23995 3383
rect 24486 3380 24492 3392
rect 24447 3352 24492 3380
rect 23937 3343 23995 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 25498 3380 25504 3392
rect 25459 3352 25504 3380
rect 25498 3340 25504 3352
rect 25556 3340 25562 3392
rect 25866 3340 25872 3392
rect 25924 3380 25930 3392
rect 26786 3380 26792 3392
rect 25924 3352 26792 3380
rect 25924 3340 25930 3352
rect 26786 3340 26792 3352
rect 26844 3340 26850 3392
rect 28074 3340 28080 3392
rect 28132 3380 28138 3392
rect 28261 3383 28319 3389
rect 28261 3380 28273 3383
rect 28132 3352 28273 3380
rect 28132 3340 28138 3352
rect 28261 3349 28273 3352
rect 28307 3349 28319 3383
rect 28994 3380 29000 3392
rect 28955 3352 29000 3380
rect 28261 3343 28319 3349
rect 28994 3340 29000 3352
rect 29052 3340 29058 3392
rect 29917 3383 29975 3389
rect 29917 3349 29929 3383
rect 29963 3380 29975 3383
rect 30116 3380 30144 3420
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 32125 3451 32183 3457
rect 32125 3417 32137 3451
rect 32171 3448 32183 3451
rect 36262 3448 36268 3460
rect 32171 3420 36268 3448
rect 32171 3417 32183 3420
rect 32125 3411 32183 3417
rect 36262 3408 36268 3420
rect 36320 3408 36326 3460
rect 29963 3352 30144 3380
rect 29963 3349 29975 3352
rect 29917 3343 29975 3349
rect 30282 3340 30288 3392
rect 30340 3380 30346 3392
rect 34422 3380 34428 3392
rect 30340 3352 34428 3380
rect 30340 3340 30346 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 38654 3380 38660 3392
rect 36228 3352 38660 3380
rect 36228 3340 36234 3352
rect 38654 3340 38660 3352
rect 38712 3340 38718 3392
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2498 3176 2504 3188
rect 1995 3148 2504 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4614 3176 4620 3188
rect 4479 3148 4620 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 7834 3176 7840 3188
rect 7795 3148 7840 3176
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3176 8631 3179
rect 8938 3176 8944 3188
rect 8619 3148 8944 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 11146 3176 11152 3188
rect 11103 3148 11152 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 17586 3176 17592 3188
rect 17547 3148 17592 3176
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 18690 3176 18696 3188
rect 18651 3148 18696 3176
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 20990 3176 20996 3188
rect 20951 3148 20996 3176
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 23550 3179 23608 3185
rect 23550 3145 23562 3179
rect 23596 3176 23608 3179
rect 24486 3176 24492 3188
rect 23596 3148 24492 3176
rect 23596 3145 23608 3148
rect 23550 3139 23608 3145
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 26142 3176 26148 3188
rect 24596 3148 26148 3176
rect 658 3068 664 3120
rect 716 3108 722 3120
rect 4246 3108 4252 3120
rect 716 3080 4252 3108
rect 716 3068 722 3080
rect 4246 3068 4252 3080
rect 4304 3068 4310 3120
rect 5166 3068 5172 3120
rect 5224 3108 5230 3120
rect 16942 3108 16948 3120
rect 5224 3080 16948 3108
rect 5224 3068 5230 3080
rect 16942 3068 16948 3080
rect 17000 3068 17006 3120
rect 17478 3111 17536 3117
rect 17478 3077 17490 3111
rect 17524 3108 17536 3111
rect 20622 3108 20628 3120
rect 17524 3080 20628 3108
rect 17524 3077 17536 3080
rect 17478 3071 17536 3077
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 23661 3111 23719 3117
rect 23661 3108 23673 3111
rect 22152 3080 23673 3108
rect 22152 3068 22158 3080
rect 23661 3077 23673 3080
rect 23707 3077 23719 3111
rect 23661 3071 23719 3077
rect 23842 3068 23848 3120
rect 23900 3108 23906 3120
rect 24596 3108 24624 3148
rect 26142 3136 26148 3148
rect 26200 3136 26206 3188
rect 26310 3179 26368 3185
rect 26310 3145 26322 3179
rect 26356 3176 26368 3179
rect 27890 3176 27896 3188
rect 26356 3148 27896 3176
rect 26356 3145 26368 3148
rect 26310 3139 26368 3145
rect 27890 3136 27896 3148
rect 27948 3136 27954 3188
rect 29362 3136 29368 3188
rect 29420 3176 29426 3188
rect 29457 3179 29515 3185
rect 29457 3176 29469 3179
rect 29420 3148 29469 3176
rect 29420 3136 29426 3148
rect 29457 3145 29469 3148
rect 29503 3145 29515 3179
rect 29457 3139 29515 3145
rect 29914 3136 29920 3188
rect 29972 3176 29978 3188
rect 30558 3176 30564 3188
rect 29972 3148 30564 3176
rect 29972 3136 29978 3148
rect 30558 3136 30564 3148
rect 30616 3136 30622 3188
rect 31662 3176 31668 3188
rect 30944 3148 31668 3176
rect 23900 3080 24624 3108
rect 23900 3068 23906 3080
rect 25222 3068 25228 3120
rect 25280 3108 25286 3120
rect 26421 3111 26479 3117
rect 26421 3108 26433 3111
rect 25280 3080 26433 3108
rect 25280 3068 25286 3080
rect 26421 3077 26433 3080
rect 26467 3077 26479 3111
rect 26786 3108 26792 3120
rect 26747 3080 26792 3108
rect 26421 3071 26479 3077
rect 26786 3068 26792 3080
rect 26844 3068 26850 3120
rect 27154 3068 27160 3120
rect 27212 3108 27218 3120
rect 30944 3108 30972 3148
rect 31662 3136 31668 3148
rect 31720 3136 31726 3188
rect 32398 3176 32404 3188
rect 32359 3148 32404 3176
rect 32398 3136 32404 3148
rect 32456 3136 32462 3188
rect 33134 3176 33140 3188
rect 33095 3148 33140 3176
rect 33134 3136 33140 3148
rect 33192 3136 33198 3188
rect 33870 3176 33876 3188
rect 33831 3148 33876 3176
rect 33870 3136 33876 3148
rect 33928 3136 33934 3188
rect 37826 3176 37832 3188
rect 33980 3148 37832 3176
rect 27212 3080 30972 3108
rect 31021 3111 31079 3117
rect 27212 3068 27218 3080
rect 31021 3077 31033 3111
rect 31067 3108 31079 3111
rect 33980 3108 34008 3148
rect 37826 3136 37832 3148
rect 37884 3136 37890 3188
rect 38010 3176 38016 3188
rect 37971 3148 38016 3176
rect 38010 3136 38016 3148
rect 38068 3136 38074 3188
rect 31067 3080 34008 3108
rect 31067 3077 31079 3080
rect 31021 3071 31079 3077
rect 35618 3068 35624 3120
rect 35676 3108 35682 3120
rect 35676 3080 38056 3108
rect 35676 3068 35682 3080
rect 38028 3052 38056 3080
rect 106 3000 112 3052
rect 164 3040 170 3052
rect 1210 3040 1216 3052
rect 164 3012 1216 3040
rect 164 3000 170 3012
rect 1210 3000 1216 3012
rect 1268 3000 1274 3052
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 6730 3040 6736 3052
rect 6691 3012 6736 3040
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13722 3040 13728 3052
rect 13219 3012 13728 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 19518 3040 19524 3052
rect 17727 3012 19524 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 22428 3012 22508 3040
rect 22428 3000 22434 3012
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 2958 2972 2964 2984
rect 2915 2944 2964 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4212 2944 4261 2972
rect 4212 2932 4218 2944
rect 4249 2941 4261 2944
rect 4295 2941 4307 2975
rect 5074 2972 5080 2984
rect 5035 2944 5080 2972
rect 4249 2935 4307 2941
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 5810 2972 5816 2984
rect 5771 2944 5816 2972
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6454 2972 6460 2984
rect 6415 2944 6460 2972
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 7650 2972 7656 2984
rect 7611 2944 7656 2972
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8260 2944 8401 2972
rect 8260 2932 8266 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 9456 2944 10241 2972
rect 9456 2932 9462 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10870 2972 10876 2984
rect 10831 2944 10876 2972
rect 10229 2935 10287 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 11790 2972 11796 2984
rect 11751 2944 11796 2972
rect 11790 2932 11796 2944
rect 11848 2932 11854 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15562 2972 15568 2984
rect 14792 2944 14964 2972
rect 15523 2944 15568 2972
rect 14792 2932 14798 2944
rect 1857 2907 1915 2913
rect 1857 2873 1869 2907
rect 1903 2904 1915 2907
rect 2774 2904 2780 2916
rect 1903 2876 2780 2904
rect 1903 2873 1915 2876
rect 1857 2867 1915 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 7926 2864 7932 2916
rect 7984 2904 7990 2916
rect 9582 2904 9588 2916
rect 7984 2876 8800 2904
rect 9543 2876 9588 2904
rect 7984 2864 7990 2876
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 5169 2839 5227 2845
rect 5169 2836 5181 2839
rect 4672 2808 5181 2836
rect 4672 2796 4678 2808
rect 5169 2805 5181 2808
rect 5215 2805 5227 2839
rect 5169 2799 5227 2805
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5684 2808 5917 2836
rect 5684 2796 5690 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 8772 2836 8800 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 14550 2904 14556 2916
rect 10428 2876 14556 2904
rect 10428 2845 10456 2876
rect 14550 2864 14556 2876
rect 14608 2864 14614 2916
rect 14826 2904 14832 2916
rect 14787 2876 14832 2904
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 14936 2904 14964 2944
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2972 16635 2975
rect 17034 2972 17040 2984
rect 16623 2944 17040 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17313 2975 17371 2981
rect 17313 2941 17325 2975
rect 17359 2972 17371 2975
rect 17954 2972 17960 2984
rect 17359 2944 17960 2972
rect 17359 2941 17371 2944
rect 17313 2935 17371 2941
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18196 2944 18521 2972
rect 18196 2932 18202 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 20070 2972 20076 2984
rect 20031 2944 20076 2972
rect 18509 2935 18567 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20806 2972 20812 2984
rect 20767 2944 20812 2972
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 21637 2975 21695 2981
rect 21637 2941 21649 2975
rect 21683 2972 21695 2975
rect 21818 2972 21824 2984
rect 21683 2944 21824 2972
rect 21683 2941 21695 2944
rect 21637 2935 21695 2941
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 18049 2907 18107 2913
rect 18049 2904 18061 2907
rect 14936 2876 18061 2904
rect 18049 2873 18061 2876
rect 18095 2873 18107 2907
rect 18049 2867 18107 2873
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 22094 2904 22100 2916
rect 20312 2876 22100 2904
rect 20312 2864 20318 2876
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 22370 2904 22376 2916
rect 22331 2876 22376 2904
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 22480 2904 22508 3012
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 22612 3012 23765 3040
rect 22612 3000 22618 3012
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 26510 3040 26516 3052
rect 23753 3003 23811 3009
rect 24044 3012 26372 3040
rect 26471 3012 26516 3040
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2972 23443 2975
rect 23934 2972 23940 2984
rect 23431 2944 23940 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23934 2932 23940 2944
rect 23992 2932 23998 2984
rect 24044 2904 24072 3012
rect 25314 2972 25320 2984
rect 25275 2944 25320 2972
rect 25314 2932 25320 2944
rect 25372 2932 25378 2984
rect 26145 2975 26203 2981
rect 26145 2941 26157 2975
rect 26191 2972 26203 2975
rect 26234 2972 26240 2984
rect 26191 2944 26240 2972
rect 26191 2941 26203 2944
rect 26145 2935 26203 2941
rect 26234 2932 26240 2944
rect 26292 2932 26298 2984
rect 26344 2972 26372 3012
rect 26510 3000 26516 3012
rect 26568 3000 26574 3052
rect 31478 3040 31484 3052
rect 26620 3012 31484 3040
rect 26620 2972 26648 3012
rect 31478 3000 31484 3012
rect 31536 3000 31542 3052
rect 31757 3043 31815 3049
rect 31757 3009 31769 3043
rect 31803 3040 31815 3043
rect 35986 3040 35992 3052
rect 31803 3012 35894 3040
rect 35947 3012 35992 3040
rect 31803 3009 31815 3012
rect 31757 3003 31815 3009
rect 26344 2944 26648 2972
rect 27433 2975 27491 2981
rect 27433 2941 27445 2975
rect 27479 2972 27491 2975
rect 27522 2972 27528 2984
rect 27479 2944 27528 2972
rect 27479 2941 27491 2944
rect 27433 2935 27491 2941
rect 27522 2932 27528 2944
rect 27580 2932 27586 2984
rect 28166 2972 28172 2984
rect 28127 2944 28172 2972
rect 28166 2932 28172 2944
rect 28224 2932 28230 2984
rect 29273 2975 29331 2981
rect 29273 2941 29285 2975
rect 29319 2972 29331 2975
rect 29546 2972 29552 2984
rect 29319 2944 29552 2972
rect 29319 2941 29331 2944
rect 29273 2935 29331 2941
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 30837 2975 30895 2981
rect 30837 2941 30849 2975
rect 30883 2972 30895 2975
rect 32214 2972 32220 2984
rect 30883 2944 31754 2972
rect 32175 2944 32220 2972
rect 30883 2941 30895 2944
rect 30837 2935 30895 2941
rect 22480 2876 24072 2904
rect 26326 2864 26332 2916
rect 26384 2904 26390 2916
rect 27617 2907 27675 2913
rect 27617 2904 27629 2907
rect 26384 2876 27629 2904
rect 26384 2864 26390 2876
rect 27617 2873 27629 2876
rect 27663 2873 27675 2907
rect 30466 2904 30472 2916
rect 27617 2867 27675 2873
rect 27724 2876 30472 2904
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 8772 2808 9689 2836
rect 5905 2799 5963 2805
rect 9677 2805 9689 2808
rect 9723 2805 9735 2839
rect 9677 2799 9735 2805
rect 10413 2839 10471 2845
rect 10413 2805 10425 2839
rect 10459 2805 10471 2839
rect 10413 2799 10471 2805
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 13228 2808 14933 2836
rect 13228 2796 13234 2808
rect 14921 2805 14933 2808
rect 14967 2805 14979 2839
rect 14921 2799 14979 2805
rect 16761 2839 16819 2845
rect 16761 2805 16773 2839
rect 16807 2836 16819 2839
rect 17770 2836 17776 2848
rect 16807 2808 17776 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 19334 2796 19340 2848
rect 19392 2836 19398 2848
rect 20165 2839 20223 2845
rect 20165 2836 20177 2839
rect 19392 2808 20177 2836
rect 19392 2796 19398 2808
rect 20165 2805 20177 2808
rect 20211 2805 20223 2839
rect 20165 2799 20223 2805
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21729 2839 21787 2845
rect 21729 2836 21741 2839
rect 21140 2808 21741 2836
rect 21140 2796 21146 2808
rect 21729 2805 21741 2808
rect 21775 2805 21787 2839
rect 21729 2799 21787 2805
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 22465 2839 22523 2845
rect 22465 2836 22477 2839
rect 22060 2808 22477 2836
rect 22060 2796 22066 2808
rect 22465 2805 22477 2808
rect 22511 2805 22523 2839
rect 22465 2799 22523 2805
rect 22922 2796 22928 2848
rect 22980 2836 22986 2848
rect 24029 2839 24087 2845
rect 24029 2836 24041 2839
rect 22980 2808 24041 2836
rect 22980 2796 22986 2808
rect 24029 2805 24041 2808
rect 24075 2805 24087 2839
rect 24029 2799 24087 2805
rect 24578 2796 24584 2848
rect 24636 2836 24642 2848
rect 25409 2839 25467 2845
rect 25409 2836 25421 2839
rect 24636 2808 25421 2836
rect 24636 2796 24642 2808
rect 25409 2805 25421 2808
rect 25455 2805 25467 2839
rect 25409 2799 25467 2805
rect 25590 2796 25596 2848
rect 25648 2836 25654 2848
rect 27724 2836 27752 2876
rect 30466 2864 30472 2876
rect 30524 2864 30530 2916
rect 31110 2864 31116 2916
rect 31168 2904 31174 2916
rect 31573 2907 31631 2913
rect 31573 2904 31585 2907
rect 31168 2876 31585 2904
rect 31168 2864 31174 2876
rect 31573 2873 31585 2876
rect 31619 2873 31631 2907
rect 31726 2904 31754 2944
rect 32214 2932 32220 2944
rect 32272 2932 32278 2984
rect 32490 2932 32496 2984
rect 32548 2972 32554 2984
rect 32953 2975 33011 2981
rect 32953 2972 32965 2975
rect 32548 2944 32965 2972
rect 32548 2932 32554 2944
rect 32953 2941 32965 2944
rect 32999 2941 33011 2975
rect 32953 2935 33011 2941
rect 33042 2932 33048 2984
rect 33100 2972 33106 2984
rect 33689 2975 33747 2981
rect 33689 2972 33701 2975
rect 33100 2944 33701 2972
rect 33100 2932 33106 2944
rect 33689 2941 33701 2944
rect 33735 2941 33747 2975
rect 34422 2972 34428 2984
rect 34383 2944 34428 2972
rect 33689 2935 33747 2941
rect 34422 2932 34428 2944
rect 34480 2932 34486 2984
rect 35250 2932 35256 2984
rect 35308 2972 35314 2984
rect 35713 2975 35771 2981
rect 35713 2972 35725 2975
rect 35308 2944 35725 2972
rect 35308 2932 35314 2944
rect 35713 2941 35725 2944
rect 35759 2941 35771 2975
rect 35866 2972 35894 3012
rect 35986 3000 35992 3012
rect 36044 3000 36050 3052
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 37369 3043 37427 3049
rect 37369 3040 37381 3043
rect 37332 3012 37381 3040
rect 37332 3000 37338 3012
rect 37369 3009 37381 3012
rect 37415 3009 37427 3043
rect 37369 3003 37427 3009
rect 38010 3000 38016 3052
rect 38068 3000 38074 3052
rect 37734 2972 37740 2984
rect 35866 2944 37740 2972
rect 35713 2935 35771 2941
rect 37734 2932 37740 2944
rect 37792 2932 37798 2984
rect 35342 2904 35348 2916
rect 31726 2876 35348 2904
rect 31573 2867 31631 2873
rect 35342 2864 35348 2876
rect 35400 2864 35406 2916
rect 36722 2864 36728 2916
rect 36780 2904 36786 2916
rect 37185 2907 37243 2913
rect 37185 2904 37197 2907
rect 36780 2876 37197 2904
rect 36780 2864 36786 2876
rect 37185 2873 37197 2876
rect 37231 2873 37243 2907
rect 37918 2904 37924 2916
rect 37879 2876 37924 2904
rect 37185 2867 37243 2873
rect 37918 2864 37924 2876
rect 37976 2864 37982 2916
rect 28258 2836 28264 2848
rect 25648 2808 27752 2836
rect 28219 2808 28264 2836
rect 25648 2796 25654 2808
rect 28258 2796 28264 2808
rect 28316 2796 28322 2848
rect 28442 2796 28448 2848
rect 28500 2836 28506 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 28500 2808 34621 2836
rect 28500 2796 28506 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 37826 2796 37832 2848
rect 37884 2836 37890 2848
rect 39758 2836 39764 2848
rect 37884 2808 39764 2836
rect 37884 2796 37890 2808
rect 39758 2796 39764 2808
rect 39816 2796 39822 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 4304 2604 5365 2632
rect 4304 2592 4310 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 8573 2635 8631 2641
rect 5592 2604 7696 2632
rect 5592 2592 5598 2604
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 2961 2567 3019 2573
rect 2961 2564 2973 2567
rect 2924 2536 2973 2564
rect 2924 2524 2930 2536
rect 2961 2533 2973 2536
rect 3007 2533 3019 2567
rect 2961 2527 3019 2533
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 4706 2564 4712 2576
rect 4571 2536 4712 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5258 2564 5264 2576
rect 5219 2536 5264 2564
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 7190 2564 7196 2576
rect 7151 2536 7196 2564
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 382 2456 388 2508
rect 440 2496 446 2508
rect 1489 2499 1547 2505
rect 1489 2496 1501 2499
rect 440 2468 1501 2496
rect 440 2456 446 2468
rect 1489 2465 1501 2468
rect 1535 2465 1547 2499
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 1489 2459 1547 2465
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 3936 2468 4261 2496
rect 3936 2456 3942 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6236 2468 6929 2496
rect 6236 2456 6242 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 7668 2428 7696 2604
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 8662 2632 8668 2644
rect 8619 2604 8668 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2632 20499 2635
rect 20990 2632 20996 2644
rect 20487 2604 20996 2632
rect 20487 2601 20499 2604
rect 20441 2595 20499 2601
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 24581 2635 24639 2641
rect 24581 2632 24593 2635
rect 22152 2604 24593 2632
rect 22152 2592 22158 2604
rect 24581 2601 24593 2604
rect 24627 2601 24639 2635
rect 24581 2595 24639 2601
rect 29365 2635 29423 2641
rect 29365 2601 29377 2635
rect 29411 2632 29423 2635
rect 29822 2632 29828 2644
rect 29411 2604 29828 2632
rect 29411 2601 29423 2604
rect 29365 2595 29423 2601
rect 29822 2592 29828 2604
rect 29880 2592 29886 2644
rect 32122 2632 32128 2644
rect 32083 2604 32128 2632
rect 32122 2592 32128 2604
rect 32180 2592 32186 2644
rect 33778 2632 33784 2644
rect 33739 2604 33784 2632
rect 33778 2592 33784 2604
rect 33836 2592 33842 2644
rect 35526 2592 35532 2644
rect 35584 2632 35590 2644
rect 37921 2635 37979 2641
rect 37921 2632 37933 2635
rect 35584 2604 37933 2632
rect 35584 2592 35590 2604
rect 37921 2601 37933 2604
rect 37967 2601 37979 2635
rect 37921 2595 37979 2601
rect 10134 2524 10140 2576
rect 10192 2564 10198 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 10192 2536 10241 2564
rect 10192 2524 10198 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 12434 2524 12440 2576
rect 12492 2564 12498 2576
rect 12897 2567 12955 2573
rect 12897 2564 12909 2567
rect 12492 2536 12909 2564
rect 12492 2524 12498 2536
rect 12897 2533 12909 2536
rect 12943 2533 12955 2567
rect 12897 2527 12955 2533
rect 13817 2567 13875 2573
rect 13817 2533 13829 2567
rect 13863 2564 13875 2567
rect 13906 2564 13912 2576
rect 13863 2536 13912 2564
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 15197 2567 15255 2573
rect 15197 2533 15209 2567
rect 15243 2564 15255 2567
rect 15286 2564 15292 2576
rect 15243 2536 15292 2564
rect 15243 2533 15255 2536
rect 15197 2527 15255 2533
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 17126 2564 17132 2576
rect 16163 2536 17132 2564
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 17865 2567 17923 2573
rect 17865 2564 17877 2567
rect 17460 2536 17877 2564
rect 17460 2524 17466 2536
rect 17865 2533 17877 2536
rect 17911 2533 17923 2567
rect 17865 2527 17923 2533
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 19153 2567 19211 2573
rect 19153 2564 19165 2567
rect 19116 2536 19165 2564
rect 19116 2524 19122 2536
rect 19153 2533 19165 2536
rect 19199 2533 19211 2567
rect 19153 2527 19211 2533
rect 23658 2524 23664 2576
rect 23716 2564 23722 2576
rect 23753 2567 23811 2573
rect 23753 2564 23765 2567
rect 23716 2536 23765 2564
rect 23716 2524 23722 2536
rect 23753 2533 23765 2536
rect 23799 2533 23811 2567
rect 23753 2527 23811 2533
rect 24489 2567 24547 2573
rect 24489 2533 24501 2567
rect 24535 2564 24547 2567
rect 25682 2564 25688 2576
rect 24535 2536 25688 2564
rect 24535 2533 24547 2536
rect 24489 2527 24547 2533
rect 25682 2524 25688 2536
rect 25740 2524 25746 2576
rect 27341 2567 27399 2573
rect 27341 2533 27353 2567
rect 27387 2564 27399 2567
rect 32674 2564 32680 2576
rect 27387 2536 32680 2564
rect 27387 2533 27399 2536
rect 27341 2527 27399 2533
rect 32674 2524 32680 2536
rect 32732 2524 32738 2576
rect 34698 2524 34704 2576
rect 34756 2564 34762 2576
rect 35069 2567 35127 2573
rect 35069 2564 35081 2567
rect 34756 2536 35081 2564
rect 34756 2524 34762 2536
rect 35069 2533 35081 2536
rect 35115 2533 35127 2567
rect 35069 2527 35127 2533
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 9122 2496 9128 2508
rect 8435 2468 9128 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 9950 2496 9956 2508
rect 9911 2468 9956 2496
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10318 2456 10324 2508
rect 10376 2496 10382 2508
rect 10873 2499 10931 2505
rect 10873 2496 10885 2499
rect 10376 2468 10885 2496
rect 10376 2456 10382 2468
rect 10873 2465 10885 2468
rect 10919 2465 10931 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 10873 2459 10931 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13538 2496 13544 2508
rect 13499 2468 13544 2496
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 14921 2459 14979 2465
rect 15304 2468 15853 2496
rect 15304 2440 15332 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17368 2468 17601 2496
rect 17368 2456 17374 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2496 18935 2499
rect 18923 2468 19104 2496
rect 18923 2465 18935 2468
rect 18877 2459 18935 2465
rect 19076 2440 19104 2468
rect 19886 2456 19892 2508
rect 19944 2496 19950 2508
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 19944 2468 20269 2496
rect 19944 2456 19950 2468
rect 20257 2465 20269 2468
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2496 21603 2499
rect 21634 2496 21640 2508
rect 21591 2468 21640 2496
rect 21591 2465 21603 2468
rect 21545 2459 21603 2465
rect 21634 2456 21640 2468
rect 21692 2456 21698 2508
rect 23474 2496 23480 2508
rect 23435 2468 23480 2496
rect 23474 2456 23480 2468
rect 23532 2456 23538 2508
rect 24302 2456 24308 2508
rect 24360 2496 24366 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 24360 2468 25605 2496
rect 24360 2456 24366 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 26970 2496 26976 2508
rect 26931 2468 26976 2496
rect 25593 2459 25651 2465
rect 26970 2456 26976 2468
rect 27028 2456 27034 2508
rect 27798 2456 27804 2508
rect 27856 2496 27862 2508
rect 28353 2499 28411 2505
rect 28353 2496 28365 2499
rect 27856 2468 28365 2496
rect 27856 2456 27862 2468
rect 28353 2465 28365 2468
rect 28399 2465 28411 2499
rect 28353 2459 28411 2465
rect 28718 2456 28724 2508
rect 28776 2496 28782 2508
rect 29181 2499 29239 2505
rect 29181 2496 29193 2499
rect 28776 2468 29193 2496
rect 28776 2456 28782 2468
rect 29181 2465 29193 2468
rect 29227 2465 29239 2499
rect 29181 2459 29239 2465
rect 30466 2456 30472 2508
rect 30524 2496 30530 2508
rect 31021 2499 31079 2505
rect 31021 2496 31033 2499
rect 30524 2468 31033 2496
rect 30524 2456 30530 2468
rect 31021 2465 31033 2468
rect 31067 2465 31079 2499
rect 31938 2496 31944 2508
rect 31899 2468 31944 2496
rect 31021 2459 31079 2465
rect 31938 2456 31944 2468
rect 31996 2456 32002 2508
rect 32766 2456 32772 2508
rect 32824 2496 32830 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 32824 2468 33609 2496
rect 32824 2456 32830 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 34790 2496 34796 2508
rect 34751 2468 34796 2496
rect 33597 2459 33655 2465
rect 34790 2456 34796 2468
rect 34848 2456 34854 2508
rect 36538 2496 36544 2508
rect 36499 2468 36544 2496
rect 36538 2456 36544 2468
rect 36596 2456 36602 2508
rect 37737 2499 37795 2505
rect 37737 2465 37749 2499
rect 37783 2496 37795 2499
rect 38286 2496 38292 2508
rect 37783 2468 38292 2496
rect 37783 2465 37795 2468
rect 37737 2459 37795 2465
rect 38286 2456 38292 2468
rect 38344 2456 38350 2508
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 7668 2400 11069 2428
rect 2041 2391 2099 2397
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 2056 2360 2084 2391
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 19058 2388 19064 2440
rect 19116 2388 19122 2440
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 21729 2431 21787 2437
rect 21729 2428 21741 2431
rect 19208 2400 21741 2428
rect 19208 2388 19214 2400
rect 21729 2397 21741 2400
rect 21775 2397 21787 2431
rect 21729 2391 21787 2397
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2428 25927 2431
rect 28534 2428 28540 2440
rect 25915 2400 28540 2428
rect 25915 2397 25927 2400
rect 25869 2391 25927 2397
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 28629 2431 28687 2437
rect 28629 2397 28641 2431
rect 28675 2428 28687 2431
rect 29638 2428 29644 2440
rect 28675 2400 29644 2428
rect 28675 2397 28687 2400
rect 28629 2391 28687 2397
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 32582 2388 32588 2440
rect 32640 2428 32646 2440
rect 36725 2431 36783 2437
rect 36725 2428 36737 2431
rect 32640 2400 36737 2428
rect 32640 2388 32646 2400
rect 36725 2397 36737 2400
rect 36771 2397 36783 2431
rect 36725 2391 36783 2397
rect 7834 2360 7840 2372
rect 2056 2332 7840 2360
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 21266 2320 21272 2372
rect 21324 2360 21330 2372
rect 31205 2363 31263 2369
rect 31205 2360 31217 2363
rect 21324 2332 31217 2360
rect 21324 2320 21330 2332
rect 31205 2329 31217 2332
rect 31251 2329 31263 2363
rect 31205 2323 31263 2329
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 27246 1436 27252 1488
rect 27304 1476 27310 1488
rect 28258 1476 28264 1488
rect 27304 1448 28264 1476
rect 27304 1436 27310 1448
rect 28258 1436 28264 1448
rect 28316 1436 28322 1488
<< via1 >>
rect 25504 117920 25556 117972
rect 31116 117920 31168 117972
rect 35256 117920 35308 117972
rect 24860 117716 24912 117768
rect 29828 117716 29880 117768
rect 4344 117648 4396 117700
rect 4896 117648 4948 117700
rect 20352 117648 20404 117700
rect 24676 117648 24728 117700
rect 35256 117648 35308 117700
rect 18512 117580 18564 117632
rect 19064 117580 19116 117632
rect 21640 117580 21692 117632
rect 27252 117580 27304 117632
rect 4246 117478 4298 117530
rect 4310 117478 4362 117530
rect 4374 117478 4426 117530
rect 4438 117478 4490 117530
rect 34966 117478 35018 117530
rect 35030 117478 35082 117530
rect 35094 117478 35146 117530
rect 35158 117478 35210 117530
rect 296 117376 348 117428
rect 16580 117376 16632 117428
rect 1124 117308 1176 117360
rect 112 117240 164 117292
rect 664 117172 716 117224
rect 12808 117308 12860 117360
rect 8300 117240 8352 117292
rect 8944 117240 8996 117292
rect 10232 117240 10284 117292
rect 11520 117240 11572 117292
rect 14004 117308 14056 117360
rect 15384 117308 15436 117360
rect 19800 117376 19852 117428
rect 20260 117376 20312 117428
rect 20996 117376 21048 117428
rect 19064 117308 19116 117360
rect 19892 117308 19944 117360
rect 22376 117376 22428 117428
rect 27252 117419 27304 117428
rect 27252 117385 27261 117419
rect 27261 117385 27295 117419
rect 27295 117385 27304 117419
rect 27252 117376 27304 117385
rect 29828 117376 29880 117428
rect 31116 117419 31168 117428
rect 31116 117385 31125 117419
rect 31125 117385 31159 117419
rect 31159 117385 31168 117419
rect 31116 117376 31168 117385
rect 34152 117376 34204 117428
rect 22928 117308 22980 117360
rect 34336 117240 34388 117292
rect 36268 117240 36320 117292
rect 36544 117283 36596 117292
rect 36544 117249 36553 117283
rect 36553 117249 36587 117283
rect 36587 117249 36596 117283
rect 36544 117240 36596 117249
rect 1860 117147 1912 117156
rect 1860 117113 1869 117147
rect 1869 117113 1903 117147
rect 1903 117113 1912 117147
rect 1860 117104 1912 117113
rect 3608 117104 3660 117156
rect 940 117036 992 117088
rect 7840 117215 7892 117224
rect 7840 117181 7849 117215
rect 7849 117181 7883 117215
rect 7883 117181 7892 117215
rect 7840 117172 7892 117181
rect 9588 117172 9640 117224
rect 10876 117172 10928 117224
rect 5080 117147 5132 117156
rect 5080 117113 5089 117147
rect 5089 117113 5123 117147
rect 5123 117113 5132 117147
rect 5080 117104 5132 117113
rect 6736 117104 6788 117156
rect 8116 117104 8168 117156
rect 8392 117147 8444 117156
rect 8392 117113 8401 117147
rect 8401 117113 8435 117147
rect 8435 117113 8444 117147
rect 8392 117104 8444 117113
rect 9496 117104 9548 117156
rect 9772 117104 9824 117156
rect 11152 117147 11204 117156
rect 11152 117113 11161 117147
rect 11161 117113 11195 117147
rect 11195 117113 11204 117147
rect 11152 117104 11204 117113
rect 11336 117104 11388 117156
rect 13084 117147 13136 117156
rect 13084 117113 13093 117147
rect 13093 117113 13127 117147
rect 13127 117113 13136 117147
rect 13084 117104 13136 117113
rect 5264 117036 5316 117088
rect 5908 117036 5960 117088
rect 12164 117036 12216 117088
rect 14096 117172 14148 117224
rect 15844 117172 15896 117224
rect 17776 117172 17828 117224
rect 19340 117172 19392 117224
rect 20444 117172 20496 117224
rect 21640 117172 21692 117224
rect 13820 117147 13872 117156
rect 13820 117113 13829 117147
rect 13829 117113 13863 117147
rect 13863 117113 13872 117147
rect 13820 117104 13872 117113
rect 15016 117147 15068 117156
rect 15016 117113 15025 117147
rect 15025 117113 15059 117147
rect 15059 117113 15068 117147
rect 15016 117104 15068 117113
rect 15936 117104 15988 117156
rect 16580 117104 16632 117156
rect 19064 117104 19116 117156
rect 13452 117036 13504 117088
rect 16304 117036 16356 117088
rect 17868 117036 17920 117088
rect 19892 117104 19944 117156
rect 20536 117104 20588 117156
rect 21364 117104 21416 117156
rect 22008 117172 22060 117224
rect 23204 117147 23256 117156
rect 21732 117036 21784 117088
rect 23204 117113 23213 117147
rect 23213 117113 23247 117147
rect 23247 117113 23256 117147
rect 23204 117104 23256 117113
rect 23296 117104 23348 117156
rect 26700 117172 26752 117224
rect 24124 117104 24176 117156
rect 24768 117104 24820 117156
rect 27160 117147 27212 117156
rect 27160 117113 27169 117147
rect 27169 117113 27203 117147
rect 27203 117113 27212 117147
rect 27160 117104 27212 117113
rect 28356 117147 28408 117156
rect 28356 117113 28365 117147
rect 28365 117113 28399 117147
rect 28399 117113 28408 117147
rect 28356 117104 28408 117113
rect 23940 117036 23992 117088
rect 24676 117036 24728 117088
rect 25964 117036 26016 117088
rect 30656 117104 30708 117156
rect 31760 117147 31812 117156
rect 31760 117113 31769 117147
rect 31769 117113 31803 117147
rect 31803 117113 31812 117147
rect 31760 117104 31812 117113
rect 32312 117104 32364 117156
rect 34244 117147 34296 117156
rect 34244 117113 34253 117147
rect 34253 117113 34287 117147
rect 34287 117113 34296 117147
rect 34244 117104 34296 117113
rect 29184 117079 29236 117088
rect 29184 117045 29193 117079
rect 29193 117045 29227 117079
rect 29227 117045 29236 117079
rect 34980 117172 35032 117224
rect 35624 117104 35676 117156
rect 37096 117172 37148 117224
rect 37740 117172 37792 117224
rect 37924 117147 37976 117156
rect 29184 117036 29236 117045
rect 36452 117036 36504 117088
rect 37924 117113 37933 117147
rect 37933 117113 37967 117147
rect 37967 117113 37976 117147
rect 37924 117104 37976 117113
rect 39028 117036 39080 117088
rect 19606 116934 19658 116986
rect 19670 116934 19722 116986
rect 19734 116934 19786 116986
rect 19798 116934 19850 116986
rect 1308 116832 1360 116884
rect 2596 116832 2648 116884
rect 6460 116832 6512 116884
rect 7104 116832 7156 116884
rect 8576 116832 8628 116884
rect 9312 116832 9364 116884
rect 11704 116832 11756 116884
rect 12440 116832 12492 116884
rect 13636 116832 13688 116884
rect 14740 116832 14792 116884
rect 16764 116832 16816 116884
rect 17592 116832 17644 116884
rect 18696 116832 18748 116884
rect 20444 116875 20496 116884
rect 20444 116841 20453 116875
rect 20453 116841 20487 116875
rect 20487 116841 20496 116875
rect 20444 116832 20496 116841
rect 20720 116832 20772 116884
rect 22284 116832 22336 116884
rect 2136 116764 2188 116816
rect 3240 116764 3292 116816
rect 7840 116764 7892 116816
rect 9680 116764 9732 116816
rect 13176 116764 13228 116816
rect 14280 116764 14332 116816
rect 16028 116764 16080 116816
rect 17868 116764 17920 116816
rect 18052 116764 18104 116816
rect 19156 116764 19208 116816
rect 22376 116764 22428 116816
rect 22652 116807 22704 116816
rect 22652 116773 22678 116807
rect 22678 116773 22704 116807
rect 22652 116764 22704 116773
rect 2596 116739 2648 116748
rect 2596 116705 2605 116739
rect 2605 116705 2639 116739
rect 2639 116705 2648 116739
rect 2596 116696 2648 116705
rect 3792 116696 3844 116748
rect 4068 116739 4120 116748
rect 4068 116705 4077 116739
rect 4077 116705 4111 116739
rect 4111 116705 4120 116739
rect 4068 116696 4120 116705
rect 4804 116739 4856 116748
rect 4804 116705 4813 116739
rect 4813 116705 4847 116739
rect 4847 116705 4856 116739
rect 4804 116696 4856 116705
rect 5540 116739 5592 116748
rect 5540 116705 5549 116739
rect 5549 116705 5583 116739
rect 5583 116705 5592 116739
rect 5540 116696 5592 116705
rect 6920 116739 6972 116748
rect 6920 116705 6929 116739
rect 6929 116705 6963 116739
rect 6963 116705 6972 116739
rect 6920 116696 6972 116705
rect 7012 116696 7064 116748
rect 8576 116696 8628 116748
rect 9864 116739 9916 116748
rect 9864 116705 9873 116739
rect 9873 116705 9907 116739
rect 9907 116705 9916 116739
rect 9864 116696 9916 116705
rect 10600 116739 10652 116748
rect 10600 116705 10609 116739
rect 10609 116705 10643 116739
rect 10643 116705 10652 116739
rect 10600 116696 10652 116705
rect 12164 116739 12216 116748
rect 12164 116705 12173 116739
rect 12173 116705 12207 116739
rect 12207 116705 12216 116739
rect 12164 116696 12216 116705
rect 12900 116739 12952 116748
rect 12900 116705 12909 116739
rect 12909 116705 12943 116739
rect 12943 116705 12952 116739
rect 12900 116696 12952 116705
rect 12992 116696 13044 116748
rect 14372 116739 14424 116748
rect 14372 116705 14381 116739
rect 14381 116705 14415 116739
rect 14415 116705 14424 116739
rect 14372 116696 14424 116705
rect 15108 116739 15160 116748
rect 15108 116705 15117 116739
rect 15117 116705 15151 116739
rect 15151 116705 15160 116739
rect 15108 116696 15160 116705
rect 15568 116696 15620 116748
rect 17408 116739 17460 116748
rect 17408 116705 17417 116739
rect 17417 116705 17451 116739
rect 17451 116705 17460 116739
rect 17408 116696 17460 116705
rect 18144 116739 18196 116748
rect 18144 116705 18153 116739
rect 18153 116705 18187 116739
rect 18187 116705 18196 116739
rect 18144 116696 18196 116705
rect 18880 116739 18932 116748
rect 18880 116705 18889 116739
rect 18889 116705 18923 116739
rect 18923 116705 18932 116739
rect 18880 116696 18932 116705
rect 19340 116696 19392 116748
rect 20352 116739 20404 116748
rect 20352 116705 20361 116739
rect 20361 116705 20395 116739
rect 20395 116705 20404 116739
rect 20352 116696 20404 116705
rect 23664 116832 23716 116884
rect 24216 116832 24268 116884
rect 24492 116832 24544 116884
rect 25688 116832 25740 116884
rect 26792 116832 26844 116884
rect 29092 116832 29144 116884
rect 30012 116832 30064 116884
rect 26056 116764 26108 116816
rect 26148 116764 26200 116816
rect 28540 116764 28592 116816
rect 34612 116832 34664 116884
rect 34888 116832 34940 116884
rect 31024 116764 31076 116816
rect 33048 116764 33100 116816
rect 34980 116764 35032 116816
rect 35348 116764 35400 116816
rect 24308 116739 24360 116748
rect 24308 116705 24317 116739
rect 24317 116705 24351 116739
rect 24351 116705 24360 116739
rect 24308 116696 24360 116705
rect 25596 116696 25648 116748
rect 25780 116739 25832 116748
rect 25780 116705 25789 116739
rect 25789 116705 25823 116739
rect 25823 116705 25832 116739
rect 25780 116696 25832 116705
rect 26516 116739 26568 116748
rect 26516 116705 26525 116739
rect 26525 116705 26559 116739
rect 26559 116705 26568 116739
rect 26516 116696 26568 116705
rect 3884 116628 3936 116680
rect 14648 116628 14700 116680
rect 16304 116628 16356 116680
rect 17224 116628 17276 116680
rect 19064 116628 19116 116680
rect 20076 116628 20128 116680
rect 22008 116628 22060 116680
rect 22100 116628 22152 116680
rect 6552 116560 6604 116612
rect 17960 116560 18012 116612
rect 21732 116560 21784 116612
rect 21824 116560 21876 116612
rect 30196 116696 30248 116748
rect 31668 116696 31720 116748
rect 32772 116696 32824 116748
rect 34704 116739 34756 116748
rect 29644 116671 29696 116680
rect 29644 116637 29653 116671
rect 29653 116637 29687 116671
rect 29687 116637 29696 116671
rect 29644 116628 29696 116637
rect 31024 116628 31076 116680
rect 33416 116628 33468 116680
rect 34704 116705 34713 116739
rect 34713 116705 34747 116739
rect 34747 116705 34756 116739
rect 34704 116696 34756 116705
rect 34612 116628 34664 116680
rect 35900 116696 35952 116748
rect 35532 116628 35584 116680
rect 28816 116560 28868 116612
rect 38844 116560 38896 116612
rect 3424 116535 3476 116544
rect 3424 116501 3433 116535
rect 3433 116501 3467 116535
rect 3467 116501 3476 116535
rect 3424 116492 3476 116501
rect 7656 116492 7708 116544
rect 21088 116492 21140 116544
rect 22376 116492 22428 116544
rect 22468 116492 22520 116544
rect 25044 116492 25096 116544
rect 29368 116492 29420 116544
rect 29552 116535 29604 116544
rect 29552 116501 29561 116535
rect 29561 116501 29595 116535
rect 29595 116501 29604 116535
rect 29552 116492 29604 116501
rect 30932 116492 30984 116544
rect 31208 116535 31260 116544
rect 31208 116501 31217 116535
rect 31217 116501 31251 116535
rect 31251 116501 31260 116535
rect 31208 116492 31260 116501
rect 33140 116492 33192 116544
rect 33600 116492 33652 116544
rect 35440 116492 35492 116544
rect 4246 116390 4298 116442
rect 4310 116390 4362 116442
rect 4374 116390 4426 116442
rect 4438 116390 4490 116442
rect 34966 116390 35018 116442
rect 35030 116390 35082 116442
rect 35094 116390 35146 116442
rect 35158 116390 35210 116442
rect 2228 116288 2280 116340
rect 2780 116288 2832 116340
rect 4620 116288 4672 116340
rect 5816 116288 5868 116340
rect 6644 116288 6696 116340
rect 10416 116288 10468 116340
rect 11060 116288 11112 116340
rect 15660 116288 15712 116340
rect 19984 116288 20036 116340
rect 21272 116288 21324 116340
rect 22100 116288 22152 116340
rect 22652 116288 22704 116340
rect 22928 116288 22980 116340
rect 23112 116288 23164 116340
rect 23756 116288 23808 116340
rect 25872 116288 25924 116340
rect 26608 116288 26660 116340
rect 28172 116288 28224 116340
rect 35256 116288 35308 116340
rect 1860 116220 1912 116272
rect 3608 116152 3660 116204
rect 4528 116152 4580 116204
rect 5172 116220 5224 116272
rect 6000 116220 6052 116272
rect 16120 116220 16172 116272
rect 9496 116195 9548 116204
rect 9496 116161 9505 116195
rect 9505 116161 9539 116195
rect 9539 116161 9548 116195
rect 9496 116152 9548 116161
rect 13084 116152 13136 116204
rect 15016 116152 15068 116204
rect 19892 116152 19944 116204
rect 5172 116084 5224 116136
rect 13820 116084 13872 116136
rect 15936 116084 15988 116136
rect 21364 116220 21416 116272
rect 22376 116220 22428 116272
rect 24768 116220 24820 116272
rect 26700 116220 26752 116272
rect 26976 116220 27028 116272
rect 30748 116263 30800 116272
rect 30748 116229 30757 116263
rect 30757 116229 30791 116263
rect 30791 116229 30800 116263
rect 30748 116220 30800 116229
rect 23112 116152 23164 116204
rect 26240 116152 26292 116204
rect 2320 116059 2372 116068
rect 2320 116025 2329 116059
rect 2329 116025 2363 116059
rect 2363 116025 2372 116059
rect 2320 116016 2372 116025
rect 3056 116059 3108 116068
rect 3056 116025 3065 116059
rect 3065 116025 3099 116059
rect 3099 116025 3108 116059
rect 3056 116016 3108 116025
rect 5448 116016 5500 116068
rect 5724 116016 5776 116068
rect 6276 116059 6328 116068
rect 6276 116025 6285 116059
rect 6285 116025 6319 116059
rect 6319 116025 6328 116059
rect 6276 116016 6328 116025
rect 7564 116016 7616 116068
rect 7748 116059 7800 116068
rect 7748 116025 7757 116059
rect 7757 116025 7791 116059
rect 7791 116025 7800 116059
rect 7748 116016 7800 116025
rect 10968 116016 11020 116068
rect 11244 116059 11296 116068
rect 11244 116025 11253 116059
rect 11253 116025 11287 116059
rect 11287 116025 11296 116059
rect 11244 116016 11296 116025
rect 15660 116059 15712 116068
rect 15660 116025 15669 116059
rect 15669 116025 15703 116059
rect 15703 116025 15712 116059
rect 15660 116016 15712 116025
rect 16396 116059 16448 116068
rect 16396 116025 16405 116059
rect 16405 116025 16439 116059
rect 16439 116025 16448 116059
rect 16396 116016 16448 116025
rect 20536 116016 20588 116068
rect 23020 116016 23072 116068
rect 25320 116084 25372 116136
rect 28816 116152 28868 116204
rect 30564 116152 30616 116204
rect 31484 116220 31536 116272
rect 31944 116263 31996 116272
rect 31944 116229 31953 116263
rect 31953 116229 31987 116263
rect 31987 116229 31996 116263
rect 31944 116220 31996 116229
rect 33140 116263 33192 116272
rect 33140 116229 33149 116263
rect 33149 116229 33183 116263
rect 33183 116229 33192 116263
rect 33140 116220 33192 116229
rect 35716 116220 35768 116272
rect 31116 116152 31168 116204
rect 33876 116152 33928 116204
rect 38200 116220 38252 116272
rect 37832 116195 37884 116204
rect 37832 116161 37841 116195
rect 37841 116161 37875 116195
rect 37875 116161 37884 116195
rect 37832 116152 37884 116161
rect 32128 116084 32180 116136
rect 32404 116084 32456 116136
rect 35716 116084 35768 116136
rect 37648 116127 37700 116136
rect 37648 116093 37657 116127
rect 37657 116093 37691 116127
rect 37691 116093 37700 116127
rect 37648 116084 37700 116093
rect 25872 116016 25924 116068
rect 5080 115948 5132 116000
rect 5632 115948 5684 116000
rect 20720 115948 20772 116000
rect 26148 116016 26200 116068
rect 27528 116059 27580 116068
rect 27528 116025 27537 116059
rect 27537 116025 27571 116059
rect 27571 116025 27580 116059
rect 27528 116016 27580 116025
rect 28264 116059 28316 116068
rect 28264 116025 28273 116059
rect 28273 116025 28307 116059
rect 28307 116025 28316 116059
rect 28264 116016 28316 116025
rect 29000 116059 29052 116068
rect 29000 116025 29009 116059
rect 29009 116025 29043 116059
rect 29043 116025 29052 116059
rect 29000 116016 29052 116025
rect 30656 116016 30708 116068
rect 32680 116016 32732 116068
rect 32864 116059 32916 116068
rect 32864 116025 32873 116059
rect 32873 116025 32907 116059
rect 32907 116025 32916 116059
rect 32864 116016 32916 116025
rect 34060 116016 34112 116068
rect 35256 116016 35308 116068
rect 27344 115948 27396 116000
rect 29828 115948 29880 116000
rect 19606 115846 19658 115898
rect 19670 115846 19722 115898
rect 19734 115846 19786 115898
rect 19798 115846 19850 115898
rect 1676 115744 1728 115796
rect 2412 115744 2464 115796
rect 480 115676 532 115728
rect 3424 115744 3476 115796
rect 3516 115744 3568 115796
rect 4712 115744 4764 115796
rect 7288 115744 7340 115796
rect 8392 115744 8444 115796
rect 9772 115744 9824 115796
rect 11152 115744 11204 115796
rect 14096 115744 14148 115796
rect 15844 115744 15896 115796
rect 20076 115744 20128 115796
rect 2964 115676 3016 115728
rect 2504 115608 2556 115660
rect 3608 115651 3660 115660
rect 3608 115617 3617 115651
rect 3617 115617 3651 115651
rect 3651 115617 3660 115651
rect 3608 115608 3660 115617
rect 3976 115676 4028 115728
rect 8668 115676 8720 115728
rect 11336 115676 11388 115728
rect 16580 115676 16632 115728
rect 23296 115744 23348 115796
rect 23572 115744 23624 115796
rect 24676 115744 24728 115796
rect 25964 115744 26016 115796
rect 26332 115744 26384 115796
rect 27252 115744 27304 115796
rect 29460 115744 29512 115796
rect 29736 115744 29788 115796
rect 31024 115744 31076 115796
rect 31208 115744 31260 115796
rect 35808 115744 35860 115796
rect 36084 115744 36136 115796
rect 4620 115608 4672 115660
rect 5080 115651 5132 115660
rect 5080 115617 5089 115651
rect 5089 115617 5123 115651
rect 5123 115617 5132 115651
rect 5080 115608 5132 115617
rect 6920 115608 6972 115660
rect 1584 115540 1636 115592
rect 5908 115540 5960 115592
rect 4528 115472 4580 115524
rect 4712 115472 4764 115524
rect 12164 115608 12216 115660
rect 12900 115651 12952 115660
rect 12900 115617 12909 115651
rect 12909 115617 12943 115651
rect 12943 115617 12952 115651
rect 12900 115608 12952 115617
rect 17408 115608 17460 115660
rect 21088 115608 21140 115660
rect 21640 115608 21692 115660
rect 22928 115608 22980 115660
rect 23020 115608 23072 115660
rect 23848 115608 23900 115660
rect 25412 115676 25464 115728
rect 24308 115608 24360 115660
rect 25504 115651 25556 115660
rect 25504 115617 25513 115651
rect 25513 115617 25547 115651
rect 25547 115617 25556 115651
rect 25504 115608 25556 115617
rect 26424 115651 26476 115660
rect 26424 115617 26433 115651
rect 26433 115617 26467 115651
rect 26467 115617 26476 115651
rect 26424 115608 26476 115617
rect 28724 115651 28776 115660
rect 17776 115540 17828 115592
rect 22008 115540 22060 115592
rect 22560 115540 22612 115592
rect 28724 115617 28733 115651
rect 28733 115617 28767 115651
rect 28767 115617 28776 115651
rect 28724 115608 28776 115617
rect 28816 115608 28868 115660
rect 31852 115676 31904 115728
rect 34520 115676 34572 115728
rect 35348 115719 35400 115728
rect 35348 115685 35357 115719
rect 35357 115685 35391 115719
rect 35391 115685 35400 115719
rect 35348 115676 35400 115685
rect 31576 115608 31628 115660
rect 33784 115608 33836 115660
rect 34336 115608 34388 115660
rect 34520 115540 34572 115592
rect 34888 115540 34940 115592
rect 36268 115608 36320 115660
rect 36636 115651 36688 115660
rect 36636 115617 36645 115651
rect 36645 115617 36679 115651
rect 36679 115617 36688 115651
rect 36636 115608 36688 115617
rect 35348 115540 35400 115592
rect 1952 115447 2004 115456
rect 1952 115413 1961 115447
rect 1961 115413 1995 115447
rect 1995 115413 2004 115447
rect 1952 115404 2004 115413
rect 10048 115404 10100 115456
rect 10876 115404 10928 115456
rect 21640 115472 21692 115524
rect 23204 115472 23256 115524
rect 24124 115472 24176 115524
rect 24676 115472 24728 115524
rect 25136 115404 25188 115456
rect 25872 115472 25924 115524
rect 39488 115472 39540 115524
rect 29184 115404 29236 115456
rect 29736 115404 29788 115456
rect 33416 115404 33468 115456
rect 4246 115302 4298 115354
rect 4310 115302 4362 115354
rect 4374 115302 4426 115354
rect 4438 115302 4490 115354
rect 34966 115302 35018 115354
rect 35030 115302 35082 115354
rect 35094 115302 35146 115354
rect 35158 115302 35210 115354
rect 1400 115200 1452 115252
rect 4068 115200 4120 115252
rect 5540 115200 5592 115252
rect 6276 115200 6328 115252
rect 7932 115200 7984 115252
rect 9864 115200 9916 115252
rect 10600 115200 10652 115252
rect 10968 115243 11020 115252
rect 10968 115209 10977 115243
rect 10977 115209 11011 115243
rect 11011 115209 11020 115243
rect 10968 115200 11020 115209
rect 11244 115200 11296 115252
rect 12992 115243 13044 115252
rect 12992 115209 13001 115243
rect 13001 115209 13035 115243
rect 13035 115209 13044 115243
rect 12992 115200 13044 115209
rect 14372 115200 14424 115252
rect 15108 115200 15160 115252
rect 15568 115243 15620 115252
rect 15568 115209 15577 115243
rect 15577 115209 15611 115243
rect 15611 115209 15620 115243
rect 15568 115200 15620 115209
rect 15660 115200 15712 115252
rect 16396 115200 16448 115252
rect 18144 115200 18196 115252
rect 19340 115200 19392 115252
rect 20352 115200 20404 115252
rect 20720 115200 20772 115252
rect 21640 115243 21692 115252
rect 21640 115209 21649 115243
rect 21649 115209 21683 115243
rect 21683 115209 21692 115243
rect 21640 115200 21692 115209
rect 22100 115243 22152 115252
rect 22100 115209 22109 115243
rect 22109 115209 22143 115243
rect 22143 115209 22152 115243
rect 22100 115200 22152 115209
rect 25780 115200 25832 115252
rect 26516 115200 26568 115252
rect 27620 115200 27672 115252
rect 28908 115200 28960 115252
rect 31116 115243 31168 115252
rect 2872 115132 2924 115184
rect 5356 115132 5408 115184
rect 5448 115064 5500 115116
rect 9864 115064 9916 115116
rect 18696 115132 18748 115184
rect 10692 115064 10744 115116
rect 2688 114996 2740 115048
rect 6276 114996 6328 115048
rect 10968 114996 11020 115048
rect 18880 115064 18932 115116
rect 19340 115064 19392 115116
rect 26424 115132 26476 115184
rect 15292 114996 15344 115048
rect 27528 115064 27580 115116
rect 28356 115064 28408 115116
rect 1860 114971 1912 114980
rect 1860 114937 1869 114971
rect 1869 114937 1903 114971
rect 1903 114937 1912 114971
rect 1860 114928 1912 114937
rect 5632 114971 5684 114980
rect 5632 114937 5641 114971
rect 5641 114937 5675 114971
rect 5675 114937 5684 114971
rect 5632 114928 5684 114937
rect 8024 114971 8076 114980
rect 8024 114937 8033 114971
rect 8033 114937 8067 114971
rect 8067 114937 8076 114971
rect 8024 114928 8076 114937
rect 9404 114928 9456 114980
rect 10508 114928 10560 114980
rect 11888 114928 11940 114980
rect 12900 114928 12952 114980
rect 17316 114928 17368 114980
rect 26700 115039 26752 115048
rect 8392 114860 8444 114912
rect 12532 114860 12584 114912
rect 13544 114860 13596 114912
rect 18880 114860 18932 114912
rect 20904 114860 20956 114912
rect 20996 114860 21048 114912
rect 23112 114928 23164 114980
rect 26700 115005 26709 115039
rect 26709 115005 26743 115039
rect 26743 115005 26752 115039
rect 26700 114996 26752 115005
rect 27804 114996 27856 115048
rect 31116 115209 31125 115243
rect 31125 115209 31159 115243
rect 31159 115209 31168 115243
rect 31116 115200 31168 115209
rect 31668 115200 31720 115252
rect 32404 115243 32456 115252
rect 32404 115209 32413 115243
rect 32413 115209 32447 115243
rect 32447 115209 32456 115243
rect 32404 115200 32456 115209
rect 36912 115200 36964 115252
rect 37096 115243 37148 115252
rect 37096 115209 37105 115243
rect 37105 115209 37139 115243
rect 37139 115209 37148 115243
rect 37096 115200 37148 115209
rect 32588 115132 32640 115184
rect 34520 115132 34572 115184
rect 38016 115132 38068 115184
rect 37556 115064 37608 115116
rect 32036 114996 32088 115048
rect 33968 114996 34020 115048
rect 35072 114996 35124 115048
rect 36728 114996 36780 115048
rect 37648 115039 37700 115048
rect 37648 115005 37657 115039
rect 37657 115005 37691 115039
rect 37691 115005 37700 115039
rect 37648 114996 37700 115005
rect 27712 114971 27764 114980
rect 23296 114860 23348 114912
rect 26056 114860 26108 114912
rect 27712 114937 27721 114971
rect 27721 114937 27755 114971
rect 27755 114937 27764 114971
rect 27712 114928 27764 114937
rect 29092 114928 29144 114980
rect 32404 114928 32456 114980
rect 33416 114928 33468 114980
rect 34520 114928 34572 114980
rect 35992 114928 36044 114980
rect 36912 114928 36964 114980
rect 38292 114928 38344 114980
rect 27896 114860 27948 114912
rect 30472 114903 30524 114912
rect 30472 114869 30481 114903
rect 30481 114869 30515 114903
rect 30515 114869 30524 114903
rect 30472 114860 30524 114869
rect 19606 114758 19658 114810
rect 19670 114758 19722 114810
rect 19734 114758 19786 114810
rect 19798 114758 19850 114810
rect 6644 114656 6696 114708
rect 10416 114656 10468 114708
rect 3516 114588 3568 114640
rect 14464 114656 14516 114708
rect 2412 114520 2464 114572
rect 3700 114520 3752 114572
rect 4988 114520 5040 114572
rect 5540 114520 5592 114572
rect 6552 114520 6604 114572
rect 2044 114495 2096 114504
rect 2044 114461 2053 114495
rect 2053 114461 2087 114495
rect 2087 114461 2096 114495
rect 2044 114452 2096 114461
rect 3240 114452 3292 114504
rect 4804 114452 4856 114504
rect 5724 114452 5776 114504
rect 7012 114495 7064 114504
rect 7012 114461 7021 114495
rect 7021 114461 7055 114495
rect 7055 114461 7064 114495
rect 7012 114452 7064 114461
rect 7564 114452 7616 114504
rect 3332 114316 3384 114368
rect 5080 114316 5132 114368
rect 8208 114520 8260 114572
rect 8576 114495 8628 114504
rect 8576 114461 8585 114495
rect 8585 114461 8619 114495
rect 8619 114461 8628 114495
rect 8576 114452 8628 114461
rect 10508 114563 10560 114572
rect 10508 114529 10517 114563
rect 10517 114529 10551 114563
rect 10551 114529 10560 114563
rect 10508 114520 10560 114529
rect 10876 114520 10928 114572
rect 11428 114520 11480 114572
rect 12900 114563 12952 114572
rect 12900 114529 12909 114563
rect 12909 114529 12943 114563
rect 12943 114529 12952 114563
rect 12900 114520 12952 114529
rect 13268 114520 13320 114572
rect 13544 114563 13596 114572
rect 13544 114529 13553 114563
rect 13553 114529 13587 114563
rect 13587 114529 13596 114563
rect 13544 114520 13596 114529
rect 13912 114520 13964 114572
rect 14924 114520 14976 114572
rect 17316 114699 17368 114708
rect 17316 114665 17325 114699
rect 17325 114665 17359 114699
rect 17359 114665 17368 114699
rect 17316 114656 17368 114665
rect 20720 114656 20772 114708
rect 21364 114656 21416 114708
rect 21732 114656 21784 114708
rect 22560 114699 22612 114708
rect 22560 114665 22569 114699
rect 22569 114665 22603 114699
rect 22603 114665 22612 114699
rect 22560 114656 22612 114665
rect 23664 114656 23716 114708
rect 17040 114520 17092 114572
rect 18052 114563 18104 114572
rect 18052 114529 18061 114563
rect 18061 114529 18095 114563
rect 18095 114529 18104 114563
rect 18052 114520 18104 114529
rect 18696 114563 18748 114572
rect 18696 114529 18705 114563
rect 18705 114529 18739 114563
rect 18739 114529 18748 114563
rect 18696 114520 18748 114529
rect 19432 114588 19484 114640
rect 18972 114520 19024 114572
rect 20260 114520 20312 114572
rect 20904 114520 20956 114572
rect 21824 114588 21876 114640
rect 22192 114588 22244 114640
rect 22284 114588 22336 114640
rect 22744 114563 22796 114572
rect 20720 114452 20772 114504
rect 22744 114529 22753 114563
rect 22753 114529 22787 114563
rect 22787 114529 22796 114563
rect 22744 114520 22796 114529
rect 23848 114520 23900 114572
rect 27896 114656 27948 114708
rect 29092 114656 29144 114708
rect 29552 114656 29604 114708
rect 30932 114656 30984 114708
rect 28632 114588 28684 114640
rect 8300 114384 8352 114436
rect 15292 114427 15344 114436
rect 15292 114393 15301 114427
rect 15301 114393 15335 114427
rect 15335 114393 15344 114427
rect 15292 114384 15344 114393
rect 18880 114427 18932 114436
rect 18880 114393 18889 114427
rect 18889 114393 18923 114427
rect 18923 114393 18932 114427
rect 18880 114384 18932 114393
rect 19340 114427 19392 114436
rect 19340 114393 19349 114427
rect 19349 114393 19383 114427
rect 19383 114393 19392 114427
rect 19340 114384 19392 114393
rect 26424 114563 26476 114572
rect 26424 114529 26433 114563
rect 26433 114529 26467 114563
rect 26467 114529 26476 114563
rect 26424 114520 26476 114529
rect 27988 114520 28040 114572
rect 28448 114520 28500 114572
rect 29920 114588 29972 114640
rect 30012 114520 30064 114572
rect 30288 114520 30340 114572
rect 30472 114452 30524 114504
rect 25320 114384 25372 114436
rect 26240 114427 26292 114436
rect 26240 114393 26249 114427
rect 26249 114393 26283 114427
rect 26283 114393 26292 114427
rect 26240 114384 26292 114393
rect 26700 114384 26752 114436
rect 30196 114384 30248 114436
rect 9864 114359 9916 114368
rect 9864 114325 9873 114359
rect 9873 114325 9907 114359
rect 9907 114325 9916 114359
rect 9864 114316 9916 114325
rect 10968 114359 11020 114368
rect 10968 114325 10977 114359
rect 10977 114325 11011 114359
rect 11011 114325 11020 114359
rect 10968 114316 11020 114325
rect 13360 114359 13412 114368
rect 13360 114325 13369 114359
rect 13369 114325 13403 114359
rect 13403 114325 13412 114359
rect 13360 114316 13412 114325
rect 14648 114359 14700 114368
rect 14648 114325 14657 114359
rect 14657 114325 14691 114359
rect 14691 114325 14700 114359
rect 14648 114316 14700 114325
rect 28632 114359 28684 114368
rect 28632 114325 28641 114359
rect 28641 114325 28675 114359
rect 28675 114325 28684 114359
rect 28632 114316 28684 114325
rect 30288 114316 30340 114368
rect 32772 114588 32824 114640
rect 34152 114588 34204 114640
rect 39212 114588 39264 114640
rect 32220 114520 32272 114572
rect 33232 114520 33284 114572
rect 32772 114452 32824 114504
rect 34796 114520 34848 114572
rect 36176 114520 36228 114572
rect 37096 114563 37148 114572
rect 35072 114452 35124 114504
rect 36728 114452 36780 114504
rect 37096 114529 37105 114563
rect 37105 114529 37139 114563
rect 37139 114529 37148 114563
rect 37096 114520 37148 114529
rect 39672 114452 39724 114504
rect 37372 114384 37424 114436
rect 37280 114359 37332 114368
rect 37280 114325 37289 114359
rect 37289 114325 37323 114359
rect 37323 114325 37332 114359
rect 37280 114316 37332 114325
rect 4246 114214 4298 114266
rect 4310 114214 4362 114266
rect 4374 114214 4426 114266
rect 4438 114214 4490 114266
rect 34966 114214 35018 114266
rect 35030 114214 35082 114266
rect 35094 114214 35146 114266
rect 35158 114214 35210 114266
rect 2596 114112 2648 114164
rect 4620 114112 4672 114164
rect 5632 114112 5684 114164
rect 7748 114112 7800 114164
rect 18052 114112 18104 114164
rect 20260 114112 20312 114164
rect 24492 114112 24544 114164
rect 25412 114112 25464 114164
rect 25596 114112 25648 114164
rect 28724 114112 28776 114164
rect 29644 114112 29696 114164
rect 31484 114112 31536 114164
rect 31944 114112 31996 114164
rect 32864 114112 32916 114164
rect 3608 114044 3660 114096
rect 5448 114044 5500 114096
rect 10416 113976 10468 114028
rect 22744 114044 22796 114096
rect 29368 114044 29420 114096
rect 36820 114044 36872 114096
rect 37188 114112 37240 114164
rect 38384 114044 38436 114096
rect 20720 113976 20772 114028
rect 30380 113976 30432 114028
rect 2136 113840 2188 113892
rect 8760 113908 8812 113960
rect 15752 113908 15804 113960
rect 16488 113908 16540 113960
rect 17684 113908 17736 113960
rect 18236 113908 18288 113960
rect 20168 113951 20220 113960
rect 20168 113917 20177 113951
rect 20177 113917 20211 113951
rect 20211 113917 20220 113951
rect 20168 113908 20220 113917
rect 20812 113951 20864 113960
rect 20812 113917 20821 113951
rect 20821 113917 20855 113951
rect 20855 113917 20864 113951
rect 20812 113908 20864 113917
rect 22192 113951 22244 113960
rect 8392 113840 8444 113892
rect 22192 113917 22201 113951
rect 22201 113917 22235 113951
rect 22235 113917 22244 113951
rect 22192 113908 22244 113917
rect 22836 113951 22888 113960
rect 22836 113917 22845 113951
rect 22845 113917 22879 113951
rect 22879 113917 22888 113951
rect 22836 113908 22888 113917
rect 23388 113908 23440 113960
rect 24032 113908 24084 113960
rect 26148 113908 26200 113960
rect 28632 113908 28684 113960
rect 29276 113908 29328 113960
rect 30104 113908 30156 113960
rect 33048 113976 33100 114028
rect 33968 113976 34020 114028
rect 35808 113976 35860 114028
rect 37372 114019 37424 114028
rect 37372 113985 37381 114019
rect 37381 113985 37415 114019
rect 37415 113985 37424 114019
rect 37372 113976 37424 113985
rect 32496 113908 32548 113960
rect 33692 113908 33744 113960
rect 35532 113908 35584 113960
rect 1952 113815 2004 113824
rect 1952 113781 1961 113815
rect 1961 113781 1995 113815
rect 1995 113781 2004 113815
rect 1952 113772 2004 113781
rect 3884 113772 3936 113824
rect 31576 113840 31628 113892
rect 35348 113840 35400 113892
rect 37464 113840 37516 113892
rect 25412 113772 25464 113824
rect 34060 113772 34112 113824
rect 19606 113670 19658 113722
rect 19670 113670 19722 113722
rect 19734 113670 19786 113722
rect 19798 113670 19850 113722
rect 5172 113568 5224 113620
rect 5264 113568 5316 113620
rect 1768 113432 1820 113484
rect 2320 113475 2372 113484
rect 2320 113441 2329 113475
rect 2329 113441 2363 113475
rect 2363 113441 2372 113475
rect 2320 113432 2372 113441
rect 3056 113432 3108 113484
rect 3148 113432 3200 113484
rect 6644 113500 6696 113552
rect 6276 113432 6328 113484
rect 8300 113568 8352 113620
rect 30748 113611 30800 113620
rect 30748 113577 30757 113611
rect 30757 113577 30791 113611
rect 30791 113577 30800 113611
rect 30748 113568 30800 113577
rect 32680 113568 32732 113620
rect 38568 113568 38620 113620
rect 7472 113500 7524 113552
rect 8208 113500 8260 113552
rect 14648 113500 14700 113552
rect 36360 113500 36412 113552
rect 37004 113500 37056 113552
rect 8392 113432 8444 113484
rect 24584 113475 24636 113484
rect 24584 113441 24593 113475
rect 24593 113441 24627 113475
rect 24627 113441 24636 113475
rect 24584 113432 24636 113441
rect 25228 113475 25280 113484
rect 25228 113441 25237 113475
rect 25237 113441 25271 113475
rect 25271 113441 25280 113475
rect 25228 113432 25280 113441
rect 30840 113432 30892 113484
rect 31300 113432 31352 113484
rect 32956 113432 33008 113484
rect 33600 113432 33652 113484
rect 34520 113432 34572 113484
rect 35716 113475 35768 113484
rect 35716 113441 35725 113475
rect 35725 113441 35759 113475
rect 35759 113441 35768 113475
rect 35716 113432 35768 113441
rect 36084 113432 36136 113484
rect 13360 113364 13412 113416
rect 21640 113364 21692 113416
rect 4712 113296 4764 113348
rect 6736 113296 6788 113348
rect 8116 113339 8168 113348
rect 8116 113305 8125 113339
rect 8125 113305 8159 113339
rect 8159 113305 8168 113339
rect 8116 113296 8168 113305
rect 30656 113296 30708 113348
rect 32128 113296 32180 113348
rect 37372 113339 37424 113348
rect 37372 113305 37381 113339
rect 37381 113305 37415 113339
rect 37415 113305 37424 113339
rect 37372 113296 37424 113305
rect 4246 113126 4298 113178
rect 4310 113126 4362 113178
rect 4374 113126 4426 113178
rect 4438 113126 4490 113178
rect 34966 113126 35018 113178
rect 35030 113126 35082 113178
rect 35094 113126 35146 113178
rect 35158 113126 35210 113178
rect 30564 113024 30616 113076
rect 33140 113024 33192 113076
rect 33876 113024 33928 113076
rect 36544 113067 36596 113076
rect 36544 113033 36553 113067
rect 36553 113033 36587 113067
rect 36587 113033 36596 113067
rect 36544 113024 36596 113033
rect 6828 112956 6880 113008
rect 28540 112956 28592 113008
rect 1676 112888 1728 112940
rect 1860 112863 1912 112872
rect 1860 112829 1869 112863
rect 1869 112829 1903 112863
rect 1903 112829 1912 112863
rect 1860 112820 1912 112829
rect 3792 112820 3844 112872
rect 4896 112863 4948 112872
rect 4896 112829 4905 112863
rect 4905 112829 4939 112863
rect 4939 112829 4948 112863
rect 4896 112820 4948 112829
rect 5540 112863 5592 112872
rect 5540 112829 5549 112863
rect 5549 112829 5583 112863
rect 5583 112829 5592 112863
rect 5540 112820 5592 112829
rect 5816 112820 5868 112872
rect 6276 112820 6328 112872
rect 31024 112888 31076 112940
rect 28172 112863 28224 112872
rect 28172 112829 28181 112863
rect 28181 112829 28215 112863
rect 28215 112829 28224 112863
rect 28172 112820 28224 112829
rect 29828 112820 29880 112872
rect 31392 112820 31444 112872
rect 33324 112820 33376 112872
rect 33600 112820 33652 112872
rect 31944 112752 31996 112804
rect 36360 112752 36412 112804
rect 37372 112795 37424 112804
rect 37372 112761 37381 112795
rect 37381 112761 37415 112795
rect 37415 112761 37424 112795
rect 37372 112752 37424 112761
rect 38108 112795 38160 112804
rect 38108 112761 38117 112795
rect 38117 112761 38151 112795
rect 38151 112761 38160 112795
rect 38108 112752 38160 112761
rect 16028 112684 16080 112736
rect 26240 112684 26292 112736
rect 33140 112684 33192 112736
rect 34244 112684 34296 112736
rect 19606 112582 19658 112634
rect 19670 112582 19722 112634
rect 19734 112582 19786 112634
rect 19798 112582 19850 112634
rect 35808 112480 35860 112532
rect 20720 112412 20772 112464
rect 12716 112344 12768 112396
rect 23572 112412 23624 112464
rect 35992 112412 36044 112464
rect 39856 112412 39908 112464
rect 34428 112208 34480 112260
rect 1952 112183 2004 112192
rect 1952 112149 1961 112183
rect 1961 112149 1995 112183
rect 1995 112149 2004 112183
rect 1952 112140 2004 112149
rect 23296 112140 23348 112192
rect 36820 112344 36872 112396
rect 4246 112038 4298 112090
rect 4310 112038 4362 112090
rect 4374 112038 4426 112090
rect 4438 112038 4490 112090
rect 34966 112038 35018 112090
rect 35030 112038 35082 112090
rect 35094 112038 35146 112090
rect 35158 112038 35210 112090
rect 35532 111800 35584 111852
rect 35808 111800 35860 111852
rect 37648 111775 37700 111784
rect 37648 111741 37657 111775
rect 37657 111741 37691 111775
rect 37691 111741 37700 111775
rect 37648 111732 37700 111741
rect 35532 111664 35584 111716
rect 19606 111494 19658 111546
rect 19670 111494 19722 111546
rect 19734 111494 19786 111546
rect 19798 111494 19850 111546
rect 33784 111392 33836 111444
rect 36544 111435 36596 111444
rect 36544 111401 36553 111435
rect 36553 111401 36587 111435
rect 36587 111401 36596 111435
rect 36544 111392 36596 111401
rect 25320 111324 25372 111376
rect 34520 111324 34572 111376
rect 1400 111299 1452 111308
rect 1400 111265 1409 111299
rect 1409 111265 1443 111299
rect 1443 111265 1452 111299
rect 1400 111256 1452 111265
rect 31484 111256 31536 111308
rect 36452 111299 36504 111308
rect 36452 111265 36461 111299
rect 36461 111265 36495 111299
rect 36495 111265 36504 111299
rect 36452 111256 36504 111265
rect 7656 111188 7708 111240
rect 31116 111188 31168 111240
rect 26792 111120 26844 111172
rect 37372 111163 37424 111172
rect 34612 111052 34664 111104
rect 35900 111052 35952 111104
rect 37372 111129 37381 111163
rect 37381 111129 37415 111163
rect 37415 111129 37424 111163
rect 37372 111120 37424 111129
rect 37464 111052 37516 111104
rect 4246 110950 4298 111002
rect 4310 110950 4362 111002
rect 4374 110950 4426 111002
rect 4438 110950 4490 111002
rect 34966 110950 35018 111002
rect 35030 110950 35082 111002
rect 35094 110950 35146 111002
rect 35158 110950 35210 111002
rect 28264 110848 28316 110900
rect 36452 110848 36504 110900
rect 36268 110712 36320 110764
rect 36452 110712 36504 110764
rect 37464 110687 37516 110696
rect 37464 110653 37473 110687
rect 37473 110653 37507 110687
rect 37507 110653 37516 110687
rect 37464 110644 37516 110653
rect 2228 110576 2280 110628
rect 37832 110619 37884 110628
rect 37832 110585 37841 110619
rect 37841 110585 37875 110619
rect 37875 110585 37884 110619
rect 37832 110576 37884 110585
rect 1952 110551 2004 110560
rect 1952 110517 1961 110551
rect 1961 110517 1995 110551
rect 1995 110517 2004 110551
rect 1952 110508 2004 110517
rect 19606 110406 19658 110458
rect 19670 110406 19722 110458
rect 19734 110406 19786 110458
rect 19798 110406 19850 110458
rect 37188 110211 37240 110220
rect 37188 110177 37197 110211
rect 37197 110177 37231 110211
rect 37231 110177 37240 110211
rect 37188 110168 37240 110177
rect 22560 110032 22612 110084
rect 32772 110032 32824 110084
rect 38200 110032 38252 110084
rect 26700 109964 26752 110016
rect 36912 109964 36964 110016
rect 4246 109862 4298 109914
rect 4310 109862 4362 109914
rect 4374 109862 4426 109914
rect 4438 109862 4490 109914
rect 34966 109862 35018 109914
rect 35030 109862 35082 109914
rect 35094 109862 35146 109914
rect 35158 109862 35210 109914
rect 24676 109760 24728 109812
rect 37832 109760 37884 109812
rect 5264 109692 5316 109744
rect 26240 109692 26292 109744
rect 27620 109692 27672 109744
rect 36176 109692 36228 109744
rect 2044 109599 2096 109608
rect 2044 109565 2053 109599
rect 2053 109565 2087 109599
rect 2087 109565 2096 109599
rect 2044 109556 2096 109565
rect 37188 109599 37240 109608
rect 37188 109565 37197 109599
rect 37197 109565 37231 109599
rect 37231 109565 37240 109599
rect 37188 109556 37240 109565
rect 11060 109488 11112 109540
rect 37924 109531 37976 109540
rect 37924 109497 37933 109531
rect 37933 109497 37967 109531
rect 37967 109497 37976 109531
rect 37924 109488 37976 109497
rect 38660 109488 38712 109540
rect 38384 109420 38436 109472
rect 19606 109318 19658 109370
rect 19670 109318 19722 109370
rect 19734 109318 19786 109370
rect 19798 109318 19850 109370
rect 8668 109259 8720 109268
rect 8668 109225 8677 109259
rect 8677 109225 8711 109259
rect 8711 109225 8720 109259
rect 8668 109216 8720 109225
rect 13084 109080 13136 109132
rect 37188 109123 37240 109132
rect 37188 109089 37197 109123
rect 37197 109089 37231 109123
rect 37231 109089 37240 109123
rect 37188 109080 37240 109089
rect 2504 109012 2556 109064
rect 3424 109012 3476 109064
rect 32680 109012 32732 109064
rect 4246 108774 4298 108826
rect 4310 108774 4362 108826
rect 4374 108774 4426 108826
rect 4438 108774 4490 108826
rect 34966 108774 35018 108826
rect 35030 108774 35082 108826
rect 35094 108774 35146 108826
rect 35158 108774 35210 108826
rect 1952 108715 2004 108724
rect 1952 108681 1961 108715
rect 1961 108681 1995 108715
rect 1995 108681 2004 108715
rect 1952 108672 2004 108681
rect 32772 108468 32824 108520
rect 7564 108400 7616 108452
rect 21548 108400 21600 108452
rect 33232 108400 33284 108452
rect 37924 108443 37976 108452
rect 37924 108409 37933 108443
rect 37933 108409 37967 108443
rect 37967 108409 37976 108443
rect 37924 108400 37976 108409
rect 23112 108332 23164 108384
rect 31944 108332 31996 108384
rect 19606 108230 19658 108282
rect 19670 108230 19722 108282
rect 19734 108230 19786 108282
rect 19798 108230 19850 108282
rect 13452 107992 13504 108044
rect 37188 108035 37240 108044
rect 37188 108001 37197 108035
rect 37197 108001 37231 108035
rect 37231 108001 37240 108035
rect 37188 107992 37240 108001
rect 2044 107899 2096 107908
rect 2044 107865 2053 107899
rect 2053 107865 2087 107899
rect 2087 107865 2096 107899
rect 2044 107856 2096 107865
rect 33232 107788 33284 107840
rect 4246 107686 4298 107738
rect 4310 107686 4362 107738
rect 4374 107686 4426 107738
rect 4438 107686 4490 107738
rect 34966 107686 35018 107738
rect 35030 107686 35082 107738
rect 35094 107686 35146 107738
rect 35158 107686 35210 107738
rect 32956 107584 33008 107636
rect 37372 107584 37424 107636
rect 37188 107423 37240 107432
rect 37188 107389 37197 107423
rect 37197 107389 37231 107423
rect 37231 107389 37240 107423
rect 37188 107380 37240 107389
rect 37556 107312 37608 107364
rect 37924 107355 37976 107364
rect 37924 107321 37933 107355
rect 37933 107321 37967 107355
rect 37967 107321 37976 107355
rect 37924 107312 37976 107321
rect 36912 107244 36964 107296
rect 19606 107142 19658 107194
rect 19670 107142 19722 107194
rect 19734 107142 19786 107194
rect 19798 107142 19850 107194
rect 1952 107083 2004 107092
rect 1952 107049 1961 107083
rect 1961 107049 1995 107083
rect 1995 107049 2004 107083
rect 1952 107040 2004 107049
rect 24032 106972 24084 107024
rect 37832 106972 37884 107024
rect 7748 106904 7800 106956
rect 22468 106904 22520 106956
rect 32404 106904 32456 106956
rect 37188 106947 37240 106956
rect 37188 106913 37197 106947
rect 37197 106913 37231 106947
rect 37231 106913 37240 106947
rect 37188 106904 37240 106913
rect 38476 106768 38528 106820
rect 4246 106598 4298 106650
rect 4310 106598 4362 106650
rect 4374 106598 4426 106650
rect 4438 106598 4490 106650
rect 34966 106598 35018 106650
rect 35030 106598 35082 106650
rect 35094 106598 35146 106650
rect 35158 106598 35210 106650
rect 1768 106335 1820 106344
rect 1768 106301 1777 106335
rect 1777 106301 1811 106335
rect 1811 106301 1820 106335
rect 1768 106292 1820 106301
rect 29644 106360 29696 106412
rect 36544 106360 36596 106412
rect 32864 106292 32916 106344
rect 33232 106292 33284 106344
rect 37280 106335 37332 106344
rect 37280 106301 37289 106335
rect 37289 106301 37323 106335
rect 37323 106301 37332 106335
rect 37280 106292 37332 106301
rect 19606 106054 19658 106106
rect 19670 106054 19722 106106
rect 19734 106054 19786 106106
rect 19798 106054 19850 106106
rect 37188 105859 37240 105868
rect 37188 105825 37197 105859
rect 37197 105825 37231 105859
rect 37231 105825 37240 105859
rect 37188 105816 37240 105825
rect 25964 105680 26016 105732
rect 35808 105680 35860 105732
rect 33324 105612 33376 105664
rect 4246 105510 4298 105562
rect 4310 105510 4362 105562
rect 4374 105510 4426 105562
rect 4438 105510 4490 105562
rect 34966 105510 35018 105562
rect 35030 105510 35082 105562
rect 35094 105510 35146 105562
rect 35158 105510 35210 105562
rect 27620 105408 27672 105460
rect 36084 105408 36136 105460
rect 1400 105247 1452 105256
rect 1400 105213 1409 105247
rect 1409 105213 1443 105247
rect 1443 105213 1452 105247
rect 1400 105204 1452 105213
rect 24860 105204 24912 105256
rect 26056 105247 26108 105256
rect 20628 105136 20680 105188
rect 26056 105213 26065 105247
rect 26065 105213 26099 105247
rect 26099 105213 26108 105247
rect 26056 105204 26108 105213
rect 32036 105247 32088 105256
rect 32036 105213 32045 105247
rect 32045 105213 32079 105247
rect 32079 105213 32088 105247
rect 32036 105204 32088 105213
rect 37188 105247 37240 105256
rect 37188 105213 37197 105247
rect 37197 105213 37231 105247
rect 37231 105213 37240 105247
rect 37188 105204 37240 105213
rect 37924 105179 37976 105188
rect 37924 105145 37933 105179
rect 37933 105145 37967 105179
rect 37967 105145 37976 105179
rect 37924 105136 37976 105145
rect 8944 105068 8996 105120
rect 34152 105068 34204 105120
rect 38016 105111 38068 105120
rect 38016 105077 38025 105111
rect 38025 105077 38059 105111
rect 38059 105077 38068 105111
rect 38016 105068 38068 105077
rect 19606 104966 19658 105018
rect 19670 104966 19722 105018
rect 19734 104966 19786 105018
rect 19798 104966 19850 105018
rect 25964 104907 26016 104916
rect 25964 104873 25973 104907
rect 25973 104873 26007 104907
rect 26007 104873 26016 104907
rect 25964 104864 26016 104873
rect 20444 104796 20496 104848
rect 1860 104771 1912 104780
rect 1860 104737 1869 104771
rect 1869 104737 1903 104771
rect 1903 104737 1912 104771
rect 1860 104728 1912 104737
rect 24860 104771 24912 104780
rect 24860 104737 24869 104771
rect 24869 104737 24903 104771
rect 24903 104737 24912 104771
rect 24860 104728 24912 104737
rect 26056 104796 26108 104848
rect 37188 104771 37240 104780
rect 21272 104660 21324 104712
rect 37188 104737 37197 104771
rect 37197 104737 37231 104771
rect 37231 104737 37240 104771
rect 37188 104728 37240 104737
rect 10324 104524 10376 104576
rect 37004 104524 37056 104576
rect 4246 104422 4298 104474
rect 4310 104422 4362 104474
rect 4374 104422 4426 104474
rect 4438 104422 4490 104474
rect 34966 104422 35018 104474
rect 35030 104422 35082 104474
rect 35094 104422 35146 104474
rect 35158 104422 35210 104474
rect 35348 104320 35400 104372
rect 24952 104184 25004 104236
rect 31392 104184 31444 104236
rect 26884 104116 26936 104168
rect 34244 104116 34296 104168
rect 38016 104116 38068 104168
rect 37188 104091 37240 104100
rect 37188 104057 37197 104091
rect 37197 104057 37231 104091
rect 37231 104057 37240 104091
rect 37188 104048 37240 104057
rect 37372 104091 37424 104100
rect 37372 104057 37381 104091
rect 37381 104057 37415 104091
rect 37415 104057 37424 104091
rect 37372 104048 37424 104057
rect 37924 104091 37976 104100
rect 37924 104057 37933 104091
rect 37933 104057 37967 104091
rect 37967 104057 37976 104091
rect 37924 104048 37976 104057
rect 38016 104023 38068 104032
rect 38016 103989 38025 104023
rect 38025 103989 38059 104023
rect 38059 103989 38068 104023
rect 38016 103980 38068 103989
rect 19606 103878 19658 103930
rect 19670 103878 19722 103930
rect 19734 103878 19786 103930
rect 19798 103878 19850 103930
rect 11060 103776 11112 103828
rect 21272 103819 21324 103828
rect 1860 103751 1912 103760
rect 1860 103717 1869 103751
rect 1869 103717 1903 103751
rect 1903 103717 1912 103751
rect 1860 103708 1912 103717
rect 12532 103683 12584 103692
rect 12532 103649 12541 103683
rect 12541 103649 12575 103683
rect 12575 103649 12584 103683
rect 12532 103640 12584 103649
rect 12624 103640 12676 103692
rect 21272 103785 21281 103819
rect 21281 103785 21315 103819
rect 21315 103785 21324 103819
rect 21272 103776 21324 103785
rect 21640 103819 21692 103828
rect 21640 103785 21649 103819
rect 21649 103785 21683 103819
rect 21683 103785 21692 103819
rect 21640 103776 21692 103785
rect 18328 103708 18380 103760
rect 20444 103708 20496 103760
rect 20536 103708 20588 103760
rect 24860 103708 24912 103760
rect 26792 103708 26844 103760
rect 14464 103640 14516 103692
rect 37188 103683 37240 103692
rect 37188 103649 37197 103683
rect 37197 103649 37231 103683
rect 37231 103649 37240 103683
rect 37188 103640 37240 103649
rect 18052 103572 18104 103624
rect 9036 103504 9088 103556
rect 31208 103572 31260 103624
rect 32312 103504 32364 103556
rect 36912 103504 36964 103556
rect 13544 103436 13596 103488
rect 16580 103436 16632 103488
rect 18328 103436 18380 103488
rect 19340 103436 19392 103488
rect 4246 103334 4298 103386
rect 4310 103334 4362 103386
rect 4374 103334 4426 103386
rect 4438 103334 4490 103386
rect 34966 103334 35018 103386
rect 35030 103334 35082 103386
rect 35094 103334 35146 103386
rect 35158 103334 35210 103386
rect 3516 103232 3568 103284
rect 2044 103164 2096 103216
rect 31300 103164 31352 103216
rect 36084 103096 36136 103148
rect 6184 103071 6236 103080
rect 6184 103037 6193 103071
rect 6193 103037 6227 103071
rect 6227 103037 6236 103071
rect 6184 103028 6236 103037
rect 6828 103071 6880 103080
rect 6828 103037 6837 103071
rect 6837 103037 6871 103071
rect 6871 103037 6880 103071
rect 6828 103028 6880 103037
rect 37280 103071 37332 103080
rect 37280 103037 37289 103071
rect 37289 103037 37323 103071
rect 37323 103037 37332 103071
rect 37280 103028 37332 103037
rect 1860 103003 1912 103012
rect 1860 102969 1869 103003
rect 1869 102969 1903 103003
rect 1903 102969 1912 103003
rect 1860 102960 1912 102969
rect 4804 102960 4856 103012
rect 15200 102960 15252 103012
rect 19606 102790 19658 102842
rect 19670 102790 19722 102842
rect 19734 102790 19786 102842
rect 19798 102790 19850 102842
rect 2688 102688 2740 102740
rect 12440 102731 12492 102740
rect 12440 102697 12449 102731
rect 12449 102697 12483 102731
rect 12483 102697 12492 102731
rect 12440 102688 12492 102697
rect 13544 102688 13596 102740
rect 26792 102731 26844 102740
rect 26792 102697 26801 102731
rect 26801 102697 26835 102731
rect 26835 102697 26844 102731
rect 26792 102688 26844 102697
rect 12624 102620 12676 102672
rect 13176 102552 13228 102604
rect 26700 102595 26752 102604
rect 26700 102561 26709 102595
rect 26709 102561 26743 102595
rect 26743 102561 26752 102595
rect 26700 102552 26752 102561
rect 37188 102595 37240 102604
rect 37188 102561 37197 102595
rect 37197 102561 37231 102595
rect 37231 102561 37240 102595
rect 37188 102552 37240 102561
rect 12072 102527 12124 102536
rect 12072 102493 12081 102527
rect 12081 102493 12115 102527
rect 12115 102493 12124 102527
rect 12072 102484 12124 102493
rect 12532 102527 12584 102536
rect 12532 102493 12566 102527
rect 12566 102493 12584 102527
rect 12532 102484 12584 102493
rect 7564 102416 7616 102468
rect 13360 102348 13412 102400
rect 37280 102391 37332 102400
rect 37280 102357 37289 102391
rect 37289 102357 37323 102391
rect 37323 102357 37332 102391
rect 37280 102348 37332 102357
rect 4246 102246 4298 102298
rect 4310 102246 4362 102298
rect 4374 102246 4426 102298
rect 4438 102246 4490 102298
rect 34966 102246 35018 102298
rect 35030 102246 35082 102298
rect 35094 102246 35146 102298
rect 35158 102246 35210 102298
rect 32496 102144 32548 102196
rect 36544 102144 36596 102196
rect 36912 102144 36964 102196
rect 38016 102144 38068 102196
rect 7748 102076 7800 102128
rect 13452 102119 13504 102128
rect 13452 102085 13461 102119
rect 13461 102085 13495 102119
rect 13495 102085 13504 102119
rect 13452 102076 13504 102085
rect 12624 102008 12676 102060
rect 13544 102008 13596 102060
rect 1860 101983 1912 101992
rect 1860 101949 1869 101983
rect 1869 101949 1903 101983
rect 1903 101949 1912 101983
rect 1860 101940 1912 101949
rect 12072 101940 12124 101992
rect 18052 101940 18104 101992
rect 2044 101915 2096 101924
rect 2044 101881 2053 101915
rect 2053 101881 2087 101915
rect 2087 101881 2096 101915
rect 2044 101872 2096 101881
rect 12256 101872 12308 101924
rect 19432 101872 19484 101924
rect 37924 101915 37976 101924
rect 37924 101881 37933 101915
rect 37933 101881 37967 101915
rect 37967 101881 37976 101915
rect 37924 101872 37976 101881
rect 12440 101804 12492 101856
rect 12624 101804 12676 101856
rect 20628 101804 20680 101856
rect 30472 101804 30524 101856
rect 19606 101702 19658 101754
rect 19670 101702 19722 101754
rect 19734 101702 19786 101754
rect 19798 101702 19850 101754
rect 2136 101600 2188 101652
rect 12440 101643 12492 101652
rect 12440 101609 12449 101643
rect 12449 101609 12483 101643
rect 12483 101609 12492 101643
rect 12716 101643 12768 101652
rect 12440 101600 12492 101609
rect 12716 101609 12725 101643
rect 12725 101609 12759 101643
rect 12759 101609 12768 101643
rect 12716 101600 12768 101609
rect 23296 101643 23348 101652
rect 23296 101609 23305 101643
rect 23305 101609 23339 101643
rect 23339 101609 23348 101643
rect 23296 101600 23348 101609
rect 12624 101532 12676 101584
rect 1860 101507 1912 101516
rect 1860 101473 1869 101507
rect 1869 101473 1903 101507
rect 1903 101473 1912 101507
rect 1860 101464 1912 101473
rect 5724 101507 5776 101516
rect 5724 101473 5733 101507
rect 5733 101473 5767 101507
rect 5767 101473 5776 101507
rect 5724 101464 5776 101473
rect 12900 101464 12952 101516
rect 17224 101464 17276 101516
rect 37188 101507 37240 101516
rect 37188 101473 37197 101507
rect 37197 101473 37231 101507
rect 37231 101473 37240 101507
rect 37188 101464 37240 101473
rect 2412 101396 2464 101448
rect 10876 101396 10928 101448
rect 12532 101439 12584 101448
rect 12532 101405 12566 101439
rect 12566 101405 12584 101439
rect 12532 101396 12584 101405
rect 21456 101396 21508 101448
rect 31116 101396 31168 101448
rect 35348 101396 35400 101448
rect 36636 101396 36688 101448
rect 4068 101328 4120 101380
rect 36544 101260 36596 101312
rect 4246 101158 4298 101210
rect 4310 101158 4362 101210
rect 4374 101158 4426 101210
rect 4438 101158 4490 101210
rect 34966 101158 35018 101210
rect 35030 101158 35082 101210
rect 35094 101158 35146 101210
rect 35158 101158 35210 101210
rect 32128 100920 32180 100972
rect 37372 100920 37424 100972
rect 19432 100852 19484 100904
rect 20536 100852 20588 100904
rect 37924 100895 37976 100904
rect 37924 100861 37933 100895
rect 37933 100861 37967 100895
rect 37967 100861 37976 100895
rect 37924 100852 37976 100861
rect 37188 100827 37240 100836
rect 37188 100793 37197 100827
rect 37197 100793 37231 100827
rect 37231 100793 37240 100827
rect 37188 100784 37240 100793
rect 37648 100784 37700 100836
rect 36728 100716 36780 100768
rect 19606 100614 19658 100666
rect 19670 100614 19722 100666
rect 19734 100614 19786 100666
rect 19798 100614 19850 100666
rect 23112 100555 23164 100564
rect 23112 100521 23121 100555
rect 23121 100521 23155 100555
rect 23155 100521 23164 100555
rect 23112 100512 23164 100521
rect 1860 100487 1912 100496
rect 1860 100453 1869 100487
rect 1869 100453 1903 100487
rect 1903 100453 1912 100487
rect 1860 100444 1912 100453
rect 15936 100376 15988 100428
rect 37188 100419 37240 100428
rect 37188 100385 37197 100419
rect 37197 100385 37231 100419
rect 37231 100385 37240 100419
rect 37188 100376 37240 100385
rect 17316 100172 17368 100224
rect 31116 100172 31168 100224
rect 4246 100070 4298 100122
rect 4310 100070 4362 100122
rect 4374 100070 4426 100122
rect 4438 100070 4490 100122
rect 34966 100070 35018 100122
rect 35030 100070 35082 100122
rect 35094 100070 35146 100122
rect 35158 100070 35210 100122
rect 5724 99968 5776 100020
rect 12072 99968 12124 100020
rect 32220 99968 32272 100020
rect 35624 99900 35676 99952
rect 29644 99764 29696 99816
rect 1860 99739 1912 99748
rect 1860 99705 1869 99739
rect 1869 99705 1903 99739
rect 1903 99705 1912 99739
rect 1860 99696 1912 99705
rect 6276 99696 6328 99748
rect 18604 99696 18656 99748
rect 31024 99696 31076 99748
rect 33600 99739 33652 99748
rect 33600 99705 33609 99739
rect 33609 99705 33643 99739
rect 33643 99705 33652 99739
rect 33600 99696 33652 99705
rect 34428 99739 34480 99748
rect 34428 99705 34437 99739
rect 34437 99705 34471 99739
rect 34471 99705 34480 99739
rect 34428 99696 34480 99705
rect 37924 99739 37976 99748
rect 37924 99705 37933 99739
rect 37933 99705 37967 99739
rect 37967 99705 37976 99739
rect 37924 99696 37976 99705
rect 37832 99628 37884 99680
rect 19606 99526 19658 99578
rect 19670 99526 19722 99578
rect 19734 99526 19786 99578
rect 19798 99526 19850 99578
rect 13728 99356 13780 99408
rect 15200 99356 15252 99408
rect 29644 99356 29696 99408
rect 29920 99356 29972 99408
rect 16396 99288 16448 99340
rect 37188 99331 37240 99340
rect 37188 99297 37197 99331
rect 37197 99297 37231 99331
rect 37231 99297 37240 99331
rect 37188 99288 37240 99297
rect 12900 99263 12952 99272
rect 12900 99229 12909 99263
rect 12909 99229 12943 99263
rect 12943 99229 12952 99263
rect 12900 99220 12952 99229
rect 13176 99263 13228 99272
rect 13176 99229 13185 99263
rect 13185 99229 13219 99263
rect 13219 99229 13228 99263
rect 13176 99220 13228 99229
rect 15200 99220 15252 99272
rect 20076 99152 20128 99204
rect 3424 99084 3476 99136
rect 31576 99084 31628 99136
rect 4246 98982 4298 99034
rect 4310 98982 4362 99034
rect 4374 98982 4426 99034
rect 4438 98982 4490 99034
rect 34966 98982 35018 99034
rect 35030 98982 35082 99034
rect 35094 98982 35146 99034
rect 35158 98982 35210 99034
rect 21456 98855 21508 98864
rect 21456 98821 21465 98855
rect 21465 98821 21499 98855
rect 21499 98821 21508 98855
rect 21456 98812 21508 98821
rect 28264 98812 28316 98864
rect 1860 98719 1912 98728
rect 1860 98685 1869 98719
rect 1869 98685 1903 98719
rect 1903 98685 1912 98719
rect 1860 98676 1912 98685
rect 13820 98676 13872 98728
rect 26700 98676 26752 98728
rect 37188 98719 37240 98728
rect 37188 98685 37197 98719
rect 37197 98685 37231 98719
rect 37231 98685 37240 98719
rect 37188 98676 37240 98685
rect 3516 98608 3568 98660
rect 21272 98651 21324 98660
rect 21272 98617 21281 98651
rect 21281 98617 21315 98651
rect 21315 98617 21324 98651
rect 21272 98608 21324 98617
rect 22008 98651 22060 98660
rect 22008 98617 22017 98651
rect 22017 98617 22051 98651
rect 22051 98617 22060 98651
rect 22008 98608 22060 98617
rect 23664 98608 23716 98660
rect 31484 98608 31536 98660
rect 37740 98608 37792 98660
rect 37924 98651 37976 98660
rect 37924 98617 37933 98651
rect 37933 98617 37967 98651
rect 37967 98617 37976 98651
rect 37924 98608 37976 98617
rect 36636 98540 36688 98592
rect 19606 98438 19658 98490
rect 19670 98438 19722 98490
rect 19734 98438 19786 98490
rect 19798 98438 19850 98490
rect 2228 98336 2280 98388
rect 1860 98243 1912 98252
rect 1860 98209 1869 98243
rect 1869 98209 1903 98243
rect 1903 98209 1912 98243
rect 1860 98200 1912 98209
rect 4988 98243 5040 98252
rect 4988 98209 4997 98243
rect 4997 98209 5031 98243
rect 5031 98209 5040 98243
rect 4988 98200 5040 98209
rect 37188 98243 37240 98252
rect 37188 98209 37197 98243
rect 37197 98209 37231 98243
rect 37231 98209 37240 98243
rect 37188 98200 37240 98209
rect 9128 98064 9180 98116
rect 32404 98064 32456 98116
rect 33324 98064 33376 98116
rect 35624 98064 35676 98116
rect 36820 98064 36872 98116
rect 29460 97996 29512 98048
rect 4246 97894 4298 97946
rect 4310 97894 4362 97946
rect 4374 97894 4426 97946
rect 4438 97894 4490 97946
rect 34966 97894 35018 97946
rect 35030 97894 35082 97946
rect 35094 97894 35146 97946
rect 35158 97894 35210 97946
rect 16580 97767 16632 97776
rect 16580 97733 16589 97767
rect 16589 97733 16623 97767
rect 16623 97733 16632 97767
rect 16580 97724 16632 97733
rect 16396 97631 16448 97640
rect 16396 97597 16405 97631
rect 16405 97597 16439 97631
rect 16439 97597 16448 97631
rect 16396 97588 16448 97597
rect 18236 97588 18288 97640
rect 37924 97631 37976 97640
rect 37924 97597 37933 97631
rect 37933 97597 37967 97631
rect 37967 97597 37976 97631
rect 37924 97588 37976 97597
rect 15200 97520 15252 97572
rect 15844 97520 15896 97572
rect 12532 97452 12584 97504
rect 15108 97495 15160 97504
rect 15108 97461 15117 97495
rect 15117 97461 15151 97495
rect 15151 97461 15160 97495
rect 15108 97452 15160 97461
rect 33508 97452 33560 97504
rect 19606 97350 19658 97402
rect 19670 97350 19722 97402
rect 19734 97350 19786 97402
rect 19798 97350 19850 97402
rect 6828 97248 6880 97300
rect 14004 97248 14056 97300
rect 1860 97155 1912 97164
rect 1860 97121 1869 97155
rect 1869 97121 1903 97155
rect 1903 97121 1912 97155
rect 1860 97112 1912 97121
rect 37188 97155 37240 97164
rect 37188 97121 37197 97155
rect 37197 97121 37231 97155
rect 37231 97121 37240 97155
rect 37188 97112 37240 97121
rect 11704 96908 11756 96960
rect 31300 96908 31352 96960
rect 4246 96806 4298 96858
rect 4310 96806 4362 96858
rect 4374 96806 4426 96858
rect 4438 96806 4490 96858
rect 34966 96806 35018 96858
rect 35030 96806 35082 96858
rect 35094 96806 35146 96858
rect 35158 96806 35210 96858
rect 19340 96704 19392 96756
rect 18236 96543 18288 96552
rect 18236 96509 18245 96543
rect 18245 96509 18279 96543
rect 18279 96509 18288 96543
rect 18236 96500 18288 96509
rect 37188 96543 37240 96552
rect 37188 96509 37197 96543
rect 37197 96509 37231 96543
rect 37231 96509 37240 96543
rect 37188 96500 37240 96509
rect 37924 96543 37976 96552
rect 37924 96509 37933 96543
rect 37933 96509 37967 96543
rect 37967 96509 37976 96543
rect 37924 96500 37976 96509
rect 1860 96475 1912 96484
rect 1860 96441 1869 96475
rect 1869 96441 1903 96475
rect 1903 96441 1912 96475
rect 1860 96432 1912 96441
rect 18052 96475 18104 96484
rect 18052 96441 18061 96475
rect 18061 96441 18095 96475
rect 18095 96441 18104 96475
rect 18052 96432 18104 96441
rect 36820 96432 36872 96484
rect 16580 96364 16632 96416
rect 28908 96364 28960 96416
rect 19606 96262 19658 96314
rect 19670 96262 19722 96314
rect 19734 96262 19786 96314
rect 19798 96262 19850 96314
rect 37188 96067 37240 96076
rect 37188 96033 37197 96067
rect 37197 96033 37231 96067
rect 37231 96033 37240 96067
rect 37188 96024 37240 96033
rect 4068 95888 4120 95940
rect 28448 95888 28500 95940
rect 1952 95820 2004 95872
rect 27068 95820 27120 95872
rect 36176 95820 36228 95872
rect 4246 95718 4298 95770
rect 4310 95718 4362 95770
rect 4374 95718 4426 95770
rect 4438 95718 4490 95770
rect 34966 95718 35018 95770
rect 35030 95718 35082 95770
rect 35094 95718 35146 95770
rect 35158 95718 35210 95770
rect 1952 95659 2004 95668
rect 1952 95625 1961 95659
rect 1961 95625 1995 95659
rect 1995 95625 2004 95659
rect 1952 95616 2004 95625
rect 35992 95548 36044 95600
rect 19340 95480 19392 95532
rect 1860 95455 1912 95464
rect 1860 95421 1869 95455
rect 1869 95421 1903 95455
rect 1903 95421 1912 95455
rect 1860 95412 1912 95421
rect 15108 95412 15160 95464
rect 37280 95455 37332 95464
rect 19984 95344 20036 95396
rect 20628 95344 20680 95396
rect 37280 95421 37289 95455
rect 37289 95421 37323 95455
rect 37323 95421 37332 95455
rect 37280 95412 37332 95421
rect 37924 95455 37976 95464
rect 37924 95421 37933 95455
rect 37933 95421 37967 95455
rect 37967 95421 37976 95455
rect 37924 95412 37976 95421
rect 23940 95319 23992 95328
rect 23940 95285 23949 95319
rect 23949 95285 23983 95319
rect 23983 95285 23992 95319
rect 23940 95276 23992 95285
rect 30932 95276 30984 95328
rect 19606 95174 19658 95226
rect 19670 95174 19722 95226
rect 19734 95174 19786 95226
rect 19798 95174 19850 95226
rect 1860 94979 1912 94988
rect 1860 94945 1869 94979
rect 1869 94945 1903 94979
rect 1903 94945 1912 94979
rect 1860 94936 1912 94945
rect 37188 94979 37240 94988
rect 37188 94945 37197 94979
rect 37197 94945 37231 94979
rect 37231 94945 37240 94979
rect 37188 94936 37240 94945
rect 25504 94732 25556 94784
rect 28264 94732 28316 94784
rect 37648 94732 37700 94784
rect 38660 94732 38712 94784
rect 4246 94630 4298 94682
rect 4310 94630 4362 94682
rect 4374 94630 4426 94682
rect 4438 94630 4490 94682
rect 34966 94630 35018 94682
rect 35030 94630 35082 94682
rect 35094 94630 35146 94682
rect 35158 94630 35210 94682
rect 32772 94528 32824 94580
rect 33048 94528 33100 94580
rect 38384 94528 38436 94580
rect 38844 94528 38896 94580
rect 35900 94460 35952 94512
rect 37556 94392 37608 94444
rect 38568 94392 38620 94444
rect 37280 94367 37332 94376
rect 37280 94333 37289 94367
rect 37289 94333 37323 94367
rect 37323 94333 37332 94367
rect 37280 94324 37332 94333
rect 37924 94367 37976 94376
rect 37924 94333 37933 94367
rect 37933 94333 37967 94367
rect 37967 94333 37976 94367
rect 37924 94324 37976 94333
rect 37464 94231 37516 94240
rect 37464 94197 37473 94231
rect 37473 94197 37507 94231
rect 37507 94197 37516 94231
rect 37464 94188 37516 94197
rect 19606 94086 19658 94138
rect 19670 94086 19722 94138
rect 19734 94086 19786 94138
rect 19798 94086 19850 94138
rect 1860 93891 1912 93900
rect 1860 93857 1869 93891
rect 1869 93857 1903 93891
rect 1903 93857 1912 93891
rect 1860 93848 1912 93857
rect 26976 93848 27028 93900
rect 4246 93542 4298 93594
rect 4310 93542 4362 93594
rect 4374 93542 4426 93594
rect 4438 93542 4490 93594
rect 34966 93542 35018 93594
rect 35030 93542 35082 93594
rect 35094 93542 35146 93594
rect 35158 93542 35210 93594
rect 2044 93236 2096 93288
rect 27344 93236 27396 93288
rect 37280 93279 37332 93288
rect 37280 93245 37289 93279
rect 37289 93245 37323 93279
rect 37323 93245 37332 93279
rect 37280 93236 37332 93245
rect 1860 93211 1912 93220
rect 1860 93177 1869 93211
rect 1869 93177 1903 93211
rect 1903 93177 1912 93211
rect 1860 93168 1912 93177
rect 24860 93100 24912 93152
rect 37648 93100 37700 93152
rect 38384 93100 38436 93152
rect 19606 92998 19658 93050
rect 19670 92998 19722 93050
rect 19734 92998 19786 93050
rect 19798 92998 19850 93050
rect 37188 92803 37240 92812
rect 37188 92769 37197 92803
rect 37197 92769 37231 92803
rect 37231 92769 37240 92803
rect 37188 92760 37240 92769
rect 37372 92599 37424 92608
rect 37372 92565 37381 92599
rect 37381 92565 37415 92599
rect 37415 92565 37424 92599
rect 37372 92556 37424 92565
rect 38936 92531 38988 92540
rect 4246 92454 4298 92506
rect 4310 92454 4362 92506
rect 4374 92454 4426 92506
rect 4438 92454 4490 92506
rect 34966 92454 35018 92506
rect 35030 92454 35082 92506
rect 35094 92454 35146 92506
rect 35158 92454 35210 92506
rect 38936 92497 38945 92531
rect 38945 92497 38979 92531
rect 38979 92497 38988 92531
rect 38936 92488 38988 92497
rect 19984 92352 20036 92404
rect 35808 92284 35860 92336
rect 1860 92191 1912 92200
rect 1860 92157 1869 92191
rect 1869 92157 1903 92191
rect 1903 92157 1912 92191
rect 1860 92148 1912 92157
rect 29184 92148 29236 92200
rect 37280 92191 37332 92200
rect 37280 92157 37289 92191
rect 37289 92157 37323 92191
rect 37323 92157 37332 92191
rect 37280 92148 37332 92157
rect 37924 92191 37976 92200
rect 37924 92157 37933 92191
rect 37933 92157 37967 92191
rect 37967 92157 37976 92191
rect 37924 92148 37976 92157
rect 20076 92123 20128 92132
rect 20076 92089 20085 92123
rect 20085 92089 20119 92123
rect 20119 92089 20128 92123
rect 20076 92080 20128 92089
rect 30288 92012 30340 92064
rect 19606 91910 19658 91962
rect 19670 91910 19722 91962
rect 19734 91910 19786 91962
rect 19798 91910 19850 91962
rect 10876 91851 10928 91860
rect 10876 91817 10885 91851
rect 10885 91817 10919 91851
rect 10919 91817 10928 91851
rect 10876 91808 10928 91817
rect 15844 91851 15896 91860
rect 15844 91817 15853 91851
rect 15853 91817 15887 91851
rect 15887 91817 15896 91851
rect 15844 91808 15896 91817
rect 16028 91808 16080 91860
rect 23388 91808 23440 91860
rect 19064 91740 19116 91792
rect 26884 91740 26936 91792
rect 1860 91715 1912 91724
rect 1860 91681 1869 91715
rect 1869 91681 1903 91715
rect 1903 91681 1912 91715
rect 1860 91672 1912 91681
rect 10784 91715 10836 91724
rect 10784 91681 10793 91715
rect 10793 91681 10827 91715
rect 10827 91681 10836 91715
rect 10784 91672 10836 91681
rect 16488 91672 16540 91724
rect 1952 91511 2004 91520
rect 1952 91477 1961 91511
rect 1961 91477 1995 91511
rect 1995 91477 2004 91511
rect 1952 91468 2004 91477
rect 4246 91366 4298 91418
rect 4310 91366 4362 91418
rect 4374 91366 4426 91418
rect 4438 91366 4490 91418
rect 34966 91366 35018 91418
rect 35030 91366 35082 91418
rect 35094 91366 35146 91418
rect 35158 91366 35210 91418
rect 1952 91264 2004 91316
rect 25044 91264 25096 91316
rect 29644 91264 29696 91316
rect 28356 91103 28408 91112
rect 28356 91069 28365 91103
rect 28365 91069 28399 91103
rect 28399 91069 28408 91103
rect 28356 91060 28408 91069
rect 28448 91103 28500 91112
rect 28448 91069 28458 91103
rect 28458 91069 28492 91103
rect 28492 91069 28500 91103
rect 28632 91103 28684 91112
rect 28448 91060 28500 91069
rect 28632 91069 28641 91103
rect 28641 91069 28675 91103
rect 28675 91069 28684 91103
rect 28632 91060 28684 91069
rect 32864 91128 32916 91180
rect 37556 91196 37608 91248
rect 28724 91035 28776 91044
rect 28724 91001 28733 91035
rect 28733 91001 28767 91035
rect 28767 91001 28776 91035
rect 28724 90992 28776 91001
rect 31944 91035 31996 91044
rect 31944 91001 31953 91035
rect 31953 91001 31987 91035
rect 31987 91001 31996 91035
rect 31944 90992 31996 91001
rect 32772 91060 32824 91112
rect 37280 91103 37332 91112
rect 37280 91069 37289 91103
rect 37289 91069 37323 91103
rect 37323 91069 37332 91103
rect 37280 91060 37332 91069
rect 37464 91060 37516 91112
rect 37924 91103 37976 91112
rect 37924 91069 37933 91103
rect 37933 91069 37967 91103
rect 37967 91069 37976 91103
rect 37924 91060 37976 91069
rect 32956 90924 33008 90976
rect 19606 90822 19658 90874
rect 19670 90822 19722 90874
rect 19734 90822 19786 90874
rect 19798 90822 19850 90874
rect 13176 90720 13228 90772
rect 27344 90652 27396 90704
rect 28632 90695 28684 90704
rect 1860 90627 1912 90636
rect 1860 90593 1869 90627
rect 1869 90593 1903 90627
rect 1903 90593 1912 90627
rect 1860 90584 1912 90593
rect 19892 90584 19944 90636
rect 26792 90584 26844 90636
rect 28632 90661 28641 90695
rect 28641 90661 28675 90695
rect 28675 90661 28684 90695
rect 28632 90652 28684 90661
rect 28724 90627 28776 90636
rect 28724 90593 28733 90627
rect 28733 90593 28767 90627
rect 28767 90593 28776 90627
rect 28724 90584 28776 90593
rect 35992 90652 36044 90704
rect 29092 90516 29144 90568
rect 31852 90584 31904 90636
rect 32312 90584 32364 90636
rect 32864 90584 32916 90636
rect 33232 90584 33284 90636
rect 37188 90627 37240 90636
rect 37188 90593 37197 90627
rect 37197 90593 37231 90627
rect 37231 90593 37240 90627
rect 37188 90584 37240 90593
rect 31392 90448 31444 90500
rect 1952 90423 2004 90432
rect 1952 90389 1961 90423
rect 1961 90389 1995 90423
rect 1995 90389 2004 90423
rect 1952 90380 2004 90389
rect 29000 90423 29052 90432
rect 29000 90389 29009 90423
rect 29009 90389 29043 90423
rect 29043 90389 29052 90423
rect 29000 90380 29052 90389
rect 30564 90380 30616 90432
rect 32864 90380 32916 90432
rect 38016 90380 38068 90432
rect 4246 90278 4298 90330
rect 4310 90278 4362 90330
rect 4374 90278 4426 90330
rect 4438 90278 4490 90330
rect 34966 90278 35018 90330
rect 35030 90278 35082 90330
rect 35094 90278 35146 90330
rect 35158 90278 35210 90330
rect 1952 90176 2004 90228
rect 24124 90176 24176 90228
rect 17316 90040 17368 90092
rect 16488 89972 16540 90024
rect 27804 89972 27856 90024
rect 28632 90015 28684 90024
rect 19340 89904 19392 89956
rect 28632 89981 28641 90015
rect 28641 89981 28675 90015
rect 28675 89981 28684 90015
rect 28632 89972 28684 89981
rect 35900 90176 35952 90228
rect 33048 90108 33100 90160
rect 33324 90108 33376 90160
rect 32772 90083 32824 90092
rect 32772 90049 32781 90083
rect 32781 90049 32815 90083
rect 32815 90049 32824 90083
rect 32772 90040 32824 90049
rect 29000 89972 29052 90024
rect 32956 89972 33008 90024
rect 37280 90015 37332 90024
rect 37280 89981 37289 90015
rect 37289 89981 37323 90015
rect 37323 89981 37332 90015
rect 37280 89972 37332 89981
rect 37924 90015 37976 90024
rect 37924 89981 37933 90015
rect 37933 89981 37967 90015
rect 37967 89981 37976 90015
rect 37924 89972 37976 89981
rect 28724 89947 28776 89956
rect 28724 89913 28733 89947
rect 28733 89913 28767 89947
rect 28767 89913 28776 89947
rect 28724 89904 28776 89913
rect 32220 89904 32272 89956
rect 28448 89836 28500 89888
rect 32588 89836 32640 89888
rect 37464 89879 37516 89888
rect 37464 89845 37473 89879
rect 37473 89845 37507 89879
rect 37507 89845 37516 89879
rect 37464 89836 37516 89845
rect 19606 89734 19658 89786
rect 19670 89734 19722 89786
rect 19734 89734 19786 89786
rect 19798 89734 19850 89786
rect 29092 89632 29144 89684
rect 32312 89632 32364 89684
rect 32772 89632 32824 89684
rect 33324 89632 33376 89684
rect 33692 89632 33744 89684
rect 1860 89607 1912 89616
rect 1860 89573 1869 89607
rect 1869 89573 1903 89607
rect 1903 89573 1912 89607
rect 1860 89564 1912 89573
rect 6276 89496 6328 89548
rect 27712 89496 27764 89548
rect 28448 89496 28500 89548
rect 28632 89539 28684 89548
rect 28632 89505 28641 89539
rect 28641 89505 28675 89539
rect 28675 89505 28684 89539
rect 28632 89496 28684 89505
rect 28816 89496 28868 89548
rect 28908 89496 28960 89548
rect 31852 89496 31904 89548
rect 38476 89564 38528 89616
rect 31484 89471 31536 89480
rect 31484 89437 31493 89471
rect 31493 89437 31527 89471
rect 31527 89437 31536 89471
rect 31484 89428 31536 89437
rect 32772 89428 32824 89480
rect 3424 89360 3476 89412
rect 29828 89360 29880 89412
rect 33968 89496 34020 89548
rect 34152 89539 34204 89548
rect 34152 89505 34161 89539
rect 34161 89505 34195 89539
rect 34195 89505 34204 89539
rect 34152 89496 34204 89505
rect 36360 89428 36412 89480
rect 36636 89428 36688 89480
rect 30380 89292 30432 89344
rect 31852 89292 31904 89344
rect 32956 89292 33008 89344
rect 33324 89292 33376 89344
rect 36636 89292 36688 89344
rect 37188 89292 37240 89344
rect 4246 89190 4298 89242
rect 4310 89190 4362 89242
rect 4374 89190 4426 89242
rect 4438 89190 4490 89242
rect 34966 89190 35018 89242
rect 35030 89190 35082 89242
rect 35094 89190 35146 89242
rect 35158 89190 35210 89242
rect 28908 89131 28960 89140
rect 28908 89097 28917 89131
rect 28917 89097 28951 89131
rect 28951 89097 28960 89131
rect 28908 89088 28960 89097
rect 29000 89088 29052 89140
rect 38384 89088 38436 89140
rect 28816 89020 28868 89072
rect 31484 89020 31536 89072
rect 32772 89020 32824 89072
rect 37648 89020 37700 89072
rect 3516 88884 3568 88936
rect 23388 88884 23440 88936
rect 27896 88884 27948 88936
rect 38568 88952 38620 89004
rect 32588 88927 32640 88936
rect 1860 88859 1912 88868
rect 1860 88825 1869 88859
rect 1869 88825 1903 88859
rect 1903 88825 1912 88859
rect 1860 88816 1912 88825
rect 9220 88816 9272 88868
rect 27160 88816 27212 88868
rect 27804 88816 27856 88868
rect 28448 88816 28500 88868
rect 28632 88859 28684 88868
rect 28632 88825 28641 88859
rect 28641 88825 28675 88859
rect 28675 88825 28684 88859
rect 28632 88816 28684 88825
rect 29368 88816 29420 88868
rect 31300 88816 31352 88868
rect 31852 88816 31904 88868
rect 32588 88893 32597 88927
rect 32597 88893 32631 88927
rect 32631 88893 32640 88927
rect 32588 88884 32640 88893
rect 32772 88884 32824 88936
rect 32956 88927 33008 88936
rect 32956 88893 32965 88927
rect 32965 88893 32999 88927
rect 32999 88893 33008 88927
rect 32956 88884 33008 88893
rect 37280 88927 37332 88936
rect 37280 88893 37289 88927
rect 37289 88893 37323 88927
rect 37323 88893 37332 88927
rect 37280 88884 37332 88893
rect 37924 88927 37976 88936
rect 37924 88893 37933 88927
rect 37933 88893 37967 88927
rect 37967 88893 37976 88927
rect 37924 88884 37976 88893
rect 38108 88884 38160 88936
rect 38384 88884 38436 88936
rect 37372 88816 37424 88868
rect 30748 88748 30800 88800
rect 35808 88748 35860 88800
rect 36084 88748 36136 88800
rect 38108 88791 38160 88800
rect 38108 88757 38117 88791
rect 38117 88757 38151 88791
rect 38151 88757 38160 88791
rect 38108 88748 38160 88757
rect 19606 88646 19658 88698
rect 19670 88646 19722 88698
rect 19734 88646 19786 88698
rect 19798 88646 19850 88698
rect 9128 88544 9180 88596
rect 28172 88544 28224 88596
rect 31668 88544 31720 88596
rect 32312 88544 32364 88596
rect 32772 88544 32824 88596
rect 33048 88544 33100 88596
rect 16580 88476 16632 88528
rect 28816 88476 28868 88528
rect 29000 88476 29052 88528
rect 27436 88408 27488 88460
rect 28172 88451 28224 88460
rect 28172 88417 28182 88451
rect 28182 88417 28216 88451
rect 28216 88417 28224 88451
rect 28172 88408 28224 88417
rect 27252 88272 27304 88324
rect 28448 88451 28500 88460
rect 28448 88417 28457 88451
rect 28457 88417 28491 88451
rect 28491 88417 28500 88451
rect 28448 88408 28500 88417
rect 28908 88408 28960 88460
rect 29092 88408 29144 88460
rect 28816 88340 28868 88392
rect 30748 88408 30800 88460
rect 31392 88408 31444 88460
rect 27620 88204 27672 88256
rect 28448 88204 28500 88256
rect 29828 88340 29880 88392
rect 30840 88340 30892 88392
rect 31208 88340 31260 88392
rect 31484 88383 31536 88392
rect 31484 88349 31493 88383
rect 31493 88349 31527 88383
rect 31527 88349 31536 88383
rect 31484 88340 31536 88349
rect 32404 88408 32456 88460
rect 32588 88408 32640 88460
rect 33232 88408 33284 88460
rect 35808 88476 35860 88528
rect 38108 88476 38160 88528
rect 31024 88272 31076 88324
rect 32312 88340 32364 88392
rect 32404 88272 32456 88324
rect 33968 88408 34020 88460
rect 34244 88451 34296 88460
rect 34244 88417 34253 88451
rect 34253 88417 34287 88451
rect 34287 88417 34296 88451
rect 34244 88408 34296 88417
rect 37188 88451 37240 88460
rect 37188 88417 37197 88451
rect 37197 88417 37231 88451
rect 37231 88417 37240 88451
rect 37188 88408 37240 88417
rect 33232 88204 33284 88256
rect 4246 88102 4298 88154
rect 4310 88102 4362 88154
rect 4374 88102 4426 88154
rect 4438 88102 4490 88154
rect 34966 88102 35018 88154
rect 35030 88102 35082 88154
rect 35094 88102 35146 88154
rect 35158 88102 35210 88154
rect 24124 88000 24176 88052
rect 28172 87932 28224 87984
rect 11704 87864 11756 87916
rect 29000 88000 29052 88052
rect 28816 87932 28868 87984
rect 1860 87839 1912 87848
rect 1860 87805 1869 87839
rect 1869 87805 1903 87839
rect 1903 87805 1912 87839
rect 1860 87796 1912 87805
rect 26240 87796 26292 87848
rect 27068 87839 27120 87848
rect 27068 87805 27078 87839
rect 27078 87805 27112 87839
rect 27112 87805 27120 87839
rect 27068 87796 27120 87805
rect 27528 87796 27580 87848
rect 28080 87839 28132 87848
rect 28080 87805 28089 87839
rect 28089 87805 28123 87839
rect 28123 87805 28132 87839
rect 28080 87796 28132 87805
rect 29000 87864 29052 87916
rect 30656 87932 30708 87984
rect 32404 87932 32456 87984
rect 32496 87932 32548 87984
rect 36176 87932 36228 87984
rect 31484 87864 31536 87916
rect 30288 87796 30340 87848
rect 3516 87728 3568 87780
rect 27252 87771 27304 87780
rect 27252 87737 27261 87771
rect 27261 87737 27295 87771
rect 27295 87737 27304 87771
rect 27252 87728 27304 87737
rect 27620 87728 27672 87780
rect 28448 87771 28500 87780
rect 28448 87737 28457 87771
rect 28457 87737 28491 87771
rect 28491 87737 28500 87771
rect 28448 87728 28500 87737
rect 28816 87728 28868 87780
rect 31300 87728 31352 87780
rect 31668 87796 31720 87848
rect 32312 87796 32364 87848
rect 33968 87796 34020 87848
rect 34152 87796 34204 87848
rect 35900 87796 35952 87848
rect 37280 87839 37332 87848
rect 37280 87805 37289 87839
rect 37289 87805 37323 87839
rect 37323 87805 37332 87839
rect 37280 87796 37332 87805
rect 37924 87839 37976 87848
rect 37924 87805 37933 87839
rect 37933 87805 37967 87839
rect 37967 87805 37976 87839
rect 37924 87796 37976 87805
rect 32588 87728 32640 87780
rect 28172 87660 28224 87712
rect 32404 87660 32456 87712
rect 32496 87660 32548 87712
rect 35900 87660 35952 87712
rect 19606 87558 19658 87610
rect 19670 87558 19722 87610
rect 19734 87558 19786 87610
rect 19798 87558 19850 87610
rect 26148 87456 26200 87508
rect 9036 87388 9088 87440
rect 1860 87363 1912 87372
rect 1860 87329 1869 87363
rect 1869 87329 1903 87363
rect 1903 87329 1912 87363
rect 1860 87320 1912 87329
rect 23388 87363 23440 87372
rect 23388 87329 23397 87363
rect 23397 87329 23431 87363
rect 23431 87329 23440 87363
rect 23388 87320 23440 87329
rect 27344 87320 27396 87372
rect 28172 87388 28224 87440
rect 31208 87456 31260 87508
rect 32956 87456 33008 87508
rect 33968 87456 34020 87508
rect 37004 87456 37056 87508
rect 30932 87388 30984 87440
rect 32404 87388 32456 87440
rect 37556 87388 37608 87440
rect 29552 87320 29604 87372
rect 28908 87252 28960 87304
rect 30104 87252 30156 87304
rect 30840 87320 30892 87372
rect 28724 87184 28776 87236
rect 30748 87252 30800 87304
rect 32312 87320 32364 87372
rect 32496 87320 32548 87372
rect 32956 87320 33008 87372
rect 34612 87320 34664 87372
rect 35256 87320 35308 87372
rect 35440 87320 35492 87372
rect 31024 87252 31076 87304
rect 33968 87252 34020 87304
rect 1952 87159 2004 87168
rect 1952 87125 1961 87159
rect 1961 87125 1995 87159
rect 1995 87125 2004 87159
rect 1952 87116 2004 87125
rect 28264 87116 28316 87168
rect 28540 87116 28592 87168
rect 29276 87116 29328 87168
rect 30748 87116 30800 87168
rect 30840 87116 30892 87168
rect 34612 87184 34664 87236
rect 35164 87184 35216 87236
rect 32404 87116 32456 87168
rect 32864 87116 32916 87168
rect 35256 87116 35308 87168
rect 4246 87014 4298 87066
rect 4310 87014 4362 87066
rect 4374 87014 4426 87066
rect 4438 87014 4490 87066
rect 34966 87014 35018 87066
rect 35030 87014 35082 87066
rect 35094 87014 35146 87066
rect 35158 87014 35210 87066
rect 4804 86912 4856 86964
rect 27620 86912 27672 86964
rect 20076 86776 20128 86828
rect 19340 86708 19392 86760
rect 24860 86776 24912 86828
rect 23388 86708 23440 86760
rect 26608 86708 26660 86760
rect 27160 86751 27212 86760
rect 27160 86717 27169 86751
rect 27169 86717 27203 86751
rect 27203 86717 27212 86751
rect 27160 86708 27212 86717
rect 27528 86776 27580 86828
rect 32496 86912 32548 86964
rect 32588 86912 32640 86964
rect 28172 86844 28224 86896
rect 28264 86776 28316 86828
rect 30104 86844 30156 86896
rect 31024 86844 31076 86896
rect 19432 86640 19484 86692
rect 20168 86640 20220 86692
rect 22744 86640 22796 86692
rect 18236 86572 18288 86624
rect 19340 86572 19392 86624
rect 26700 86640 26752 86692
rect 28540 86708 28592 86760
rect 28908 86776 28960 86828
rect 31668 86844 31720 86896
rect 32772 86844 32824 86896
rect 32956 86844 33008 86896
rect 32128 86819 32180 86828
rect 32128 86785 32137 86819
rect 32137 86785 32171 86819
rect 32171 86785 32180 86819
rect 32128 86776 32180 86785
rect 28908 86640 28960 86692
rect 29828 86708 29880 86760
rect 32404 86708 32456 86760
rect 30288 86640 30340 86692
rect 30932 86640 30984 86692
rect 31208 86640 31260 86692
rect 32772 86708 32824 86760
rect 32588 86640 32640 86692
rect 33968 86912 34020 86964
rect 37464 86912 37516 86964
rect 33968 86708 34020 86760
rect 37280 86751 37332 86760
rect 37280 86717 37289 86751
rect 37289 86717 37323 86751
rect 37323 86717 37332 86751
rect 37280 86708 37332 86717
rect 37924 86751 37976 86760
rect 37924 86717 37933 86751
rect 37933 86717 37967 86751
rect 37967 86717 37976 86751
rect 37924 86708 37976 86717
rect 28540 86572 28592 86624
rect 32404 86572 32456 86624
rect 32772 86615 32824 86624
rect 32772 86581 32781 86615
rect 32781 86581 32815 86615
rect 32815 86581 32824 86615
rect 32772 86572 32824 86581
rect 34244 86572 34296 86624
rect 37556 86572 37608 86624
rect 37648 86572 37700 86624
rect 19606 86470 19658 86522
rect 19670 86470 19722 86522
rect 19734 86470 19786 86522
rect 19798 86470 19850 86522
rect 20076 86368 20128 86420
rect 27804 86368 27856 86420
rect 29276 86368 29328 86420
rect 29828 86368 29880 86420
rect 32312 86368 32364 86420
rect 1860 86343 1912 86352
rect 1860 86309 1869 86343
rect 1869 86309 1903 86343
rect 1903 86309 1912 86343
rect 1860 86300 1912 86309
rect 25504 86300 25556 86352
rect 19892 86275 19944 86284
rect 19892 86241 19901 86275
rect 19901 86241 19935 86275
rect 19935 86241 19944 86275
rect 19892 86232 19944 86241
rect 23388 86275 23440 86284
rect 23388 86241 23397 86275
rect 23397 86241 23431 86275
rect 23431 86241 23440 86275
rect 23388 86232 23440 86241
rect 26700 86275 26752 86284
rect 26700 86241 26709 86275
rect 26709 86241 26743 86275
rect 26743 86241 26752 86275
rect 26700 86232 26752 86241
rect 28816 86300 28868 86352
rect 26332 86164 26384 86216
rect 27252 86164 27304 86216
rect 2044 86139 2096 86148
rect 2044 86105 2053 86139
rect 2053 86105 2087 86139
rect 2087 86105 2096 86139
rect 2044 86096 2096 86105
rect 28264 86096 28316 86148
rect 28816 86164 28868 86216
rect 23296 86028 23348 86080
rect 26976 86028 27028 86080
rect 29277 86232 29329 86284
rect 29644 86232 29696 86284
rect 30748 86300 30800 86352
rect 35992 86300 36044 86352
rect 29828 86164 29880 86216
rect 30012 86164 30064 86216
rect 30288 86232 30340 86284
rect 32128 86232 32180 86284
rect 32496 86232 32548 86284
rect 32864 86232 32916 86284
rect 37188 86275 37240 86284
rect 37188 86241 37197 86275
rect 37197 86241 37231 86275
rect 37231 86241 37240 86275
rect 37188 86232 37240 86241
rect 37096 86164 37148 86216
rect 29276 86096 29328 86148
rect 31484 86096 31536 86148
rect 31668 86096 31720 86148
rect 31024 86071 31076 86080
rect 31024 86037 31033 86071
rect 31033 86037 31067 86071
rect 31067 86037 31076 86071
rect 31024 86028 31076 86037
rect 31208 86028 31260 86080
rect 33692 86028 33744 86080
rect 37372 86071 37424 86080
rect 37372 86037 37381 86071
rect 37381 86037 37415 86071
rect 37415 86037 37424 86071
rect 37372 86028 37424 86037
rect 4246 85926 4298 85978
rect 4310 85926 4362 85978
rect 4374 85926 4426 85978
rect 4438 85926 4490 85978
rect 34966 85926 35018 85978
rect 35030 85926 35082 85978
rect 35094 85926 35146 85978
rect 35158 85926 35210 85978
rect 1860 85663 1912 85672
rect 1860 85629 1869 85663
rect 1869 85629 1903 85663
rect 1903 85629 1912 85663
rect 1860 85620 1912 85629
rect 21824 85620 21876 85672
rect 28540 85824 28592 85876
rect 28816 85824 28868 85876
rect 29644 85824 29696 85876
rect 30748 85756 30800 85808
rect 29184 85688 29236 85740
rect 2688 85552 2740 85604
rect 10324 85552 10376 85604
rect 27804 85484 27856 85536
rect 28540 85620 28592 85672
rect 29828 85688 29880 85740
rect 28172 85595 28224 85604
rect 28172 85561 28181 85595
rect 28181 85561 28215 85595
rect 28215 85561 28224 85595
rect 28172 85552 28224 85561
rect 28816 85552 28868 85604
rect 28908 85484 28960 85536
rect 31208 85620 31260 85672
rect 30748 85595 30800 85604
rect 30748 85561 30757 85595
rect 30757 85561 30791 85595
rect 30791 85561 30800 85595
rect 30748 85552 30800 85561
rect 29368 85484 29420 85536
rect 29552 85527 29604 85536
rect 29552 85493 29561 85527
rect 29561 85493 29595 85527
rect 29595 85493 29604 85527
rect 29552 85484 29604 85493
rect 30380 85484 30432 85536
rect 31484 85663 31536 85672
rect 31484 85629 31493 85663
rect 31493 85629 31527 85663
rect 31527 85629 31536 85663
rect 32128 85688 32180 85740
rect 31484 85620 31536 85629
rect 34152 85756 34204 85808
rect 36912 85756 36964 85808
rect 32404 85688 32456 85740
rect 32680 85663 32732 85672
rect 32680 85629 32689 85663
rect 32689 85629 32723 85663
rect 32723 85629 32732 85663
rect 32680 85620 32732 85629
rect 32956 85663 33008 85672
rect 32588 85552 32640 85604
rect 32956 85629 32965 85663
rect 32965 85629 32999 85663
rect 32999 85629 33008 85663
rect 32956 85620 33008 85629
rect 33968 85620 34020 85672
rect 37280 85663 37332 85672
rect 37280 85629 37289 85663
rect 37289 85629 37323 85663
rect 37323 85629 37332 85663
rect 37280 85620 37332 85629
rect 37924 85663 37976 85672
rect 37924 85629 37933 85663
rect 37933 85629 37967 85663
rect 37967 85629 37976 85663
rect 37924 85620 37976 85629
rect 32496 85527 32548 85536
rect 32496 85493 32505 85527
rect 32505 85493 32539 85527
rect 32539 85493 32548 85527
rect 32496 85484 32548 85493
rect 33876 85484 33928 85536
rect 19606 85382 19658 85434
rect 19670 85382 19722 85434
rect 19734 85382 19786 85434
rect 19798 85382 19850 85434
rect 27252 85280 27304 85332
rect 27804 85280 27856 85332
rect 8944 85212 8996 85264
rect 28356 85280 28408 85332
rect 28816 85280 28868 85332
rect 28908 85280 28960 85332
rect 23388 85144 23440 85196
rect 26424 85144 26476 85196
rect 26700 85187 26752 85196
rect 26700 85153 26709 85187
rect 26709 85153 26743 85187
rect 26743 85153 26752 85187
rect 26700 85144 26752 85153
rect 27160 85144 27212 85196
rect 23296 85076 23348 85128
rect 29276 85280 29328 85332
rect 32956 85280 33008 85332
rect 33416 85280 33468 85332
rect 28172 85187 28224 85196
rect 28172 85153 28181 85187
rect 28181 85153 28215 85187
rect 28215 85153 28224 85187
rect 28172 85144 28224 85153
rect 28448 85144 28500 85196
rect 25872 85008 25924 85060
rect 28356 85008 28408 85060
rect 28172 84940 28224 84992
rect 28908 85187 28960 85196
rect 28908 85153 28917 85187
rect 28917 85153 28951 85187
rect 28951 85153 28960 85187
rect 28908 85144 28960 85153
rect 29000 85187 29052 85196
rect 29000 85153 29010 85187
rect 29010 85153 29044 85187
rect 29044 85153 29052 85187
rect 33048 85212 33100 85264
rect 29000 85144 29052 85153
rect 30104 85144 30156 85196
rect 32128 85144 32180 85196
rect 33416 85187 33468 85196
rect 33416 85153 33425 85187
rect 33425 85153 33459 85187
rect 33459 85153 33468 85187
rect 33416 85144 33468 85153
rect 29368 85008 29420 85060
rect 31484 85119 31536 85128
rect 31484 85085 31493 85119
rect 31493 85085 31527 85119
rect 31527 85085 31536 85119
rect 31484 85076 31536 85085
rect 36636 85076 36688 85128
rect 29828 85008 29880 85060
rect 31208 85008 31260 85060
rect 32956 84940 33008 84992
rect 4246 84838 4298 84890
rect 4310 84838 4362 84890
rect 4374 84838 4426 84890
rect 4438 84838 4490 84890
rect 34966 84838 35018 84890
rect 35030 84838 35082 84890
rect 35094 84838 35146 84890
rect 35158 84838 35210 84890
rect 27528 84668 27580 84720
rect 25044 84600 25096 84652
rect 1860 84575 1912 84584
rect 1860 84541 1869 84575
rect 1869 84541 1903 84575
rect 1903 84541 1912 84575
rect 1860 84532 1912 84541
rect 27068 84532 27120 84584
rect 36084 84736 36136 84788
rect 37740 84736 37792 84788
rect 38200 84736 38252 84788
rect 28632 84668 28684 84720
rect 30656 84668 30708 84720
rect 31484 84668 31536 84720
rect 28448 84600 28500 84652
rect 29828 84600 29880 84652
rect 30472 84600 30524 84652
rect 28632 84532 28684 84584
rect 29644 84532 29696 84584
rect 31208 84575 31260 84584
rect 31208 84541 31217 84575
rect 31217 84541 31251 84575
rect 31251 84541 31260 84575
rect 31484 84575 31536 84584
rect 31208 84532 31260 84541
rect 31484 84541 31493 84575
rect 31493 84541 31527 84575
rect 31527 84541 31536 84575
rect 31484 84532 31536 84541
rect 2596 84464 2648 84516
rect 29276 84464 29328 84516
rect 29828 84464 29880 84516
rect 29000 84396 29052 84448
rect 30472 84507 30524 84516
rect 30472 84473 30481 84507
rect 30481 84473 30515 84507
rect 30515 84473 30524 84507
rect 33968 84668 34020 84720
rect 30472 84464 30524 84473
rect 32312 84464 32364 84516
rect 36728 84532 36780 84584
rect 37280 84575 37332 84584
rect 37280 84541 37289 84575
rect 37289 84541 37323 84575
rect 37323 84541 37332 84575
rect 37280 84532 37332 84541
rect 37924 84575 37976 84584
rect 37924 84541 37933 84575
rect 37933 84541 37967 84575
rect 37967 84541 37976 84575
rect 37924 84532 37976 84541
rect 34244 84464 34296 84516
rect 38660 84464 38712 84516
rect 37740 84396 37792 84448
rect 19606 84294 19658 84346
rect 19670 84294 19722 84346
rect 19734 84294 19786 84346
rect 19798 84294 19850 84346
rect 9220 84124 9272 84176
rect 1860 84099 1912 84108
rect 1860 84065 1869 84099
rect 1869 84065 1903 84099
rect 1903 84065 1912 84099
rect 1860 84056 1912 84065
rect 27804 84099 27856 84108
rect 27804 84065 27813 84099
rect 27813 84065 27847 84099
rect 27847 84065 27856 84099
rect 27804 84056 27856 84065
rect 28724 84124 28776 84176
rect 29092 84124 29144 84176
rect 29368 84124 29420 84176
rect 4068 83920 4120 83972
rect 28448 84056 28500 84108
rect 28632 84056 28684 84108
rect 29092 83988 29144 84040
rect 29000 83852 29052 83904
rect 29276 84056 29328 84108
rect 30012 84056 30064 84108
rect 30380 84192 30432 84244
rect 31668 84192 31720 84244
rect 31484 84056 31536 84108
rect 36544 84056 36596 84108
rect 37188 84099 37240 84108
rect 37188 84065 37197 84099
rect 37197 84065 37231 84099
rect 37231 84065 37240 84099
rect 37188 84056 37240 84065
rect 30656 83988 30708 84040
rect 31208 83988 31260 84040
rect 33692 83988 33744 84040
rect 36360 83988 36412 84040
rect 35900 83920 35952 83972
rect 30380 83852 30432 83904
rect 31484 83852 31536 83904
rect 36360 83852 36412 83904
rect 4246 83750 4298 83802
rect 4310 83750 4362 83802
rect 4374 83750 4426 83802
rect 4438 83750 4490 83802
rect 34966 83750 35018 83802
rect 35030 83750 35082 83802
rect 35094 83750 35146 83802
rect 35158 83750 35210 83802
rect 25136 83648 25188 83700
rect 3424 83580 3476 83632
rect 30472 83648 30524 83700
rect 31668 83648 31720 83700
rect 26884 83444 26936 83496
rect 30656 83580 30708 83632
rect 31208 83580 31260 83632
rect 28172 83512 28224 83564
rect 28724 83512 28776 83564
rect 29000 83512 29052 83564
rect 29092 83376 29144 83428
rect 28632 83308 28684 83360
rect 29276 83487 29328 83496
rect 29276 83453 29285 83487
rect 29285 83453 29319 83487
rect 29319 83453 29328 83487
rect 29276 83444 29328 83453
rect 31208 83487 31260 83496
rect 31208 83453 31217 83487
rect 31217 83453 31251 83487
rect 31251 83453 31260 83487
rect 31208 83444 31260 83453
rect 34244 83444 34296 83496
rect 37280 83487 37332 83496
rect 37280 83453 37289 83487
rect 37289 83453 37323 83487
rect 37323 83453 37332 83487
rect 37280 83444 37332 83453
rect 37924 83487 37976 83496
rect 37924 83453 37933 83487
rect 37933 83453 37967 83487
rect 37967 83453 37976 83487
rect 37924 83444 37976 83453
rect 30104 83376 30156 83428
rect 37648 83376 37700 83428
rect 35808 83308 35860 83360
rect 37464 83351 37516 83360
rect 37464 83317 37473 83351
rect 37473 83317 37507 83351
rect 37507 83317 37516 83351
rect 37464 83308 37516 83317
rect 38108 83351 38160 83360
rect 38108 83317 38117 83351
rect 38117 83317 38151 83351
rect 38151 83317 38160 83351
rect 38108 83308 38160 83317
rect 19606 83206 19658 83258
rect 19670 83206 19722 83258
rect 19734 83206 19786 83258
rect 19798 83206 19850 83258
rect 27252 83104 27304 83156
rect 3516 83036 3568 83088
rect 28172 83104 28224 83156
rect 1400 83011 1452 83020
rect 1400 82977 1409 83011
rect 1409 82977 1443 83011
rect 1443 82977 1452 83011
rect 1400 82968 1452 82977
rect 26976 82968 27028 83020
rect 36176 83104 36228 83156
rect 30380 83036 30432 83088
rect 30656 83011 30708 83020
rect 8852 82900 8904 82952
rect 30656 82977 30665 83011
rect 30665 82977 30699 83011
rect 30699 82977 30708 83011
rect 30656 82968 30708 82977
rect 31116 83011 31168 83020
rect 31116 82977 31125 83011
rect 31125 82977 31159 83011
rect 31159 82977 31168 83011
rect 31116 82968 31168 82977
rect 31208 82900 31260 82952
rect 28264 82832 28316 82884
rect 29828 82832 29880 82884
rect 29092 82764 29144 82816
rect 4246 82662 4298 82714
rect 4310 82662 4362 82714
rect 4374 82662 4426 82714
rect 4438 82662 4490 82714
rect 34966 82662 35018 82714
rect 35030 82662 35082 82714
rect 35094 82662 35146 82714
rect 35158 82662 35210 82714
rect 29000 82560 29052 82612
rect 30656 82560 30708 82612
rect 2044 82492 2096 82544
rect 1952 82424 2004 82476
rect 26700 82356 26752 82408
rect 27528 82424 27580 82476
rect 28172 82356 28224 82408
rect 29828 82492 29880 82544
rect 30288 82492 30340 82544
rect 28724 82399 28776 82408
rect 28724 82365 28733 82399
rect 28733 82365 28767 82399
rect 28767 82365 28776 82399
rect 28724 82356 28776 82365
rect 37372 82492 37424 82544
rect 39212 82492 39264 82544
rect 31576 82467 31628 82476
rect 31576 82433 31585 82467
rect 31585 82433 31619 82467
rect 31619 82433 31628 82467
rect 31576 82424 31628 82433
rect 31116 82399 31168 82408
rect 31116 82365 31125 82399
rect 31125 82365 31159 82399
rect 31159 82365 31168 82399
rect 31116 82356 31168 82365
rect 31208 82399 31260 82408
rect 31208 82365 31217 82399
rect 31217 82365 31251 82399
rect 31251 82365 31260 82399
rect 31208 82356 31260 82365
rect 34152 82356 34204 82408
rect 37280 82399 37332 82408
rect 37280 82365 37289 82399
rect 37289 82365 37323 82399
rect 37323 82365 37332 82399
rect 37280 82356 37332 82365
rect 37924 82399 37976 82408
rect 37924 82365 37933 82399
rect 37933 82365 37967 82399
rect 37967 82365 37976 82399
rect 37924 82356 37976 82365
rect 1860 82331 1912 82340
rect 1860 82297 1869 82331
rect 1869 82297 1903 82331
rect 1903 82297 1912 82331
rect 1860 82288 1912 82297
rect 27252 82288 27304 82340
rect 29092 82288 29144 82340
rect 30012 82288 30064 82340
rect 30472 82331 30524 82340
rect 30472 82297 30481 82331
rect 30481 82297 30515 82331
rect 30515 82297 30524 82331
rect 30472 82288 30524 82297
rect 31576 82288 31628 82340
rect 22100 82220 22152 82272
rect 28724 82220 28776 82272
rect 37556 82288 37608 82340
rect 37280 82220 37332 82272
rect 19606 82118 19658 82170
rect 19670 82118 19722 82170
rect 19734 82118 19786 82170
rect 19798 82118 19850 82170
rect 28632 82016 28684 82068
rect 28724 81923 28776 81932
rect 28724 81889 28733 81923
rect 28733 81889 28767 81923
rect 28767 81889 28776 81923
rect 28724 81880 28776 81889
rect 28632 81855 28684 81864
rect 28632 81821 28641 81855
rect 28641 81821 28675 81855
rect 28675 81821 28684 81855
rect 28632 81812 28684 81821
rect 30288 82016 30340 82068
rect 33876 82016 33928 82068
rect 33048 81948 33100 82000
rect 29184 81923 29236 81932
rect 29184 81889 29193 81923
rect 29193 81889 29227 81923
rect 29227 81889 29236 81923
rect 29184 81880 29236 81889
rect 30656 81880 30708 81932
rect 31576 81880 31628 81932
rect 37188 81923 37240 81932
rect 37188 81889 37197 81923
rect 37197 81889 37231 81923
rect 37231 81889 37240 81923
rect 37188 81880 37240 81889
rect 23848 81744 23900 81796
rect 27252 81676 27304 81728
rect 38384 81812 38436 81864
rect 31208 81744 31260 81796
rect 32864 81676 32916 81728
rect 37556 81676 37608 81728
rect 4246 81574 4298 81626
rect 4310 81574 4362 81626
rect 4374 81574 4426 81626
rect 4438 81574 4490 81626
rect 34966 81574 35018 81626
rect 35030 81574 35082 81626
rect 35094 81574 35146 81626
rect 35158 81574 35210 81626
rect 31576 81472 31628 81524
rect 28172 81336 28224 81388
rect 29184 81336 29236 81388
rect 29460 81379 29512 81388
rect 29460 81345 29469 81379
rect 29469 81345 29503 81379
rect 29503 81345 29512 81379
rect 29460 81336 29512 81345
rect 1860 81311 1912 81320
rect 1860 81277 1869 81311
rect 1869 81277 1903 81311
rect 1903 81277 1912 81311
rect 1860 81268 1912 81277
rect 29000 81311 29052 81320
rect 29000 81277 29009 81311
rect 29009 81277 29043 81311
rect 29043 81277 29052 81311
rect 29000 81268 29052 81277
rect 2044 81243 2096 81252
rect 2044 81209 2053 81243
rect 2053 81209 2087 81243
rect 2087 81209 2096 81243
rect 2044 81200 2096 81209
rect 24584 81200 24636 81252
rect 28632 81200 28684 81252
rect 31116 81311 31168 81320
rect 31116 81277 31125 81311
rect 31125 81277 31159 81311
rect 31159 81277 31168 81311
rect 31116 81268 31168 81277
rect 31208 81311 31260 81320
rect 31208 81277 31217 81311
rect 31217 81277 31251 81311
rect 31251 81277 31260 81311
rect 38200 81336 38252 81388
rect 31208 81268 31260 81277
rect 32404 81268 32456 81320
rect 27344 81132 27396 81184
rect 27528 81132 27580 81184
rect 29460 81200 29512 81252
rect 30380 81200 30432 81252
rect 31576 81200 31628 81252
rect 32680 81200 32732 81252
rect 29644 81132 29696 81184
rect 33048 81268 33100 81320
rect 33508 81268 33560 81320
rect 37280 81311 37332 81320
rect 37280 81277 37289 81311
rect 37289 81277 37323 81311
rect 37323 81277 37332 81311
rect 37280 81268 37332 81277
rect 37924 81311 37976 81320
rect 37924 81277 37933 81311
rect 37933 81277 37967 81311
rect 37967 81277 37976 81311
rect 37924 81268 37976 81277
rect 39396 81200 39448 81252
rect 39304 81132 39356 81184
rect 19606 81030 19658 81082
rect 19670 81030 19722 81082
rect 19734 81030 19786 81082
rect 19798 81030 19850 81082
rect 2688 80860 2740 80912
rect 1400 80835 1452 80844
rect 1400 80801 1409 80835
rect 1409 80801 1443 80835
rect 1443 80801 1452 80835
rect 1400 80792 1452 80801
rect 25780 80792 25832 80844
rect 30104 80928 30156 80980
rect 31208 80928 31260 80980
rect 29460 80860 29512 80912
rect 25872 80724 25924 80776
rect 29184 80792 29236 80844
rect 31208 80792 31260 80844
rect 2688 80588 2740 80640
rect 29460 80724 29512 80776
rect 29644 80724 29696 80776
rect 30104 80767 30156 80776
rect 30104 80733 30113 80767
rect 30113 80733 30147 80767
rect 30147 80733 30156 80767
rect 30104 80724 30156 80733
rect 28632 80588 28684 80640
rect 29644 80631 29696 80640
rect 29644 80597 29653 80631
rect 29653 80597 29687 80631
rect 29687 80597 29696 80631
rect 29644 80588 29696 80597
rect 30656 80588 30708 80640
rect 32864 80792 32916 80844
rect 31944 80724 31996 80776
rect 32588 80656 32640 80708
rect 38016 80588 38068 80640
rect 4246 80486 4298 80538
rect 4310 80486 4362 80538
rect 4374 80486 4426 80538
rect 4438 80486 4490 80538
rect 34966 80486 35018 80538
rect 35030 80486 35082 80538
rect 35094 80486 35146 80538
rect 35158 80486 35210 80538
rect 28172 80384 28224 80436
rect 24124 80316 24176 80368
rect 28264 80316 28316 80368
rect 4068 80248 4120 80300
rect 2596 80180 2648 80232
rect 25688 80180 25740 80232
rect 28264 80223 28316 80232
rect 28264 80189 28273 80223
rect 28273 80189 28307 80223
rect 28307 80189 28316 80223
rect 28264 80180 28316 80189
rect 28632 80248 28684 80300
rect 29000 80248 29052 80300
rect 31116 80248 31168 80300
rect 30288 80180 30340 80232
rect 31392 80316 31444 80368
rect 31944 80384 31996 80436
rect 39028 80316 39080 80368
rect 25872 80044 25924 80096
rect 28632 80155 28684 80164
rect 28632 80121 28641 80155
rect 28641 80121 28675 80155
rect 28675 80121 28684 80155
rect 28632 80112 28684 80121
rect 29460 80112 29512 80164
rect 32956 80180 33008 80232
rect 37280 80223 37332 80232
rect 37280 80189 37289 80223
rect 37289 80189 37323 80223
rect 37323 80189 37332 80223
rect 37280 80180 37332 80189
rect 37924 80223 37976 80232
rect 37924 80189 37933 80223
rect 37933 80189 37967 80223
rect 37967 80189 37976 80223
rect 37924 80180 37976 80189
rect 28172 80044 28224 80096
rect 29276 80044 29328 80096
rect 31116 80087 31168 80096
rect 31116 80053 31125 80087
rect 31125 80053 31159 80087
rect 31159 80053 31168 80087
rect 31116 80044 31168 80053
rect 32588 80112 32640 80164
rect 36912 80112 36964 80164
rect 36728 80044 36780 80096
rect 19606 79942 19658 79994
rect 19670 79942 19722 79994
rect 19734 79942 19786 79994
rect 19798 79942 19850 79994
rect 8852 79840 8904 79892
rect 1400 79747 1452 79756
rect 1400 79713 1409 79747
rect 1409 79713 1443 79747
rect 1443 79713 1452 79747
rect 1400 79704 1452 79713
rect 2044 79636 2096 79688
rect 25596 79704 25648 79756
rect 26424 79772 26476 79824
rect 28172 79815 28224 79824
rect 28172 79781 28181 79815
rect 28181 79781 28215 79815
rect 28215 79781 28224 79815
rect 28632 79840 28684 79892
rect 29184 79840 29236 79892
rect 28172 79772 28224 79781
rect 29000 79772 29052 79824
rect 26056 79636 26108 79688
rect 37740 79840 37792 79892
rect 25504 79568 25556 79620
rect 30104 79704 30156 79756
rect 36820 79704 36872 79756
rect 37188 79747 37240 79756
rect 37188 79713 37197 79747
rect 37197 79713 37231 79747
rect 37231 79713 37240 79747
rect 37188 79704 37240 79713
rect 29000 79636 29052 79688
rect 33048 79636 33100 79688
rect 1584 79543 1636 79552
rect 1584 79509 1593 79543
rect 1593 79509 1627 79543
rect 1627 79509 1636 79543
rect 1584 79500 1636 79509
rect 26056 79500 26108 79552
rect 28632 79568 28684 79620
rect 31392 79568 31444 79620
rect 28172 79500 28224 79552
rect 30380 79500 30432 79552
rect 4246 79398 4298 79450
rect 4310 79398 4362 79450
rect 4374 79398 4426 79450
rect 4438 79398 4490 79450
rect 34966 79398 35018 79450
rect 35030 79398 35082 79450
rect 35094 79398 35146 79450
rect 35158 79398 35210 79450
rect 21732 79228 21784 79280
rect 25504 79296 25556 79348
rect 28632 79296 28684 79348
rect 2688 79160 2740 79212
rect 1860 79067 1912 79076
rect 1860 79033 1869 79067
rect 1869 79033 1903 79067
rect 1903 79033 1912 79067
rect 1860 79024 1912 79033
rect 2044 79067 2096 79076
rect 2044 79033 2053 79067
rect 2053 79033 2087 79067
rect 2087 79033 2096 79067
rect 2044 79024 2096 79033
rect 22100 79160 22152 79212
rect 25044 79092 25096 79144
rect 27436 79135 27488 79144
rect 27436 79101 27445 79135
rect 27445 79101 27479 79135
rect 27479 79101 27488 79135
rect 27436 79092 27488 79101
rect 28724 79228 28776 79280
rect 30288 79228 30340 79280
rect 25872 79024 25924 79076
rect 36360 79160 36412 79212
rect 28356 79092 28408 79144
rect 37464 79092 37516 79144
rect 37924 79135 37976 79144
rect 37924 79101 37933 79135
rect 37933 79101 37967 79135
rect 37967 79101 37976 79135
rect 37924 79092 37976 79101
rect 28172 78956 28224 79008
rect 28356 78956 28408 79008
rect 29276 79024 29328 79076
rect 28724 78956 28776 79008
rect 19606 78854 19658 78906
rect 19670 78854 19722 78906
rect 19734 78854 19786 78906
rect 19798 78854 19850 78906
rect 1584 78480 1636 78532
rect 26424 78684 26476 78736
rect 28172 78752 28224 78804
rect 38108 78752 38160 78804
rect 25596 78412 25648 78464
rect 27436 78412 27488 78464
rect 28172 78659 28224 78668
rect 28172 78625 28181 78659
rect 28181 78625 28215 78659
rect 28215 78625 28224 78659
rect 28172 78616 28224 78625
rect 28448 78616 28500 78668
rect 28724 78548 28776 78600
rect 30104 78684 30156 78736
rect 37188 78727 37240 78736
rect 37188 78693 37197 78727
rect 37197 78693 37231 78727
rect 37231 78693 37240 78727
rect 37188 78684 37240 78693
rect 30012 78616 30064 78668
rect 29276 78548 29328 78600
rect 28724 78412 28776 78464
rect 29184 78412 29236 78464
rect 32588 78412 32640 78464
rect 35900 78412 35952 78464
rect 4246 78310 4298 78362
rect 4310 78310 4362 78362
rect 4374 78310 4426 78362
rect 4438 78310 4490 78362
rect 34966 78310 35018 78362
rect 35030 78310 35082 78362
rect 35094 78310 35146 78362
rect 35158 78310 35210 78362
rect 28448 78208 28500 78260
rect 24216 78140 24268 78192
rect 31392 78140 31444 78192
rect 1860 78047 1912 78056
rect 1860 78013 1869 78047
rect 1869 78013 1903 78047
rect 1903 78013 1912 78047
rect 1860 78004 1912 78013
rect 29000 78004 29052 78056
rect 37188 78047 37240 78056
rect 37188 78013 37197 78047
rect 37197 78013 37231 78047
rect 37231 78013 37240 78047
rect 37188 78004 37240 78013
rect 29276 77979 29328 77988
rect 29276 77945 29285 77979
rect 29285 77945 29319 77979
rect 29319 77945 29328 77979
rect 29276 77936 29328 77945
rect 35992 77936 36044 77988
rect 37924 77979 37976 77988
rect 1952 77911 2004 77920
rect 1952 77877 1961 77911
rect 1961 77877 1995 77911
rect 1995 77877 2004 77911
rect 1952 77868 2004 77877
rect 25504 77868 25556 77920
rect 29092 77868 29144 77920
rect 37280 77911 37332 77920
rect 37280 77877 37289 77911
rect 37289 77877 37323 77911
rect 37323 77877 37332 77911
rect 37280 77868 37332 77877
rect 37924 77945 37933 77979
rect 37933 77945 37967 77979
rect 37967 77945 37976 77979
rect 37924 77936 37976 77945
rect 19606 77766 19658 77818
rect 19670 77766 19722 77818
rect 19734 77766 19786 77818
rect 19798 77766 19850 77818
rect 20168 77664 20220 77716
rect 37280 77664 37332 77716
rect 1400 77571 1452 77580
rect 1400 77537 1409 77571
rect 1409 77537 1443 77571
rect 1443 77537 1452 77571
rect 1400 77528 1452 77537
rect 37188 77571 37240 77580
rect 37188 77537 37197 77571
rect 37197 77537 37231 77571
rect 37231 77537 37240 77571
rect 37188 77528 37240 77537
rect 23756 77460 23808 77512
rect 30380 77460 30432 77512
rect 22928 77392 22980 77444
rect 30288 77392 30340 77444
rect 12256 77324 12308 77376
rect 30012 77324 30064 77376
rect 31208 77324 31260 77376
rect 36820 77324 36872 77376
rect 4246 77222 4298 77274
rect 4310 77222 4362 77274
rect 4374 77222 4426 77274
rect 4438 77222 4490 77274
rect 34966 77222 35018 77274
rect 35030 77222 35082 77274
rect 35094 77222 35146 77274
rect 35158 77222 35210 77274
rect 29000 77052 29052 77104
rect 29460 77052 29512 77104
rect 24860 76848 24912 76900
rect 29276 76848 29328 76900
rect 37924 76891 37976 76900
rect 37924 76857 37933 76891
rect 37933 76857 37967 76891
rect 37967 76857 37976 76891
rect 37924 76848 37976 76857
rect 38016 76823 38068 76832
rect 38016 76789 38025 76823
rect 38025 76789 38059 76823
rect 38059 76789 38068 76823
rect 38016 76780 38068 76789
rect 19606 76678 19658 76730
rect 19670 76678 19722 76730
rect 19734 76678 19786 76730
rect 19798 76678 19850 76730
rect 23020 76576 23072 76628
rect 38016 76576 38068 76628
rect 1400 76483 1452 76492
rect 1400 76449 1409 76483
rect 1409 76449 1443 76483
rect 1443 76449 1452 76483
rect 1400 76440 1452 76449
rect 24860 76440 24912 76492
rect 37188 76483 37240 76492
rect 37188 76449 37197 76483
rect 37197 76449 37231 76483
rect 37231 76449 37240 76483
rect 37188 76440 37240 76449
rect 8300 76236 8352 76288
rect 19248 76236 19300 76288
rect 31576 76236 31628 76288
rect 4246 76134 4298 76186
rect 4310 76134 4362 76186
rect 4374 76134 4426 76186
rect 4438 76134 4490 76186
rect 34966 76134 35018 76186
rect 35030 76134 35082 76186
rect 35094 76134 35146 76186
rect 35158 76134 35210 76186
rect 32588 75896 32640 75948
rect 38292 75896 38344 75948
rect 22744 75828 22796 75880
rect 24860 75828 24912 75880
rect 37188 75871 37240 75880
rect 37188 75837 37197 75871
rect 37197 75837 37231 75871
rect 37231 75837 37240 75871
rect 37188 75828 37240 75837
rect 1860 75803 1912 75812
rect 1860 75769 1869 75803
rect 1869 75769 1903 75803
rect 1903 75769 1912 75803
rect 1860 75760 1912 75769
rect 36084 75760 36136 75812
rect 37924 75803 37976 75812
rect 9680 75692 9732 75744
rect 26424 75692 26476 75744
rect 33968 75692 34020 75744
rect 36176 75692 36228 75744
rect 37280 75735 37332 75744
rect 37280 75701 37289 75735
rect 37289 75701 37323 75735
rect 37323 75701 37332 75735
rect 37280 75692 37332 75701
rect 37924 75769 37933 75803
rect 37933 75769 37967 75803
rect 37967 75769 37976 75803
rect 37924 75760 37976 75769
rect 19606 75590 19658 75642
rect 19670 75590 19722 75642
rect 19734 75590 19786 75642
rect 19798 75590 19850 75642
rect 19156 75488 19208 75540
rect 37280 75488 37332 75540
rect 26424 75352 26476 75404
rect 26884 75352 26936 75404
rect 29552 75352 29604 75404
rect 30288 75352 30340 75404
rect 37188 75395 37240 75404
rect 37188 75361 37197 75395
rect 37197 75361 37231 75395
rect 37231 75361 37240 75395
rect 37188 75352 37240 75361
rect 29184 75216 29236 75268
rect 29552 75216 29604 75268
rect 26516 75148 26568 75200
rect 26976 75148 27028 75200
rect 36360 75148 36412 75200
rect 4246 75046 4298 75098
rect 4310 75046 4362 75098
rect 4374 75046 4426 75098
rect 4438 75046 4490 75098
rect 34966 75046 35018 75098
rect 35030 75046 35082 75098
rect 35094 75046 35146 75098
rect 35158 75046 35210 75098
rect 1860 74783 1912 74792
rect 1860 74749 1869 74783
rect 1869 74749 1903 74783
rect 1903 74749 1912 74783
rect 1860 74740 1912 74749
rect 9220 74672 9272 74724
rect 37924 74715 37976 74724
rect 37924 74681 37933 74715
rect 37933 74681 37967 74715
rect 37967 74681 37976 74715
rect 37924 74672 37976 74681
rect 20260 74604 20312 74656
rect 19606 74502 19658 74554
rect 19670 74502 19722 74554
rect 19734 74502 19786 74554
rect 19798 74502 19850 74554
rect 1860 74307 1912 74316
rect 1860 74273 1869 74307
rect 1869 74273 1903 74307
rect 1903 74273 1912 74307
rect 1860 74264 1912 74273
rect 37188 74307 37240 74316
rect 37188 74273 37197 74307
rect 37197 74273 37231 74307
rect 37231 74273 37240 74307
rect 37188 74264 37240 74273
rect 27436 74196 27488 74248
rect 28172 74196 28224 74248
rect 8944 74128 8996 74180
rect 22192 74060 22244 74112
rect 4246 73958 4298 74010
rect 4310 73958 4362 74010
rect 4374 73958 4426 74010
rect 4438 73958 4490 74010
rect 34966 73958 35018 74010
rect 35030 73958 35082 74010
rect 35094 73958 35146 74010
rect 35158 73958 35210 74010
rect 28632 73856 28684 73908
rect 29276 73652 29328 73704
rect 37188 73695 37240 73704
rect 37188 73661 37197 73695
rect 37197 73661 37231 73695
rect 37231 73661 37240 73695
rect 37188 73652 37240 73661
rect 37924 73627 37976 73636
rect 37924 73593 37933 73627
rect 37933 73593 37967 73627
rect 37967 73593 37976 73627
rect 37924 73584 37976 73593
rect 37280 73559 37332 73568
rect 37280 73525 37289 73559
rect 37289 73525 37323 73559
rect 37323 73525 37332 73559
rect 37280 73516 37332 73525
rect 38016 73559 38068 73568
rect 38016 73525 38025 73559
rect 38025 73525 38059 73559
rect 38059 73525 38068 73559
rect 38016 73516 38068 73525
rect 19606 73414 19658 73466
rect 19670 73414 19722 73466
rect 19734 73414 19786 73466
rect 19798 73414 19850 73466
rect 20352 73312 20404 73364
rect 37280 73312 37332 73364
rect 17868 73244 17920 73296
rect 38016 73244 38068 73296
rect 1860 73219 1912 73228
rect 1860 73185 1869 73219
rect 1869 73185 1903 73219
rect 1903 73185 1912 73219
rect 1860 73176 1912 73185
rect 6276 73176 6328 73228
rect 8300 73176 8352 73228
rect 12164 73176 12216 73228
rect 37188 73219 37240 73228
rect 37188 73185 37197 73219
rect 37197 73185 37231 73219
rect 37231 73185 37240 73219
rect 37188 73176 37240 73185
rect 37096 72972 37148 73024
rect 4246 72870 4298 72922
rect 4310 72870 4362 72922
rect 4374 72870 4426 72922
rect 4438 72870 4490 72922
rect 34966 72870 35018 72922
rect 35030 72870 35082 72922
rect 35094 72870 35146 72922
rect 35158 72870 35210 72922
rect 37924 72607 37976 72616
rect 37924 72573 37933 72607
rect 37933 72573 37967 72607
rect 37967 72573 37976 72607
rect 37924 72564 37976 72573
rect 1860 72539 1912 72548
rect 1860 72505 1869 72539
rect 1869 72505 1903 72539
rect 1903 72505 1912 72539
rect 1860 72496 1912 72505
rect 4804 72496 4856 72548
rect 37648 72428 37700 72480
rect 19606 72326 19658 72378
rect 19670 72326 19722 72378
rect 19734 72326 19786 72378
rect 19798 72326 19850 72378
rect 37188 72131 37240 72140
rect 37188 72097 37197 72131
rect 37197 72097 37231 72131
rect 37231 72097 37240 72131
rect 37188 72088 37240 72097
rect 38384 71952 38436 72004
rect 4246 71782 4298 71834
rect 4310 71782 4362 71834
rect 4374 71782 4426 71834
rect 4438 71782 4490 71834
rect 34966 71782 35018 71834
rect 35030 71782 35082 71834
rect 35094 71782 35146 71834
rect 35158 71782 35210 71834
rect 33968 71723 34020 71732
rect 33968 71689 33977 71723
rect 33977 71689 34011 71723
rect 34011 71689 34020 71723
rect 33968 71680 34020 71689
rect 1860 71519 1912 71528
rect 1860 71485 1869 71519
rect 1869 71485 1903 71519
rect 1903 71485 1912 71519
rect 1860 71476 1912 71485
rect 33692 71476 33744 71528
rect 37188 71519 37240 71528
rect 37188 71485 37197 71519
rect 37197 71485 37231 71519
rect 37231 71485 37240 71519
rect 37188 71476 37240 71485
rect 39120 71476 39172 71528
rect 3516 71408 3568 71460
rect 37924 71451 37976 71460
rect 37924 71417 37933 71451
rect 37933 71417 37967 71451
rect 37967 71417 37976 71451
rect 37924 71408 37976 71417
rect 39488 71408 39540 71460
rect 19606 71238 19658 71290
rect 19670 71238 19722 71290
rect 19734 71238 19786 71290
rect 19798 71238 19850 71290
rect 1860 71043 1912 71052
rect 1860 71009 1869 71043
rect 1869 71009 1903 71043
rect 1903 71009 1912 71043
rect 1860 71000 1912 71009
rect 3700 71000 3752 71052
rect 15292 71000 15344 71052
rect 37188 71043 37240 71052
rect 37188 71009 37197 71043
rect 37197 71009 37231 71043
rect 37231 71009 37240 71043
rect 37188 71000 37240 71009
rect 6368 70864 6420 70916
rect 38292 70864 38344 70916
rect 4246 70694 4298 70746
rect 4310 70694 4362 70746
rect 4374 70694 4426 70746
rect 4438 70694 4490 70746
rect 34966 70694 35018 70746
rect 35030 70694 35082 70746
rect 35094 70694 35146 70746
rect 35158 70694 35210 70746
rect 21640 70388 21692 70440
rect 37924 70431 37976 70440
rect 37924 70397 37933 70431
rect 37933 70397 37967 70431
rect 37967 70397 37976 70431
rect 37924 70388 37976 70397
rect 19606 70150 19658 70202
rect 19670 70150 19722 70202
rect 19734 70150 19786 70202
rect 19798 70150 19850 70202
rect 1860 69955 1912 69964
rect 1860 69921 1869 69955
rect 1869 69921 1903 69955
rect 1903 69921 1912 69955
rect 1860 69912 1912 69921
rect 37188 69955 37240 69964
rect 37188 69921 37197 69955
rect 37197 69921 37231 69955
rect 37231 69921 37240 69955
rect 37188 69912 37240 69921
rect 3424 69776 3476 69828
rect 23204 69708 23256 69760
rect 4246 69606 4298 69658
rect 4310 69606 4362 69658
rect 4374 69606 4426 69658
rect 4438 69606 4490 69658
rect 34966 69606 35018 69658
rect 35030 69606 35082 69658
rect 35094 69606 35146 69658
rect 35158 69606 35210 69658
rect 18972 69300 19024 69352
rect 17776 69164 17828 69216
rect 37188 69275 37240 69284
rect 37188 69241 37197 69275
rect 37197 69241 37231 69275
rect 37231 69241 37240 69275
rect 37188 69232 37240 69241
rect 37924 69275 37976 69284
rect 37924 69241 37933 69275
rect 37933 69241 37967 69275
rect 37967 69241 37976 69275
rect 37924 69232 37976 69241
rect 19606 69062 19658 69114
rect 19670 69062 19722 69114
rect 19734 69062 19786 69114
rect 19798 69062 19850 69114
rect 1860 68935 1912 68944
rect 1860 68901 1869 68935
rect 1869 68901 1903 68935
rect 1903 68901 1912 68935
rect 1860 68892 1912 68901
rect 29184 68892 29236 68944
rect 34060 68892 34112 68944
rect 37188 68867 37240 68876
rect 37188 68833 37197 68867
rect 37197 68833 37231 68867
rect 37231 68833 37240 68867
rect 37188 68824 37240 68833
rect 2136 68688 2188 68740
rect 38844 68620 38896 68672
rect 4246 68518 4298 68570
rect 4310 68518 4362 68570
rect 4374 68518 4426 68570
rect 4438 68518 4490 68570
rect 34966 68518 35018 68570
rect 35030 68518 35082 68570
rect 35094 68518 35146 68570
rect 35158 68518 35210 68570
rect 3148 68280 3200 68332
rect 22008 68280 22060 68332
rect 1860 68255 1912 68264
rect 1860 68221 1869 68255
rect 1869 68221 1903 68255
rect 1903 68221 1912 68255
rect 1860 68212 1912 68221
rect 37280 68255 37332 68264
rect 37280 68221 37289 68255
rect 37289 68221 37323 68255
rect 37323 68221 37332 68255
rect 37280 68212 37332 68221
rect 9036 68144 9088 68196
rect 37832 68076 37884 68128
rect 38200 68076 38252 68128
rect 19606 67974 19658 68026
rect 19670 67974 19722 68026
rect 19734 67974 19786 68026
rect 19798 67974 19850 68026
rect 37188 67779 37240 67788
rect 37188 67745 37197 67779
rect 37197 67745 37231 67779
rect 37231 67745 37240 67779
rect 37188 67736 37240 67745
rect 33508 67600 33560 67652
rect 34704 67600 34756 67652
rect 37372 67643 37424 67652
rect 37372 67609 37381 67643
rect 37381 67609 37415 67643
rect 37415 67609 37424 67643
rect 37372 67600 37424 67609
rect 38936 67643 38988 67652
rect 38936 67609 38945 67643
rect 38945 67609 38979 67643
rect 38979 67609 38988 67643
rect 38936 67600 38988 67609
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 34966 67430 35018 67482
rect 35030 67430 35082 67482
rect 35094 67430 35146 67482
rect 35158 67430 35210 67482
rect 38752 67260 38804 67312
rect 1400 67167 1452 67176
rect 1400 67133 1409 67167
rect 1409 67133 1443 67167
rect 1443 67133 1452 67167
rect 1400 67124 1452 67133
rect 37280 67167 37332 67176
rect 37280 67133 37289 67167
rect 37289 67133 37323 67167
rect 37323 67133 37332 67167
rect 37280 67124 37332 67133
rect 37924 67167 37976 67176
rect 37924 67133 37933 67167
rect 37933 67133 37967 67167
rect 37967 67133 37976 67167
rect 37924 67124 37976 67133
rect 7748 66988 7800 67040
rect 38660 66988 38712 67040
rect 19606 66886 19658 66938
rect 19670 66886 19722 66938
rect 19734 66886 19786 66938
rect 19798 66886 19850 66938
rect 1400 66691 1452 66700
rect 1400 66657 1409 66691
rect 1409 66657 1443 66691
rect 1443 66657 1452 66691
rect 1400 66648 1452 66657
rect 2228 66444 2280 66496
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 34966 66342 35018 66394
rect 35030 66342 35082 66394
rect 35094 66342 35146 66394
rect 35158 66342 35210 66394
rect 38568 66172 38620 66224
rect 37280 66079 37332 66088
rect 37280 66045 37289 66079
rect 37289 66045 37323 66079
rect 37323 66045 37332 66079
rect 37280 66036 37332 66045
rect 37924 66079 37976 66088
rect 37924 66045 37933 66079
rect 37933 66045 37967 66079
rect 37967 66045 37976 66079
rect 37924 66036 37976 66045
rect 38844 65900 38896 65952
rect 19606 65798 19658 65850
rect 19670 65798 19722 65850
rect 19734 65798 19786 65850
rect 19798 65798 19850 65850
rect 1400 65603 1452 65612
rect 1400 65569 1409 65603
rect 1409 65569 1443 65603
rect 1443 65569 1452 65603
rect 1400 65560 1452 65569
rect 34704 65560 34756 65612
rect 35532 65560 35584 65612
rect 37188 65603 37240 65612
rect 37188 65569 37197 65603
rect 37197 65569 37231 65603
rect 37231 65569 37240 65603
rect 37188 65560 37240 65569
rect 1952 65492 2004 65544
rect 12992 65492 13044 65544
rect 33324 65492 33376 65544
rect 34060 65492 34112 65544
rect 32864 65424 32916 65476
rect 34796 65424 34848 65476
rect 1676 65356 1728 65408
rect 39580 65356 39632 65408
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 34966 65254 35018 65306
rect 35030 65254 35082 65306
rect 35094 65254 35146 65306
rect 35158 65254 35210 65306
rect 9128 65084 9180 65136
rect 33876 65084 33928 65136
rect 1400 64991 1452 65000
rect 1400 64957 1409 64991
rect 1409 64957 1443 64991
rect 1443 64957 1452 64991
rect 1400 64948 1452 64957
rect 34152 64948 34204 65000
rect 35256 64948 35308 65000
rect 37188 64948 37240 65000
rect 37924 64991 37976 65000
rect 37924 64957 37933 64991
rect 37933 64957 37967 64991
rect 37967 64957 37976 64991
rect 37924 64948 37976 64957
rect 19984 64880 20036 64932
rect 19606 64710 19658 64762
rect 19670 64710 19722 64762
rect 19734 64710 19786 64762
rect 19798 64710 19850 64762
rect 34612 64651 34664 64660
rect 34612 64617 34621 64651
rect 34621 64617 34655 64651
rect 34655 64617 34664 64651
rect 34612 64608 34664 64617
rect 34244 64472 34296 64524
rect 33968 64404 34020 64456
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 34966 64166 35018 64218
rect 35030 64166 35082 64218
rect 35094 64166 35146 64218
rect 35158 64166 35210 64218
rect 15292 64107 15344 64116
rect 15292 64073 15301 64107
rect 15301 64073 15335 64107
rect 15335 64073 15344 64107
rect 15292 64064 15344 64073
rect 34152 64064 34204 64116
rect 33968 63928 34020 63980
rect 1400 63903 1452 63912
rect 1400 63869 1409 63903
rect 1409 63869 1443 63903
rect 1443 63869 1452 63903
rect 1400 63860 1452 63869
rect 34152 63903 34204 63912
rect 34152 63869 34161 63903
rect 34161 63869 34195 63903
rect 34195 63869 34204 63903
rect 34152 63860 34204 63869
rect 37280 63903 37332 63912
rect 37280 63869 37289 63903
rect 37289 63869 37323 63903
rect 37323 63869 37332 63903
rect 37280 63860 37332 63869
rect 37924 63903 37976 63912
rect 37924 63869 37933 63903
rect 37933 63869 37967 63903
rect 37967 63869 37976 63903
rect 37924 63860 37976 63869
rect 15200 63835 15252 63844
rect 15200 63801 15209 63835
rect 15209 63801 15243 63835
rect 15243 63801 15252 63835
rect 15200 63792 15252 63801
rect 33324 63792 33376 63844
rect 34888 63792 34940 63844
rect 7564 63724 7616 63776
rect 34612 63724 34664 63776
rect 19606 63622 19658 63674
rect 19670 63622 19722 63674
rect 19734 63622 19786 63674
rect 19798 63622 19850 63674
rect 22008 63520 22060 63572
rect 34888 63520 34940 63572
rect 35440 63563 35492 63572
rect 35440 63529 35449 63563
rect 35449 63529 35483 63563
rect 35483 63529 35492 63563
rect 35440 63520 35492 63529
rect 36452 63563 36504 63572
rect 36452 63529 36461 63563
rect 36461 63529 36495 63563
rect 36495 63529 36504 63563
rect 36452 63520 36504 63529
rect 32956 63452 33008 63504
rect 1400 63427 1452 63436
rect 1400 63393 1409 63427
rect 1409 63393 1443 63427
rect 1443 63393 1452 63427
rect 1400 63384 1452 63393
rect 33140 63427 33192 63436
rect 33140 63393 33149 63427
rect 33149 63393 33183 63427
rect 33183 63393 33192 63427
rect 33140 63384 33192 63393
rect 33508 63384 33560 63436
rect 33876 63384 33928 63436
rect 34520 63452 34572 63504
rect 20904 63316 20956 63368
rect 20536 63248 20588 63300
rect 35256 63384 35308 63436
rect 37188 63427 37240 63436
rect 37188 63393 37197 63427
rect 37197 63393 37231 63427
rect 37231 63393 37240 63427
rect 37188 63384 37240 63393
rect 9496 63180 9548 63232
rect 32404 63180 32456 63232
rect 34704 63180 34756 63232
rect 38476 63180 38528 63232
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 34966 63078 35018 63130
rect 35030 63078 35082 63130
rect 35094 63078 35146 63130
rect 35158 63078 35210 63130
rect 29092 62976 29144 63028
rect 32404 62976 32456 63028
rect 33048 63019 33100 63028
rect 33048 62985 33057 63019
rect 33057 62985 33091 63019
rect 33091 62985 33100 63019
rect 33048 62976 33100 62985
rect 31760 62908 31812 62960
rect 8944 62840 8996 62892
rect 10048 62840 10100 62892
rect 33048 62840 33100 62892
rect 34152 62840 34204 62892
rect 34980 62840 35032 62892
rect 35256 62840 35308 62892
rect 8024 62772 8076 62824
rect 21456 62772 21508 62824
rect 24584 62772 24636 62824
rect 24768 62772 24820 62824
rect 32956 62815 33008 62824
rect 32956 62781 32965 62815
rect 32965 62781 32999 62815
rect 32999 62781 33008 62815
rect 32956 62772 33008 62781
rect 37280 62815 37332 62824
rect 37280 62781 37289 62815
rect 37289 62781 37323 62815
rect 37323 62781 37332 62815
rect 37280 62772 37332 62781
rect 37924 62815 37976 62824
rect 37924 62781 37933 62815
rect 37933 62781 37967 62815
rect 37967 62781 37976 62815
rect 37924 62772 37976 62781
rect 32128 62704 32180 62756
rect 32404 62636 32456 62688
rect 33968 62636 34020 62688
rect 34152 62636 34204 62688
rect 37464 62679 37516 62688
rect 37464 62645 37473 62679
rect 37473 62645 37507 62679
rect 37507 62645 37516 62679
rect 37464 62636 37516 62645
rect 38108 62679 38160 62688
rect 38108 62645 38117 62679
rect 38117 62645 38151 62679
rect 38151 62645 38160 62679
rect 38108 62636 38160 62645
rect 19606 62534 19658 62586
rect 19670 62534 19722 62586
rect 19734 62534 19786 62586
rect 19798 62534 19850 62586
rect 32956 62432 33008 62484
rect 22836 62364 22888 62416
rect 31760 62364 31812 62416
rect 1400 62339 1452 62348
rect 1400 62305 1409 62339
rect 1409 62305 1443 62339
rect 1443 62305 1452 62339
rect 1400 62296 1452 62305
rect 24308 62296 24360 62348
rect 29920 62339 29972 62348
rect 29920 62305 29929 62339
rect 29929 62305 29963 62339
rect 29963 62305 29972 62339
rect 29920 62296 29972 62305
rect 33048 62296 33100 62348
rect 33784 62364 33836 62416
rect 34980 62339 35032 62348
rect 21180 62228 21232 62280
rect 34980 62305 34989 62339
rect 34989 62305 35023 62339
rect 35023 62305 35032 62339
rect 34980 62296 35032 62305
rect 35348 62339 35400 62348
rect 35348 62305 35357 62339
rect 35357 62305 35391 62339
rect 35391 62305 35400 62339
rect 35348 62296 35400 62305
rect 23112 62160 23164 62212
rect 38108 62160 38160 62212
rect 7840 62092 7892 62144
rect 33876 62092 33928 62144
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 34966 61990 35018 62042
rect 35030 61990 35082 62042
rect 35094 61990 35146 62042
rect 35158 61990 35210 62042
rect 1400 61727 1452 61736
rect 1400 61693 1409 61727
rect 1409 61693 1443 61727
rect 1443 61693 1452 61727
rect 1400 61684 1452 61693
rect 37280 61727 37332 61736
rect 37280 61693 37289 61727
rect 37289 61693 37323 61727
rect 37323 61693 37332 61727
rect 37280 61684 37332 61693
rect 37924 61727 37976 61736
rect 37924 61693 37933 61727
rect 37933 61693 37967 61727
rect 37967 61693 37976 61727
rect 37924 61684 37976 61693
rect 8484 61548 8536 61600
rect 35348 61548 35400 61600
rect 38108 61591 38160 61600
rect 38108 61557 38117 61591
rect 38117 61557 38151 61591
rect 38151 61557 38160 61591
rect 38108 61548 38160 61557
rect 19606 61446 19658 61498
rect 19670 61446 19722 61498
rect 19734 61446 19786 61498
rect 19798 61446 19850 61498
rect 23388 61276 23440 61328
rect 38108 61276 38160 61328
rect 37188 61251 37240 61260
rect 37188 61217 37197 61251
rect 37197 61217 37231 61251
rect 37231 61217 37240 61251
rect 37188 61208 37240 61217
rect 34796 61004 34848 61056
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 34966 60902 35018 60954
rect 35030 60902 35082 60954
rect 35094 60902 35146 60954
rect 35158 60902 35210 60954
rect 1400 60639 1452 60648
rect 1400 60605 1409 60639
rect 1409 60605 1443 60639
rect 1443 60605 1452 60639
rect 1400 60596 1452 60605
rect 28632 60800 28684 60852
rect 35716 60800 35768 60852
rect 26516 60639 26568 60648
rect 24400 60528 24452 60580
rect 6552 60460 6604 60512
rect 25872 60460 25924 60512
rect 26516 60605 26525 60639
rect 26525 60605 26559 60639
rect 26559 60605 26568 60639
rect 26516 60596 26568 60605
rect 30104 60596 30156 60648
rect 37280 60639 37332 60648
rect 37280 60605 37289 60639
rect 37289 60605 37323 60639
rect 37323 60605 37332 60639
rect 37280 60596 37332 60605
rect 37924 60639 37976 60648
rect 37924 60605 37933 60639
rect 37933 60605 37967 60639
rect 37967 60605 37976 60639
rect 37924 60596 37976 60605
rect 29552 60528 29604 60580
rect 37464 60503 37516 60512
rect 37464 60469 37473 60503
rect 37473 60469 37507 60503
rect 37507 60469 37516 60503
rect 37464 60460 37516 60469
rect 38108 60503 38160 60512
rect 38108 60469 38117 60503
rect 38117 60469 38151 60503
rect 38151 60469 38160 60503
rect 38108 60460 38160 60469
rect 19606 60358 19658 60410
rect 19670 60358 19722 60410
rect 19734 60358 19786 60410
rect 19798 60358 19850 60410
rect 18328 60256 18380 60308
rect 38108 60256 38160 60308
rect 18512 60188 18564 60240
rect 37464 60188 37516 60240
rect 1400 60163 1452 60172
rect 1400 60129 1409 60163
rect 1409 60129 1443 60163
rect 1443 60129 1452 60163
rect 1400 60120 1452 60129
rect 37188 60163 37240 60172
rect 37188 60129 37197 60163
rect 37197 60129 37231 60163
rect 37231 60129 37240 60163
rect 37188 60120 37240 60129
rect 26332 59984 26384 60036
rect 27436 59984 27488 60036
rect 37280 59984 37332 60036
rect 39212 59984 39264 60036
rect 8944 59916 8996 59968
rect 19984 59916 20036 59968
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 34966 59814 35018 59866
rect 35030 59814 35082 59866
rect 35094 59814 35146 59866
rect 35158 59814 35210 59866
rect 18788 59576 18840 59628
rect 23296 59576 23348 59628
rect 26240 59551 26292 59560
rect 26240 59517 26249 59551
rect 26249 59517 26283 59551
rect 26283 59517 26292 59551
rect 26240 59508 26292 59517
rect 36728 59712 36780 59764
rect 36544 59576 36596 59628
rect 36820 59576 36872 59628
rect 36912 59551 36964 59560
rect 24492 59372 24544 59424
rect 36912 59517 36921 59551
rect 36921 59517 36955 59551
rect 36955 59517 36964 59551
rect 36912 59508 36964 59517
rect 37280 59508 37332 59560
rect 37740 59551 37792 59560
rect 37740 59517 37749 59551
rect 37749 59517 37783 59551
rect 37783 59517 37792 59551
rect 37740 59508 37792 59517
rect 38016 59508 38068 59560
rect 36728 59440 36780 59492
rect 36268 59372 36320 59424
rect 36820 59372 36872 59424
rect 19606 59270 19658 59322
rect 19670 59270 19722 59322
rect 19734 59270 19786 59322
rect 19798 59270 19850 59322
rect 7288 59100 7340 59152
rect 7656 59100 7708 59152
rect 1400 59075 1452 59084
rect 1400 59041 1409 59075
rect 1409 59041 1443 59075
rect 1443 59041 1452 59075
rect 1400 59032 1452 59041
rect 12256 59075 12308 59084
rect 12256 59041 12265 59075
rect 12265 59041 12299 59075
rect 12299 59041 12308 59075
rect 12256 59032 12308 59041
rect 36452 59075 36504 59084
rect 36452 59041 36461 59075
rect 36461 59041 36495 59075
rect 36495 59041 36504 59075
rect 36452 59032 36504 59041
rect 37188 59075 37240 59084
rect 37188 59041 37197 59075
rect 37197 59041 37231 59075
rect 37231 59041 37240 59075
rect 37188 59032 37240 59041
rect 11980 58964 12032 59016
rect 36360 58964 36412 59016
rect 37004 58964 37056 59016
rect 33968 58896 34020 58948
rect 34336 58896 34388 58948
rect 35256 58896 35308 58948
rect 1584 58871 1636 58880
rect 1584 58837 1593 58871
rect 1593 58837 1627 58871
rect 1627 58837 1636 58871
rect 1584 58828 1636 58837
rect 17316 58828 17368 58880
rect 20812 58828 20864 58880
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 34966 58726 35018 58778
rect 35030 58726 35082 58778
rect 35094 58726 35146 58778
rect 35158 58726 35210 58778
rect 27160 58667 27212 58676
rect 2044 58488 2096 58540
rect 1400 58463 1452 58472
rect 1400 58429 1409 58463
rect 1409 58429 1443 58463
rect 1443 58429 1452 58463
rect 1400 58420 1452 58429
rect 11980 58352 12032 58404
rect 26240 58488 26292 58540
rect 12992 58463 13044 58472
rect 12992 58429 13001 58463
rect 13001 58429 13035 58463
rect 13035 58429 13044 58463
rect 12992 58420 13044 58429
rect 27160 58633 27169 58667
rect 27169 58633 27203 58667
rect 27203 58633 27212 58667
rect 27160 58624 27212 58633
rect 35900 58624 35952 58676
rect 38016 58624 38068 58676
rect 34336 58556 34388 58608
rect 37004 58556 37056 58608
rect 26516 58488 26568 58540
rect 36728 58488 36780 58540
rect 26240 58352 26292 58404
rect 1768 58284 1820 58336
rect 12348 58327 12400 58336
rect 12348 58293 12357 58327
rect 12357 58293 12391 58327
rect 12391 58293 12400 58327
rect 12348 58284 12400 58293
rect 17500 58284 17552 58336
rect 18052 58284 18104 58336
rect 35992 58420 36044 58472
rect 36360 58420 36412 58472
rect 36452 58420 36504 58472
rect 36912 58463 36964 58472
rect 36912 58429 36921 58463
rect 36921 58429 36955 58463
rect 36955 58429 36964 58463
rect 37556 58463 37608 58472
rect 36912 58420 36964 58429
rect 37556 58429 37565 58463
rect 37565 58429 37599 58463
rect 37599 58429 37608 58463
rect 37556 58420 37608 58429
rect 37740 58395 37792 58404
rect 37740 58361 37749 58395
rect 37749 58361 37783 58395
rect 37783 58361 37792 58395
rect 37740 58352 37792 58361
rect 35992 58284 36044 58336
rect 38108 58327 38160 58336
rect 38108 58293 38117 58327
rect 38117 58293 38151 58327
rect 38151 58293 38160 58327
rect 38108 58284 38160 58293
rect 19606 58182 19658 58234
rect 19670 58182 19722 58234
rect 19734 58182 19786 58234
rect 19798 58182 19850 58234
rect 26792 58080 26844 58132
rect 27160 58080 27212 58132
rect 11980 57944 12032 57996
rect 12164 57944 12216 57996
rect 12440 57987 12492 57996
rect 12440 57953 12449 57987
rect 12449 57953 12483 57987
rect 12483 57953 12492 57987
rect 36452 57987 36504 57996
rect 12440 57944 12492 57953
rect 36452 57953 36461 57987
rect 36461 57953 36495 57987
rect 36495 57953 36504 57987
rect 36452 57944 36504 57953
rect 36728 57944 36780 57996
rect 37004 57944 37056 57996
rect 37188 57987 37240 57996
rect 37188 57953 37197 57987
rect 37197 57953 37231 57987
rect 37231 57953 37240 57987
rect 37188 57944 37240 57953
rect 9036 57876 9088 57928
rect 10508 57876 10560 57928
rect 20168 57876 20220 57928
rect 20628 57876 20680 57928
rect 22284 57876 22336 57928
rect 28540 57876 28592 57928
rect 25228 57808 25280 57860
rect 27436 57808 27488 57860
rect 18880 57740 18932 57792
rect 36544 57783 36596 57792
rect 36544 57749 36553 57783
rect 36553 57749 36587 57783
rect 36587 57749 36596 57783
rect 36544 57740 36596 57749
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 21824 57536 21876 57588
rect 27436 57536 27488 57588
rect 36544 57536 36596 57588
rect 20536 57468 20588 57520
rect 26516 57400 26568 57452
rect 1400 57375 1452 57384
rect 1400 57341 1409 57375
rect 1409 57341 1443 57375
rect 1443 57341 1452 57375
rect 1400 57332 1452 57341
rect 25596 57332 25648 57384
rect 17224 57264 17276 57316
rect 3608 57196 3660 57248
rect 26240 57264 26292 57316
rect 28632 57400 28684 57452
rect 34704 57400 34756 57452
rect 29368 57264 29420 57316
rect 32588 57332 32640 57384
rect 37004 57332 37056 57384
rect 39396 57400 39448 57452
rect 38016 57332 38068 57384
rect 37280 57264 37332 57316
rect 37740 57307 37792 57316
rect 37740 57273 37749 57307
rect 37749 57273 37783 57307
rect 37783 57273 37792 57307
rect 37740 57264 37792 57273
rect 39212 57264 39264 57316
rect 37556 57196 37608 57248
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 1584 56992 1636 57044
rect 5080 56992 5132 57044
rect 7012 56992 7064 57044
rect 8300 56924 8352 56976
rect 17224 56924 17276 56976
rect 1400 56899 1452 56908
rect 1400 56865 1409 56899
rect 1409 56865 1443 56899
rect 1443 56865 1452 56899
rect 1400 56856 1452 56865
rect 26516 56992 26568 57044
rect 27528 56992 27580 57044
rect 35808 56992 35860 57044
rect 38108 56992 38160 57044
rect 26884 56924 26936 56976
rect 26516 56856 26568 56908
rect 18236 56720 18288 56772
rect 1584 56695 1636 56704
rect 1584 56661 1593 56695
rect 1593 56661 1627 56695
rect 1627 56661 1636 56695
rect 1584 56652 1636 56661
rect 26516 56652 26568 56704
rect 27528 56856 27580 56908
rect 34520 56924 34572 56976
rect 36452 56967 36504 56976
rect 36452 56933 36461 56967
rect 36461 56933 36495 56967
rect 36495 56933 36504 56967
rect 36452 56924 36504 56933
rect 37188 56899 37240 56908
rect 37188 56865 37197 56899
rect 37197 56865 37231 56899
rect 37231 56865 37240 56899
rect 37188 56856 37240 56865
rect 28540 56788 28592 56840
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 9128 56448 9180 56500
rect 9772 56448 9824 56500
rect 26884 56312 26936 56364
rect 27620 56448 27672 56500
rect 32956 56448 33008 56500
rect 37280 56448 37332 56500
rect 27528 56380 27580 56432
rect 28816 56380 28868 56432
rect 29920 56312 29972 56364
rect 26240 56176 26292 56228
rect 26884 56219 26936 56228
rect 26884 56185 26893 56219
rect 26893 56185 26927 56219
rect 26927 56185 26936 56219
rect 26884 56176 26936 56185
rect 8392 56108 8444 56160
rect 28632 56244 28684 56296
rect 27620 56176 27672 56228
rect 34060 56176 34112 56228
rect 36544 56380 36596 56432
rect 37188 56380 37240 56432
rect 35808 56244 35860 56296
rect 35716 56176 35768 56228
rect 36360 56244 36412 56296
rect 37832 56244 37884 56296
rect 36544 56219 36596 56228
rect 36544 56185 36553 56219
rect 36553 56185 36587 56219
rect 36587 56185 36596 56219
rect 36544 56176 36596 56185
rect 39396 56108 39448 56160
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 26884 55904 26936 55956
rect 28632 55904 28684 55956
rect 36268 55904 36320 55956
rect 6736 55836 6788 55888
rect 17132 55836 17184 55888
rect 33324 55836 33376 55888
rect 33508 55836 33560 55888
rect 34060 55836 34112 55888
rect 35256 55836 35308 55888
rect 1400 55811 1452 55820
rect 1400 55777 1409 55811
rect 1409 55777 1443 55811
rect 1443 55777 1452 55811
rect 1400 55768 1452 55777
rect 34888 55768 34940 55820
rect 1584 55700 1636 55752
rect 6460 55700 6512 55752
rect 21916 55700 21968 55752
rect 36268 55811 36320 55820
rect 36268 55777 36278 55811
rect 36278 55777 36312 55811
rect 36312 55777 36320 55811
rect 36544 55811 36596 55820
rect 36268 55768 36320 55777
rect 36544 55777 36553 55811
rect 36553 55777 36587 55811
rect 36587 55777 36596 55811
rect 36544 55768 36596 55777
rect 38936 55904 38988 55956
rect 36820 55768 36872 55820
rect 29000 55632 29052 55684
rect 4896 55564 4948 55616
rect 35256 55564 35308 55616
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 28632 55360 28684 55412
rect 36452 55360 36504 55412
rect 20076 55292 20128 55344
rect 22100 55292 22152 55344
rect 36360 55292 36412 55344
rect 35716 55224 35768 55276
rect 36452 55224 36504 55276
rect 36912 55292 36964 55344
rect 1400 55199 1452 55208
rect 1400 55165 1409 55199
rect 1409 55165 1443 55199
rect 1443 55165 1452 55199
rect 1400 55156 1452 55165
rect 29092 55199 29144 55208
rect 29092 55165 29101 55199
rect 29101 55165 29135 55199
rect 29135 55165 29144 55199
rect 29092 55156 29144 55165
rect 35440 55156 35492 55208
rect 35992 55156 36044 55208
rect 36360 55199 36412 55208
rect 36360 55165 36367 55199
rect 36367 55165 36412 55199
rect 36360 55156 36412 55165
rect 37188 55224 37240 55276
rect 20628 55088 20680 55140
rect 22284 55088 22336 55140
rect 37372 55156 37424 55208
rect 37924 55199 37976 55208
rect 37924 55165 37933 55199
rect 37933 55165 37967 55199
rect 37967 55165 37976 55199
rect 37924 55156 37976 55165
rect 39304 55156 39356 55208
rect 36544 55131 36596 55140
rect 36544 55097 36553 55131
rect 36553 55097 36587 55131
rect 36587 55097 36596 55131
rect 37740 55131 37792 55140
rect 36544 55088 36596 55097
rect 37740 55097 37749 55131
rect 37749 55097 37783 55131
rect 37783 55097 37792 55131
rect 37740 55088 37792 55097
rect 37832 55131 37884 55140
rect 37832 55097 37841 55131
rect 37841 55097 37875 55131
rect 37875 55097 37884 55131
rect 37832 55088 37884 55097
rect 1584 55063 1636 55072
rect 1584 55029 1593 55063
rect 1593 55029 1627 55063
rect 1627 55029 1636 55063
rect 1584 55020 1636 55029
rect 35164 55020 35216 55072
rect 35440 55020 35492 55072
rect 37464 55020 37516 55072
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 19984 54816 20036 54868
rect 20628 54816 20680 54868
rect 34336 54816 34388 54868
rect 35716 54680 35768 54732
rect 35992 54612 36044 54664
rect 37188 54748 37240 54800
rect 36544 54723 36596 54732
rect 36544 54689 36553 54723
rect 36553 54689 36587 54723
rect 36587 54689 36596 54723
rect 36544 54680 36596 54689
rect 38200 54680 38252 54732
rect 37556 54612 37608 54664
rect 2872 54476 2924 54528
rect 21272 54544 21324 54596
rect 35164 54544 35216 54596
rect 38936 54544 38988 54596
rect 24584 54476 24636 54528
rect 32680 54476 32732 54528
rect 33048 54476 33100 54528
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 36268 54315 36320 54324
rect 36268 54281 36277 54315
rect 36277 54281 36311 54315
rect 36311 54281 36320 54315
rect 36268 54272 36320 54281
rect 35900 54204 35952 54256
rect 1400 54111 1452 54120
rect 1400 54077 1409 54111
rect 1409 54077 1443 54111
rect 1443 54077 1452 54111
rect 1400 54068 1452 54077
rect 25596 54068 25648 54120
rect 31392 54068 31444 54120
rect 35808 54068 35860 54120
rect 37096 54111 37148 54120
rect 37096 54077 37105 54111
rect 37105 54077 37139 54111
rect 37139 54077 37148 54111
rect 37096 54068 37148 54077
rect 39028 54136 39080 54188
rect 38200 54068 38252 54120
rect 36268 54000 36320 54052
rect 36912 54000 36964 54052
rect 37740 54043 37792 54052
rect 37740 54009 37749 54043
rect 37749 54009 37783 54043
rect 37783 54009 37792 54043
rect 37740 54000 37792 54009
rect 37832 54043 37884 54052
rect 37832 54009 37841 54043
rect 37841 54009 37875 54043
rect 37875 54009 37884 54043
rect 37832 54000 37884 54009
rect 1952 53932 2004 53984
rect 35440 53932 35492 53984
rect 35716 53932 35768 53984
rect 35900 53932 35952 53984
rect 37188 53932 37240 53984
rect 37556 53932 37608 53984
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 31760 53728 31812 53780
rect 33968 53728 34020 53780
rect 36452 53728 36504 53780
rect 36728 53728 36780 53780
rect 1400 53635 1452 53644
rect 1400 53601 1409 53635
rect 1409 53601 1443 53635
rect 1443 53601 1452 53635
rect 1400 53592 1452 53601
rect 36728 53635 36780 53644
rect 36728 53601 36737 53635
rect 36737 53601 36771 53635
rect 36771 53601 36780 53635
rect 36728 53592 36780 53601
rect 37372 53635 37424 53644
rect 37372 53601 37381 53635
rect 37381 53601 37415 53635
rect 37415 53601 37424 53635
rect 37372 53592 37424 53601
rect 7932 53388 7984 53440
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 27160 53184 27212 53236
rect 24216 53116 24268 53168
rect 34704 53116 34756 53168
rect 3424 53048 3476 53100
rect 9956 53048 10008 53100
rect 35440 53048 35492 53100
rect 8024 52912 8076 52964
rect 34060 52980 34112 53032
rect 34704 52980 34756 53032
rect 35808 52980 35860 53032
rect 36636 52980 36688 53032
rect 36912 53023 36964 53032
rect 36912 52989 36921 53023
rect 36921 52989 36955 53023
rect 36955 52989 36964 53023
rect 36912 52980 36964 52989
rect 37740 53023 37792 53032
rect 37740 52989 37749 53023
rect 37749 52989 37783 53023
rect 37783 52989 37792 53023
rect 37740 52980 37792 52989
rect 38108 52980 38160 53032
rect 26332 52844 26384 52896
rect 26792 52955 26844 52964
rect 26792 52921 26801 52955
rect 26801 52921 26835 52955
rect 26835 52921 26844 52955
rect 36728 52955 36780 52964
rect 26792 52912 26844 52921
rect 36728 52921 36737 52955
rect 36737 52921 36771 52955
rect 36771 52921 36780 52955
rect 36728 52912 36780 52921
rect 37832 52955 37884 52964
rect 37832 52921 37841 52955
rect 37841 52921 37875 52955
rect 37875 52921 37884 52955
rect 37832 52912 37884 52921
rect 36636 52844 36688 52896
rect 37188 52844 37240 52896
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 36360 52640 36412 52692
rect 36820 52640 36872 52692
rect 1860 52547 1912 52556
rect 1860 52513 1869 52547
rect 1869 52513 1903 52547
rect 1903 52513 1912 52547
rect 1860 52504 1912 52513
rect 7840 52504 7892 52556
rect 8760 52504 8812 52556
rect 20168 52504 20220 52556
rect 28540 52504 28592 52556
rect 36728 52547 36780 52556
rect 36728 52513 36737 52547
rect 36737 52513 36771 52547
rect 36771 52513 36780 52547
rect 36728 52504 36780 52513
rect 37188 52504 37240 52556
rect 18052 52436 18104 52488
rect 34520 52368 34572 52420
rect 36820 52368 36872 52420
rect 21732 52300 21784 52352
rect 27160 52300 27212 52352
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 21732 52096 21784 52148
rect 28816 52096 28868 52148
rect 8300 52028 8352 52080
rect 27528 52028 27580 52080
rect 34336 51960 34388 52012
rect 26792 51935 26844 51944
rect 26792 51901 26801 51935
rect 26801 51901 26835 51935
rect 26835 51901 26844 51935
rect 26792 51892 26844 51901
rect 1860 51867 1912 51876
rect 1860 51833 1869 51867
rect 1869 51833 1903 51867
rect 1903 51833 1912 51867
rect 1860 51824 1912 51833
rect 26332 51824 26384 51876
rect 22192 51756 22244 51808
rect 27160 51892 27212 51944
rect 39028 51892 39080 51944
rect 37740 51867 37792 51876
rect 37740 51833 37749 51867
rect 37749 51833 37783 51867
rect 37783 51833 37792 51867
rect 37740 51824 37792 51833
rect 37832 51867 37884 51876
rect 37832 51833 37841 51867
rect 37841 51833 37875 51867
rect 37875 51833 37884 51867
rect 37832 51824 37884 51833
rect 36452 51756 36504 51808
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 21548 51552 21600 51604
rect 22468 51552 22520 51604
rect 24952 51595 25004 51604
rect 24952 51561 24961 51595
rect 24961 51561 24995 51595
rect 24995 51561 25004 51595
rect 24952 51552 25004 51561
rect 7656 51484 7708 51536
rect 3424 51348 3476 51400
rect 21272 51416 21324 51468
rect 11060 51280 11112 51332
rect 27528 51552 27580 51604
rect 29092 51552 29144 51604
rect 29184 51552 29236 51604
rect 35992 51552 36044 51604
rect 26792 51484 26844 51536
rect 28816 51527 28868 51536
rect 28816 51493 28825 51527
rect 28825 51493 28859 51527
rect 28859 51493 28868 51527
rect 28816 51484 28868 51493
rect 28540 51416 28592 51468
rect 30196 51484 30248 51536
rect 35532 51484 35584 51536
rect 29368 51416 29420 51468
rect 29092 51348 29144 51400
rect 29552 51348 29604 51400
rect 36544 51459 36596 51468
rect 36544 51425 36553 51459
rect 36553 51425 36587 51459
rect 36587 51425 36596 51459
rect 36544 51416 36596 51425
rect 37372 51459 37424 51468
rect 37372 51425 37381 51459
rect 37381 51425 37415 51459
rect 37415 51425 37424 51459
rect 37372 51416 37424 51425
rect 27988 51212 28040 51264
rect 29736 51212 29788 51264
rect 36268 51280 36320 51332
rect 36544 51280 36596 51332
rect 36820 51280 36872 51332
rect 33324 51212 33376 51264
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 1676 51008 1728 51060
rect 8300 51008 8352 51060
rect 20720 51051 20772 51060
rect 20720 51017 20729 51051
rect 20729 51017 20763 51051
rect 20763 51017 20772 51051
rect 20720 51008 20772 51017
rect 22560 51051 22612 51060
rect 22560 51017 22569 51051
rect 22569 51017 22603 51051
rect 22603 51017 22612 51051
rect 22560 51008 22612 51017
rect 23572 51051 23624 51060
rect 23572 51017 23581 51051
rect 23581 51017 23615 51051
rect 23615 51017 23624 51051
rect 23572 51008 23624 51017
rect 25412 51051 25464 51060
rect 25412 51017 25421 51051
rect 25421 51017 25455 51051
rect 25455 51017 25464 51051
rect 25412 51008 25464 51017
rect 27712 51008 27764 51060
rect 31760 51008 31812 51060
rect 32864 51051 32916 51060
rect 32864 51017 32873 51051
rect 32873 51017 32907 51051
rect 32907 51017 32916 51051
rect 32864 51008 32916 51017
rect 36268 51008 36320 51060
rect 37004 51008 37056 51060
rect 38016 51008 38068 51060
rect 7012 50940 7064 50992
rect 22468 50940 22520 50992
rect 23020 50940 23072 50992
rect 24860 50940 24912 50992
rect 1860 50847 1912 50856
rect 1860 50813 1869 50847
rect 1869 50813 1903 50847
rect 1903 50813 1912 50847
rect 1860 50804 1912 50813
rect 4068 50804 4120 50856
rect 21548 50804 21600 50856
rect 26516 50847 26568 50856
rect 26516 50813 26525 50847
rect 26525 50813 26559 50847
rect 26559 50813 26568 50847
rect 26516 50804 26568 50813
rect 34336 50940 34388 50992
rect 35900 50940 35952 50992
rect 28632 50804 28684 50856
rect 35532 50872 35584 50924
rect 36360 50872 36412 50924
rect 37280 50940 37332 50992
rect 37464 50872 37516 50924
rect 36820 50847 36872 50856
rect 36820 50813 36830 50847
rect 36830 50813 36864 50847
rect 36864 50813 36872 50847
rect 36820 50804 36872 50813
rect 38752 50872 38804 50924
rect 38108 50847 38160 50856
rect 4620 50736 4672 50788
rect 18420 50668 18472 50720
rect 23020 50736 23072 50788
rect 26332 50736 26384 50788
rect 26792 50779 26844 50788
rect 26792 50745 26801 50779
rect 26801 50745 26835 50779
rect 26835 50745 26844 50779
rect 26792 50736 26844 50745
rect 27988 50736 28040 50788
rect 32772 50779 32824 50788
rect 32772 50745 32781 50779
rect 32781 50745 32815 50779
rect 32815 50745 32824 50779
rect 32772 50736 32824 50745
rect 36912 50736 36964 50788
rect 38108 50813 38117 50847
rect 38117 50813 38151 50847
rect 38151 50813 38160 50847
rect 38108 50804 38160 50813
rect 27528 50668 27580 50720
rect 27712 50668 27764 50720
rect 37004 50668 37056 50720
rect 37372 50711 37424 50720
rect 37372 50677 37381 50711
rect 37381 50677 37415 50711
rect 37415 50677 37424 50711
rect 37372 50668 37424 50677
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 25320 50507 25372 50516
rect 25320 50473 25329 50507
rect 25329 50473 25363 50507
rect 25363 50473 25372 50507
rect 25320 50464 25372 50473
rect 36912 50464 36964 50516
rect 37004 50464 37056 50516
rect 7288 50371 7340 50380
rect 7288 50337 7297 50371
rect 7297 50337 7331 50371
rect 7331 50337 7340 50371
rect 7288 50328 7340 50337
rect 12256 50328 12308 50380
rect 35808 50328 35860 50380
rect 36912 50371 36964 50380
rect 36912 50337 36919 50371
rect 36919 50337 36964 50371
rect 20996 50260 21048 50312
rect 27988 50260 28040 50312
rect 29920 50260 29972 50312
rect 21088 50192 21140 50244
rect 7472 50167 7524 50176
rect 7472 50133 7481 50167
rect 7481 50133 7515 50167
rect 7515 50133 7524 50167
rect 7472 50124 7524 50133
rect 26516 50192 26568 50244
rect 34520 50192 34572 50244
rect 36912 50328 36964 50337
rect 38660 50328 38712 50380
rect 37556 50260 37608 50312
rect 37464 50192 37516 50244
rect 29368 50124 29420 50176
rect 32588 50124 32640 50176
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 27896 49920 27948 49972
rect 36820 49920 36872 49972
rect 8392 49852 8444 49904
rect 21364 49852 21416 49904
rect 28540 49852 28592 49904
rect 34336 49852 34388 49904
rect 37372 49920 37424 49972
rect 37924 49963 37976 49972
rect 37924 49929 37933 49963
rect 37933 49929 37967 49963
rect 37967 49929 37976 49963
rect 37924 49920 37976 49929
rect 1860 49759 1912 49768
rect 1860 49725 1869 49759
rect 1869 49725 1903 49759
rect 1903 49725 1912 49759
rect 1860 49716 1912 49725
rect 23204 49716 23256 49768
rect 34060 49784 34112 49836
rect 37096 49852 37148 49904
rect 1676 49648 1728 49700
rect 7656 49648 7708 49700
rect 7748 49648 7800 49700
rect 8392 49648 8444 49700
rect 8944 49648 8996 49700
rect 10140 49648 10192 49700
rect 26792 49691 26844 49700
rect 26792 49657 26801 49691
rect 26801 49657 26835 49691
rect 26835 49657 26844 49691
rect 26792 49648 26844 49657
rect 27528 49716 27580 49768
rect 36268 49759 36320 49768
rect 36268 49725 36277 49759
rect 36277 49725 36311 49759
rect 36311 49725 36320 49759
rect 36268 49716 36320 49725
rect 36820 49759 36872 49768
rect 36820 49725 36830 49759
rect 36830 49725 36864 49759
rect 36864 49725 36872 49759
rect 36820 49716 36872 49725
rect 37372 49784 37424 49836
rect 38568 49784 38620 49836
rect 38108 49759 38160 49768
rect 38108 49725 38117 49759
rect 38117 49725 38151 49759
rect 38151 49725 38160 49759
rect 38108 49716 38160 49725
rect 29368 49648 29420 49700
rect 37096 49691 37148 49700
rect 34152 49580 34204 49632
rect 35716 49580 35768 49632
rect 37096 49657 37105 49691
rect 37105 49657 37139 49691
rect 37139 49657 37148 49691
rect 37096 49648 37148 49657
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 8024 49308 8076 49360
rect 1860 49283 1912 49292
rect 1860 49249 1869 49283
rect 1869 49249 1903 49283
rect 1903 49249 1912 49283
rect 1860 49240 1912 49249
rect 24492 49376 24544 49428
rect 35532 49376 35584 49428
rect 37556 49376 37608 49428
rect 27712 49308 27764 49360
rect 35716 49308 35768 49360
rect 25872 49240 25924 49292
rect 35624 49283 35676 49292
rect 35624 49249 35633 49283
rect 35633 49249 35667 49283
rect 35667 49249 35676 49283
rect 35624 49240 35676 49249
rect 35808 49283 35860 49292
rect 35808 49249 35817 49283
rect 35817 49249 35851 49283
rect 35851 49249 35860 49283
rect 35808 49240 35860 49249
rect 36636 49283 36688 49292
rect 2044 49172 2096 49224
rect 22192 49172 22244 49224
rect 23480 49172 23532 49224
rect 36360 49172 36412 49224
rect 8208 49104 8260 49156
rect 35624 49104 35676 49156
rect 36636 49249 36645 49283
rect 36645 49249 36679 49283
rect 36679 49249 36688 49283
rect 36636 49240 36688 49249
rect 37372 49308 37424 49360
rect 37004 49283 37056 49292
rect 37004 49249 37013 49283
rect 37013 49249 37047 49283
rect 37047 49249 37056 49283
rect 37004 49240 37056 49249
rect 39580 49240 39632 49292
rect 36544 49036 36596 49088
rect 37280 49079 37332 49088
rect 37280 49045 37289 49079
rect 37289 49045 37323 49079
rect 37323 49045 37332 49079
rect 37280 49036 37332 49045
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 28908 48832 28960 48884
rect 29460 48832 29512 48884
rect 36912 48832 36964 48884
rect 37740 48832 37792 48884
rect 27712 48764 27764 48816
rect 37280 48764 37332 48816
rect 20076 48696 20128 48748
rect 21272 48696 21324 48748
rect 34612 48696 34664 48748
rect 35164 48696 35216 48748
rect 7288 48628 7340 48680
rect 36268 48628 36320 48680
rect 36452 48628 36504 48680
rect 34612 48560 34664 48612
rect 37372 48696 37424 48748
rect 38844 48628 38896 48680
rect 36912 48603 36964 48612
rect 36912 48569 36921 48603
rect 36921 48569 36955 48603
rect 36955 48569 36964 48603
rect 36912 48560 36964 48569
rect 37004 48603 37056 48612
rect 37004 48569 37013 48603
rect 37013 48569 37047 48603
rect 37047 48569 37056 48603
rect 37004 48560 37056 48569
rect 37740 48560 37792 48612
rect 7380 48535 7432 48544
rect 7380 48501 7389 48535
rect 7389 48501 7423 48535
rect 7423 48501 7432 48535
rect 7380 48492 7432 48501
rect 37096 48492 37148 48544
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 1860 48263 1912 48272
rect 1860 48229 1869 48263
rect 1869 48229 1903 48263
rect 1903 48229 1912 48263
rect 1860 48220 1912 48229
rect 2044 48263 2096 48272
rect 2044 48229 2053 48263
rect 2053 48229 2087 48263
rect 2087 48229 2096 48263
rect 2044 48220 2096 48229
rect 2320 48220 2372 48272
rect 19984 48220 20036 48272
rect 25228 48220 25280 48272
rect 35808 48220 35860 48272
rect 36268 48220 36320 48272
rect 37280 48220 37332 48272
rect 35532 48195 35584 48204
rect 35532 48161 35541 48195
rect 35541 48161 35575 48195
rect 35575 48161 35584 48195
rect 35532 48152 35584 48161
rect 36360 48195 36412 48204
rect 36360 48161 36369 48195
rect 36369 48161 36403 48195
rect 36403 48161 36412 48195
rect 36360 48152 36412 48161
rect 36636 48152 36688 48204
rect 38568 48152 38620 48204
rect 7472 48084 7524 48136
rect 35164 48084 35216 48136
rect 37924 48084 37976 48136
rect 22100 48016 22152 48068
rect 28540 48016 28592 48068
rect 35440 48016 35492 48068
rect 38200 48016 38252 48068
rect 14648 47948 14700 48000
rect 22284 47948 22336 48000
rect 27896 47948 27948 48000
rect 37372 47991 37424 48000
rect 37372 47957 37381 47991
rect 37381 47957 37415 47991
rect 37415 47957 37424 47991
rect 37372 47948 37424 47957
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 27344 47744 27396 47796
rect 35900 47744 35952 47796
rect 2044 47676 2096 47728
rect 23204 47676 23256 47728
rect 26240 47676 26292 47728
rect 36360 47676 36412 47728
rect 36636 47676 36688 47728
rect 37188 47676 37240 47728
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 7472 47608 7524 47660
rect 26608 47608 26660 47660
rect 27068 47608 27120 47660
rect 27344 47608 27396 47660
rect 27896 47608 27948 47660
rect 1400 47583 1452 47592
rect 1400 47549 1409 47583
rect 1409 47549 1443 47583
rect 1443 47549 1452 47583
rect 1400 47540 1452 47549
rect 7012 47540 7064 47592
rect 7288 47540 7340 47592
rect 8392 47583 8444 47592
rect 8392 47549 8401 47583
rect 8401 47549 8435 47583
rect 8435 47549 8444 47583
rect 8392 47540 8444 47549
rect 9772 47540 9824 47592
rect 2596 47472 2648 47524
rect 8208 47472 8260 47524
rect 13268 47472 13320 47524
rect 7288 47447 7340 47456
rect 7288 47413 7297 47447
rect 7297 47413 7331 47447
rect 7331 47413 7340 47447
rect 7288 47404 7340 47413
rect 10232 47404 10284 47456
rect 26424 47540 26476 47592
rect 35808 47540 35860 47592
rect 35992 47540 36044 47592
rect 36636 47540 36688 47592
rect 37280 47540 37332 47592
rect 26516 47515 26568 47524
rect 26516 47481 26525 47515
rect 26525 47481 26559 47515
rect 26559 47481 26568 47515
rect 26516 47472 26568 47481
rect 26608 47515 26660 47524
rect 26608 47481 26617 47515
rect 26617 47481 26651 47515
rect 26651 47481 26660 47515
rect 26608 47472 26660 47481
rect 36268 47472 36320 47524
rect 37188 47472 37240 47524
rect 27896 47404 27948 47456
rect 35992 47404 36044 47456
rect 36360 47404 36412 47456
rect 36452 47404 36504 47456
rect 37464 47404 37516 47456
rect 38108 47447 38160 47456
rect 38108 47413 38117 47447
rect 38117 47413 38151 47447
rect 38151 47413 38160 47447
rect 38108 47404 38160 47413
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 4804 47200 4856 47252
rect 8392 47200 8444 47252
rect 26424 47200 26476 47252
rect 26608 47200 26660 47252
rect 33324 47200 33376 47252
rect 36820 47200 36872 47252
rect 2320 46860 2372 46912
rect 34060 47132 34112 47184
rect 7564 47107 7616 47116
rect 7564 47073 7573 47107
rect 7573 47073 7607 47107
rect 7607 47073 7616 47107
rect 7564 47064 7616 47073
rect 8300 47064 8352 47116
rect 9220 47107 9272 47116
rect 9220 47073 9229 47107
rect 9229 47073 9263 47107
rect 9263 47073 9272 47107
rect 9220 47064 9272 47073
rect 10048 47107 10100 47116
rect 10048 47073 10057 47107
rect 10057 47073 10091 47107
rect 10091 47073 10100 47107
rect 10048 47064 10100 47073
rect 26240 47107 26292 47116
rect 26240 47073 26249 47107
rect 26249 47073 26283 47107
rect 26283 47073 26292 47107
rect 26240 47064 26292 47073
rect 26424 47107 26476 47116
rect 26424 47073 26433 47107
rect 26433 47073 26467 47107
rect 26467 47073 26476 47107
rect 26424 47064 26476 47073
rect 7472 46996 7524 47048
rect 9036 47039 9088 47048
rect 9036 47005 9045 47039
rect 9045 47005 9079 47039
rect 9079 47005 9088 47039
rect 9036 46996 9088 47005
rect 15108 46996 15160 47048
rect 33324 47064 33376 47116
rect 35256 47107 35308 47116
rect 35256 47073 35265 47107
rect 35265 47073 35299 47107
rect 35299 47073 35308 47107
rect 35256 47064 35308 47073
rect 35808 47064 35860 47116
rect 36636 47064 36688 47116
rect 7840 46928 7892 46980
rect 9220 46928 9272 46980
rect 17224 46928 17276 46980
rect 26240 46928 26292 46980
rect 34060 46996 34112 47048
rect 35440 46996 35492 47048
rect 37280 46996 37332 47048
rect 28080 46928 28132 46980
rect 39212 46928 39264 46980
rect 9404 46903 9456 46912
rect 9404 46869 9413 46903
rect 9413 46869 9447 46903
rect 9447 46869 9456 46903
rect 9404 46860 9456 46869
rect 22468 46860 22520 46912
rect 27988 46860 28040 46912
rect 28632 46860 28684 46912
rect 30288 46860 30340 46912
rect 36912 46860 36964 46912
rect 38016 46860 38068 46912
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 28908 46656 28960 46708
rect 35992 46656 36044 46708
rect 1400 46563 1452 46572
rect 1400 46529 1409 46563
rect 1409 46529 1443 46563
rect 1443 46529 1452 46563
rect 1400 46520 1452 46529
rect 4068 46520 4120 46572
rect 2136 46452 2188 46504
rect 15108 46588 15160 46640
rect 9404 46520 9456 46572
rect 17408 46520 17460 46572
rect 30380 46588 30432 46640
rect 36912 46588 36964 46640
rect 37832 46588 37884 46640
rect 7012 46495 7064 46504
rect 7012 46461 7021 46495
rect 7021 46461 7055 46495
rect 7055 46461 7064 46495
rect 7012 46452 7064 46461
rect 7748 46452 7800 46504
rect 8392 46495 8444 46504
rect 8392 46461 8401 46495
rect 8401 46461 8435 46495
rect 8435 46461 8444 46495
rect 8392 46452 8444 46461
rect 9680 46495 9732 46504
rect 9036 46384 9088 46436
rect 9680 46461 9689 46495
rect 9689 46461 9723 46495
rect 9723 46461 9732 46495
rect 9680 46452 9732 46461
rect 28908 46520 28960 46572
rect 29368 46520 29420 46572
rect 26424 46452 26476 46504
rect 27988 46452 28040 46504
rect 36360 46495 36412 46504
rect 36360 46461 36369 46495
rect 36369 46461 36403 46495
rect 36403 46461 36412 46495
rect 36360 46452 36412 46461
rect 37924 46495 37976 46504
rect 37924 46461 37933 46495
rect 37933 46461 37967 46495
rect 37967 46461 37976 46495
rect 37924 46452 37976 46461
rect 26516 46427 26568 46436
rect 26516 46393 26525 46427
rect 26525 46393 26559 46427
rect 26559 46393 26568 46427
rect 26516 46384 26568 46393
rect 26608 46427 26660 46436
rect 26608 46393 26617 46427
rect 26617 46393 26651 46427
rect 26651 46393 26660 46427
rect 26608 46384 26660 46393
rect 35164 46384 35216 46436
rect 37188 46384 37240 46436
rect 7196 46359 7248 46368
rect 7196 46325 7205 46359
rect 7205 46325 7239 46359
rect 7239 46325 7248 46359
rect 7196 46316 7248 46325
rect 8576 46359 8628 46368
rect 8576 46325 8585 46359
rect 8585 46325 8619 46359
rect 8619 46325 8628 46359
rect 8576 46316 8628 46325
rect 9864 46359 9916 46368
rect 9864 46325 9873 46359
rect 9873 46325 9907 46359
rect 9907 46325 9916 46359
rect 9864 46316 9916 46325
rect 26240 46316 26292 46368
rect 30748 46316 30800 46368
rect 31208 46316 31260 46368
rect 37280 46316 37332 46368
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 2780 46112 2832 46164
rect 26424 46112 26476 46164
rect 2044 46087 2096 46096
rect 2044 46053 2053 46087
rect 2053 46053 2087 46087
rect 2087 46053 2096 46087
rect 2044 46044 2096 46053
rect 6276 46044 6328 46096
rect 32864 46112 32916 46164
rect 35716 46112 35768 46164
rect 36728 46112 36780 46164
rect 1860 46019 1912 46028
rect 1860 45985 1869 46019
rect 1869 45985 1903 46019
rect 1903 45985 1912 46019
rect 1860 45976 1912 45985
rect 16304 45976 16356 46028
rect 21364 45976 21416 46028
rect 29920 46044 29972 46096
rect 38292 46112 38344 46164
rect 38660 46112 38712 46164
rect 26424 46019 26476 46028
rect 26424 45985 26433 46019
rect 26433 45985 26467 46019
rect 26467 45985 26476 46019
rect 26424 45976 26476 45985
rect 7748 45908 7800 45960
rect 26240 45840 26292 45892
rect 9312 45815 9364 45824
rect 9312 45781 9321 45815
rect 9321 45781 9355 45815
rect 9355 45781 9364 45815
rect 9312 45772 9364 45781
rect 20720 45772 20772 45824
rect 35716 45976 35768 46028
rect 35808 45976 35860 46028
rect 36544 46019 36596 46028
rect 36544 45985 36553 46019
rect 36553 45985 36587 46019
rect 36587 45985 36596 46019
rect 36544 45976 36596 45985
rect 36728 46019 36780 46028
rect 36728 45985 36735 46019
rect 36735 45985 36780 46019
rect 36728 45976 36780 45985
rect 36912 46019 36964 46028
rect 36912 45985 36921 46019
rect 36921 45985 36955 46019
rect 36955 45985 36964 46019
rect 36912 45976 36964 45985
rect 27344 45840 27396 45892
rect 31116 45840 31168 45892
rect 32680 45840 32732 45892
rect 36084 45840 36136 45892
rect 36360 45840 36412 45892
rect 36544 45840 36596 45892
rect 33968 45772 34020 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 7748 45611 7800 45620
rect 7748 45577 7757 45611
rect 7757 45577 7791 45611
rect 7791 45577 7800 45611
rect 7748 45568 7800 45577
rect 33324 45568 33376 45620
rect 33968 45568 34020 45620
rect 36084 45568 36136 45620
rect 12440 45500 12492 45552
rect 17684 45500 17736 45552
rect 7380 45432 7432 45484
rect 18696 45432 18748 45484
rect 21732 45432 21784 45484
rect 7288 45364 7340 45416
rect 9404 45364 9456 45416
rect 9496 45407 9548 45416
rect 9496 45373 9505 45407
rect 9505 45373 9539 45407
rect 9539 45373 9548 45407
rect 9496 45364 9548 45373
rect 9956 45364 10008 45416
rect 26424 45364 26476 45416
rect 28540 45500 28592 45552
rect 35716 45500 35768 45552
rect 36268 45500 36320 45552
rect 28540 45364 28592 45416
rect 35808 45407 35860 45416
rect 35808 45373 35817 45407
rect 35817 45373 35851 45407
rect 35851 45373 35860 45407
rect 35808 45364 35860 45373
rect 37188 45568 37240 45620
rect 36544 45500 36596 45552
rect 36820 45432 36872 45484
rect 37188 45432 37240 45484
rect 37740 45568 37792 45620
rect 38292 45568 38344 45620
rect 17500 45296 17552 45348
rect 21732 45296 21784 45348
rect 26516 45339 26568 45348
rect 26516 45305 26525 45339
rect 26525 45305 26559 45339
rect 26559 45305 26568 45339
rect 26516 45296 26568 45305
rect 8668 45228 8720 45280
rect 15844 45228 15896 45280
rect 26240 45228 26292 45280
rect 27436 45296 27488 45348
rect 31576 45296 31628 45348
rect 36268 45296 36320 45348
rect 36820 45339 36872 45348
rect 36820 45305 36829 45339
rect 36829 45305 36863 45339
rect 36863 45305 36872 45339
rect 36820 45296 36872 45305
rect 38200 45364 38252 45416
rect 39396 45364 39448 45416
rect 37740 45228 37792 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 6368 45024 6420 45076
rect 1860 44999 1912 45008
rect 1860 44965 1869 44999
rect 1869 44965 1903 44999
rect 1903 44965 1912 44999
rect 1860 44956 1912 44965
rect 2320 44956 2372 45008
rect 3516 44956 3568 45008
rect 2228 44888 2280 44940
rect 23480 45024 23532 45076
rect 24400 45024 24452 45076
rect 27436 45024 27488 45076
rect 28816 45024 28868 45076
rect 29092 45024 29144 45076
rect 29736 45024 29788 45076
rect 34520 45024 34572 45076
rect 37740 45024 37792 45076
rect 27528 44956 27580 45008
rect 29000 44956 29052 45008
rect 10508 44931 10560 44940
rect 10508 44897 10517 44931
rect 10517 44897 10551 44931
rect 10551 44897 10560 44931
rect 10508 44888 10560 44897
rect 11152 44888 11204 44940
rect 23020 44888 23072 44940
rect 24032 44931 24084 44940
rect 24032 44897 24041 44931
rect 24041 44897 24075 44931
rect 24075 44897 24084 44931
rect 24032 44888 24084 44897
rect 26608 44888 26660 44940
rect 30012 44956 30064 45008
rect 36084 44956 36136 45008
rect 9496 44863 9548 44872
rect 9496 44829 9505 44863
rect 9505 44829 9539 44863
rect 9539 44829 9548 44863
rect 9496 44820 9548 44829
rect 22192 44820 22244 44872
rect 24492 44820 24544 44872
rect 30288 44888 30340 44940
rect 34520 44931 34572 44940
rect 34520 44897 34529 44931
rect 34529 44897 34563 44931
rect 34563 44897 34572 44931
rect 34520 44888 34572 44897
rect 29184 44820 29236 44872
rect 35256 44888 35308 44940
rect 35808 44931 35860 44940
rect 35808 44897 35817 44931
rect 35817 44897 35851 44931
rect 35851 44897 35860 44931
rect 35808 44888 35860 44897
rect 35716 44820 35768 44872
rect 36084 44820 36136 44872
rect 11888 44752 11940 44804
rect 28816 44752 28868 44804
rect 8116 44684 8168 44736
rect 9036 44727 9088 44736
rect 9036 44693 9045 44727
rect 9045 44693 9079 44727
rect 9079 44693 9088 44727
rect 9036 44684 9088 44693
rect 10692 44727 10744 44736
rect 10692 44693 10701 44727
rect 10701 44693 10735 44727
rect 10735 44693 10744 44727
rect 10692 44684 10744 44693
rect 27528 44684 27580 44736
rect 29552 44727 29604 44736
rect 29552 44693 29561 44727
rect 29561 44693 29595 44727
rect 29595 44693 29604 44727
rect 29552 44684 29604 44693
rect 30196 44752 30248 44804
rect 35992 44727 36044 44736
rect 35992 44693 36001 44727
rect 36001 44693 36035 44727
rect 36035 44693 36044 44727
rect 35992 44684 36044 44693
rect 36544 44752 36596 44804
rect 36820 44931 36872 44940
rect 36820 44897 36829 44931
rect 36829 44897 36863 44931
rect 36863 44897 36872 44931
rect 36820 44888 36872 44897
rect 38016 44888 38068 44940
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 15108 44480 15160 44532
rect 26424 44480 26476 44532
rect 26792 44480 26844 44532
rect 2136 44412 2188 44464
rect 32956 44480 33008 44532
rect 34612 44523 34664 44532
rect 34612 44489 34621 44523
rect 34621 44489 34655 44523
rect 34655 44489 34664 44523
rect 34612 44480 34664 44489
rect 37188 44480 37240 44532
rect 36452 44412 36504 44464
rect 36912 44412 36964 44464
rect 6552 44344 6604 44396
rect 1860 44319 1912 44328
rect 1860 44285 1869 44319
rect 1869 44285 1903 44319
rect 1903 44285 1912 44319
rect 1860 44276 1912 44285
rect 7380 44319 7432 44328
rect 7380 44285 7389 44319
rect 7389 44285 7423 44319
rect 7423 44285 7432 44319
rect 7380 44276 7432 44285
rect 9864 44344 9916 44396
rect 17592 44344 17644 44396
rect 19248 44344 19300 44396
rect 33324 44344 33376 44396
rect 8208 44319 8260 44328
rect 8208 44285 8217 44319
rect 8217 44285 8251 44319
rect 8251 44285 8260 44319
rect 8208 44276 8260 44285
rect 8760 44276 8812 44328
rect 10140 44276 10192 44328
rect 22284 44276 22336 44328
rect 13452 44208 13504 44260
rect 26792 44208 26844 44260
rect 29184 44208 29236 44260
rect 1768 44140 1820 44192
rect 5540 44140 5592 44192
rect 7748 44183 7800 44192
rect 7748 44149 7757 44183
rect 7757 44149 7791 44183
rect 7791 44149 7800 44183
rect 7748 44140 7800 44149
rect 9864 44183 9916 44192
rect 9864 44149 9873 44183
rect 9873 44149 9907 44183
rect 9907 44149 9916 44183
rect 9864 44140 9916 44149
rect 27988 44140 28040 44192
rect 29000 44140 29052 44192
rect 30288 44276 30340 44328
rect 35348 44276 35400 44328
rect 37188 44344 37240 44396
rect 30656 44208 30708 44260
rect 35716 44208 35768 44260
rect 35992 44208 36044 44260
rect 31300 44140 31352 44192
rect 35900 44140 35952 44192
rect 36544 44140 36596 44192
rect 36820 44251 36872 44260
rect 36820 44217 36829 44251
rect 36829 44217 36863 44251
rect 36863 44217 36872 44251
rect 36820 44208 36872 44217
rect 37372 44140 37424 44192
rect 37740 44319 37792 44328
rect 37740 44285 37749 44319
rect 37749 44285 37783 44319
rect 37783 44285 37792 44319
rect 37740 44276 37792 44285
rect 38752 44276 38804 44328
rect 37832 44251 37884 44260
rect 37832 44217 37841 44251
rect 37841 44217 37875 44251
rect 37875 44217 37884 44251
rect 37832 44208 37884 44217
rect 38476 44140 38528 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 1952 43936 2004 43988
rect 9496 43936 9548 43988
rect 34152 43936 34204 43988
rect 34336 43936 34388 43988
rect 35900 43936 35952 43988
rect 9588 43868 9640 43920
rect 22008 43868 22060 43920
rect 35348 43868 35400 43920
rect 36544 43936 36596 43988
rect 8208 43843 8260 43852
rect 8208 43809 8217 43843
rect 8217 43809 8251 43843
rect 8251 43809 8260 43843
rect 8208 43800 8260 43809
rect 8484 43800 8536 43852
rect 7288 43732 7340 43784
rect 29184 43800 29236 43852
rect 30288 43800 30340 43852
rect 30380 43800 30432 43852
rect 31300 43800 31352 43852
rect 35072 43843 35124 43852
rect 35072 43809 35081 43843
rect 35081 43809 35115 43843
rect 35115 43809 35124 43843
rect 35072 43800 35124 43809
rect 35808 43800 35860 43852
rect 8208 43664 8260 43716
rect 31484 43732 31536 43784
rect 31116 43664 31168 43716
rect 36544 43843 36596 43852
rect 36544 43809 36551 43843
rect 36551 43809 36596 43843
rect 36544 43800 36596 43809
rect 37188 43936 37240 43988
rect 37556 43936 37608 43988
rect 38108 43868 38160 43920
rect 37556 43732 37608 43784
rect 37280 43664 37332 43716
rect 8576 43639 8628 43648
rect 8576 43605 8585 43639
rect 8585 43605 8619 43639
rect 8619 43605 8628 43639
rect 8576 43596 8628 43605
rect 30380 43596 30432 43648
rect 39028 43596 39080 43648
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 2044 43392 2096 43444
rect 20720 43392 20772 43444
rect 28632 43392 28684 43444
rect 36728 43392 36780 43444
rect 37004 43392 37056 43444
rect 26516 43324 26568 43376
rect 27344 43324 27396 43376
rect 34520 43324 34572 43376
rect 36544 43324 36596 43376
rect 2688 43256 2740 43308
rect 19156 43256 19208 43308
rect 1860 43231 1912 43240
rect 1860 43197 1869 43231
rect 1869 43197 1903 43231
rect 1903 43197 1912 43231
rect 1860 43188 1912 43197
rect 2136 43188 2188 43240
rect 26516 43231 26568 43240
rect 26516 43197 26525 43231
rect 26525 43197 26559 43231
rect 26559 43197 26568 43231
rect 26516 43188 26568 43197
rect 28080 43188 28132 43240
rect 25872 43052 25924 43104
rect 27528 43120 27580 43172
rect 27988 43052 28040 43104
rect 28908 43095 28960 43104
rect 28908 43061 28917 43095
rect 28917 43061 28951 43095
rect 28951 43061 28960 43095
rect 28908 43052 28960 43061
rect 29460 43188 29512 43240
rect 30012 43188 30064 43240
rect 30288 43188 30340 43240
rect 34980 43188 35032 43240
rect 35440 43188 35492 43240
rect 32496 43120 32548 43172
rect 34612 43120 34664 43172
rect 37464 43188 37516 43240
rect 37740 43231 37792 43240
rect 37740 43197 37749 43231
rect 37749 43197 37783 43231
rect 37783 43197 37792 43231
rect 37740 43188 37792 43197
rect 39028 43188 39080 43240
rect 37096 43120 37148 43172
rect 37832 43163 37884 43172
rect 37832 43129 37841 43163
rect 37841 43129 37875 43163
rect 37875 43129 37884 43163
rect 37832 43120 37884 43129
rect 33048 43052 33100 43104
rect 37188 43052 37240 43104
rect 38108 43095 38160 43104
rect 38108 43061 38117 43095
rect 38117 43061 38151 43095
rect 38151 43061 38160 43095
rect 38108 43052 38160 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 8484 42848 8536 42900
rect 16028 42848 16080 42900
rect 27344 42848 27396 42900
rect 34152 42848 34204 42900
rect 35348 42848 35400 42900
rect 9036 42780 9088 42832
rect 14740 42780 14792 42832
rect 25872 42780 25924 42832
rect 27528 42780 27580 42832
rect 29276 42780 29328 42832
rect 1860 42755 1912 42764
rect 1860 42721 1869 42755
rect 1869 42721 1903 42755
rect 1903 42721 1912 42755
rect 1860 42712 1912 42721
rect 2044 42755 2096 42764
rect 2044 42721 2053 42755
rect 2053 42721 2087 42755
rect 2087 42721 2096 42755
rect 2044 42712 2096 42721
rect 26516 42644 26568 42696
rect 2044 42576 2096 42628
rect 27068 42712 27120 42764
rect 30288 42712 30340 42764
rect 35348 42712 35400 42764
rect 27344 42644 27396 42696
rect 29276 42644 29328 42696
rect 35716 42755 35768 42764
rect 35716 42721 35725 42755
rect 35725 42721 35759 42755
rect 35759 42721 35768 42755
rect 35716 42712 35768 42721
rect 27896 42576 27948 42628
rect 35624 42576 35676 42628
rect 35716 42576 35768 42628
rect 36360 42712 36412 42764
rect 37740 42848 37792 42900
rect 21916 42508 21968 42560
rect 36728 42576 36780 42628
rect 36820 42576 36872 42628
rect 37832 42780 37884 42832
rect 37280 42712 37332 42764
rect 36544 42508 36596 42560
rect 37280 42508 37332 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 26240 42304 26292 42356
rect 27068 42304 27120 42356
rect 26792 42236 26844 42288
rect 3608 42100 3660 42152
rect 7196 42100 7248 42152
rect 7932 42143 7984 42152
rect 7932 42109 7941 42143
rect 7941 42109 7975 42143
rect 7975 42109 7984 42143
rect 7932 42100 7984 42109
rect 26240 42168 26292 42220
rect 26608 42168 26660 42220
rect 26424 42100 26476 42152
rect 8576 42032 8628 42084
rect 10324 42032 10376 42084
rect 27344 42236 27396 42288
rect 28448 42304 28500 42356
rect 36268 42304 36320 42356
rect 27528 42168 27580 42220
rect 27528 42032 27580 42084
rect 14556 41964 14608 42016
rect 26516 41964 26568 42016
rect 26792 41964 26844 42016
rect 27988 42143 28040 42152
rect 27988 42109 27997 42143
rect 27997 42109 28031 42143
rect 28031 42109 28040 42143
rect 27988 42100 28040 42109
rect 31576 42236 31628 42288
rect 33048 42236 33100 42288
rect 37372 42304 37424 42356
rect 33324 42168 33376 42220
rect 28540 42100 28592 42152
rect 28816 42100 28868 42152
rect 29092 42100 29144 42152
rect 34796 42143 34848 42152
rect 34796 42109 34805 42143
rect 34805 42109 34839 42143
rect 34839 42109 34848 42143
rect 34796 42100 34848 42109
rect 36176 42100 36228 42152
rect 37464 42236 37516 42288
rect 37740 42236 37792 42288
rect 36820 42168 36872 42220
rect 38200 42168 38252 42220
rect 38476 42168 38528 42220
rect 37372 42100 37424 42152
rect 37740 42100 37792 42152
rect 38200 42032 38252 42084
rect 28816 41964 28868 42016
rect 36268 41964 36320 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 2780 41760 2832 41812
rect 27344 41760 27396 41812
rect 1860 41735 1912 41744
rect 1860 41701 1869 41735
rect 1869 41701 1903 41735
rect 1903 41701 1912 41735
rect 1860 41692 1912 41701
rect 5540 41692 5592 41744
rect 5080 41624 5132 41676
rect 9496 41692 9548 41744
rect 22100 41692 22152 41744
rect 25872 41692 25924 41744
rect 26424 41735 26476 41744
rect 26424 41701 26433 41735
rect 26433 41701 26467 41735
rect 26467 41701 26476 41735
rect 26424 41692 26476 41701
rect 20076 41624 20128 41676
rect 7932 41599 7984 41608
rect 7932 41565 7941 41599
rect 7941 41565 7975 41599
rect 7975 41565 7984 41599
rect 7932 41556 7984 41565
rect 8300 41463 8352 41472
rect 8300 41429 8309 41463
rect 8309 41429 8343 41463
rect 8343 41429 8352 41463
rect 8300 41420 8352 41429
rect 15108 41556 15160 41608
rect 26516 41667 26568 41676
rect 26516 41633 26525 41667
rect 26525 41633 26559 41667
rect 26559 41633 26568 41667
rect 26516 41624 26568 41633
rect 26608 41667 26660 41676
rect 26608 41633 26622 41667
rect 26622 41633 26656 41667
rect 26656 41633 26660 41667
rect 26608 41624 26660 41633
rect 31116 41760 31168 41812
rect 34612 41803 34664 41812
rect 34612 41769 34621 41803
rect 34621 41769 34655 41803
rect 34655 41769 34664 41803
rect 34612 41760 34664 41769
rect 35900 41760 35952 41812
rect 37556 41760 37608 41812
rect 27712 41692 27764 41744
rect 27988 41692 28040 41744
rect 28632 41692 28684 41744
rect 29092 41692 29144 41744
rect 37096 41692 37148 41744
rect 29736 41624 29788 41676
rect 34796 41667 34848 41676
rect 34796 41633 34805 41667
rect 34805 41633 34839 41667
rect 34839 41633 34848 41667
rect 34796 41624 34848 41633
rect 35808 41624 35860 41676
rect 35900 41624 35952 41676
rect 36728 41667 36780 41676
rect 36728 41633 36737 41667
rect 36737 41633 36771 41667
rect 36771 41633 36780 41667
rect 36728 41624 36780 41633
rect 37004 41624 37056 41676
rect 37832 41624 37884 41676
rect 9128 41463 9180 41472
rect 9128 41429 9137 41463
rect 9137 41429 9171 41463
rect 9171 41429 9180 41463
rect 9128 41420 9180 41429
rect 20168 41420 20220 41472
rect 29092 41556 29144 41608
rect 34888 41556 34940 41608
rect 35348 41556 35400 41608
rect 35532 41556 35584 41608
rect 36820 41556 36872 41608
rect 27160 41488 27212 41540
rect 27896 41488 27948 41540
rect 35256 41488 35308 41540
rect 35808 41488 35860 41540
rect 27528 41420 27580 41472
rect 29184 41420 29236 41472
rect 29920 41420 29972 41472
rect 30288 41420 30340 41472
rect 32588 41420 32640 41472
rect 34796 41420 34848 41472
rect 35532 41420 35584 41472
rect 37372 41420 37424 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 22836 41216 22888 41268
rect 2136 41148 2188 41200
rect 23112 41148 23164 41200
rect 27436 41216 27488 41268
rect 34060 41216 34112 41268
rect 38108 41216 38160 41268
rect 6460 41080 6512 41132
rect 1860 41055 1912 41064
rect 1860 41021 1869 41055
rect 1869 41021 1903 41055
rect 1903 41021 1912 41055
rect 1860 41012 1912 41021
rect 7932 41055 7984 41064
rect 7932 41021 7941 41055
rect 7941 41021 7975 41055
rect 7975 41021 7984 41055
rect 7932 41012 7984 41021
rect 8208 41080 8260 41132
rect 36728 41148 36780 41200
rect 37372 41148 37424 41200
rect 9588 41012 9640 41064
rect 10968 40944 11020 40996
rect 22376 41012 22428 41064
rect 23112 41012 23164 41064
rect 26516 41055 26568 41064
rect 26516 41021 26525 41055
rect 26525 41021 26559 41055
rect 26559 41021 26568 41055
rect 26516 41012 26568 41021
rect 34612 41055 34664 41064
rect 34612 41021 34621 41055
rect 34621 41021 34655 41055
rect 34655 41021 34664 41055
rect 34612 41012 34664 41021
rect 36636 41080 36688 41132
rect 26424 40944 26476 40996
rect 26792 40987 26844 40996
rect 26792 40953 26801 40987
rect 26801 40953 26835 40987
rect 26835 40953 26844 40987
rect 26792 40944 26844 40953
rect 29092 40944 29144 40996
rect 30748 40944 30800 40996
rect 31576 40944 31628 40996
rect 34152 40944 34204 40996
rect 34796 40944 34848 40996
rect 35348 40944 35400 40996
rect 37372 41012 37424 41064
rect 37556 41055 37608 41064
rect 37556 41021 37565 41055
rect 37565 41021 37599 41055
rect 37599 41021 37608 41055
rect 37556 41012 37608 41021
rect 38844 41012 38896 41064
rect 36544 40987 36596 40996
rect 36544 40953 36553 40987
rect 36553 40953 36587 40987
rect 36587 40953 36596 40987
rect 36544 40944 36596 40953
rect 36636 40987 36688 40996
rect 36636 40953 36645 40987
rect 36645 40953 36679 40987
rect 36679 40953 36688 40987
rect 36636 40944 36688 40953
rect 37464 40944 37516 40996
rect 7472 40876 7524 40928
rect 9956 40876 10008 40928
rect 27896 40876 27948 40928
rect 34336 40876 34388 40928
rect 35440 40876 35492 40928
rect 36912 40919 36964 40928
rect 36912 40885 36921 40919
rect 36921 40885 36955 40919
rect 36955 40885 36964 40919
rect 36912 40876 36964 40885
rect 37096 40876 37148 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 1584 40672 1636 40724
rect 24860 40715 24912 40724
rect 4896 40604 4948 40656
rect 8208 40536 8260 40588
rect 24860 40681 24869 40715
rect 24869 40681 24903 40715
rect 24903 40681 24912 40715
rect 24860 40672 24912 40681
rect 26516 40672 26568 40724
rect 34060 40672 34112 40724
rect 24308 40604 24360 40656
rect 29000 40647 29052 40656
rect 29000 40613 29034 40647
rect 29034 40613 29052 40647
rect 29000 40604 29052 40613
rect 24676 40579 24728 40588
rect 7932 40468 7984 40520
rect 24676 40545 24685 40579
rect 24685 40545 24719 40579
rect 24719 40545 24728 40579
rect 24676 40536 24728 40545
rect 26516 40536 26568 40588
rect 28816 40536 28868 40588
rect 29276 40536 29328 40588
rect 30012 40536 30064 40588
rect 35164 40579 35216 40588
rect 35164 40545 35173 40579
rect 35173 40545 35207 40579
rect 35207 40545 35216 40579
rect 35164 40536 35216 40545
rect 35808 40579 35860 40588
rect 35808 40545 35817 40579
rect 35817 40545 35851 40579
rect 35851 40545 35860 40579
rect 35808 40536 35860 40545
rect 22836 40511 22888 40520
rect 22836 40477 22845 40511
rect 22845 40477 22879 40511
rect 22879 40477 22888 40511
rect 22836 40468 22888 40477
rect 23020 40468 23072 40520
rect 8576 40400 8628 40452
rect 21548 40400 21600 40452
rect 7932 40332 7984 40384
rect 8116 40332 8168 40384
rect 13544 40332 13596 40384
rect 21364 40332 21416 40384
rect 27436 40468 27488 40520
rect 34888 40468 34940 40520
rect 35440 40468 35492 40520
rect 37004 40672 37056 40724
rect 36544 40647 36596 40656
rect 36544 40613 36553 40647
rect 36553 40613 36587 40647
rect 36587 40613 36596 40647
rect 36544 40604 36596 40613
rect 36360 40579 36412 40588
rect 36360 40545 36370 40579
rect 36370 40545 36404 40579
rect 36404 40545 36412 40579
rect 36636 40579 36688 40588
rect 36360 40536 36412 40545
rect 36636 40545 36645 40579
rect 36645 40545 36679 40579
rect 36679 40545 36688 40579
rect 36636 40536 36688 40545
rect 36728 40579 36780 40588
rect 36728 40545 36742 40579
rect 36742 40545 36776 40579
rect 36776 40545 36780 40579
rect 36728 40536 36780 40545
rect 38568 40468 38620 40520
rect 29736 40400 29788 40452
rect 33968 40400 34020 40452
rect 36084 40400 36136 40452
rect 30656 40332 30708 40384
rect 32956 40332 33008 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 20260 40128 20312 40180
rect 37556 40128 37608 40180
rect 37832 40128 37884 40180
rect 38568 40128 38620 40180
rect 26792 40060 26844 40112
rect 27804 40060 27856 40112
rect 29276 40060 29328 40112
rect 32220 40060 32272 40112
rect 2044 40035 2096 40044
rect 2044 40001 2053 40035
rect 2053 40001 2087 40035
rect 2087 40001 2096 40035
rect 2044 39992 2096 40001
rect 8024 40035 8076 40044
rect 8024 40001 8033 40035
rect 8033 40001 8067 40035
rect 8067 40001 8076 40035
rect 8024 39992 8076 40001
rect 9864 39992 9916 40044
rect 11704 39992 11756 40044
rect 17316 39992 17368 40044
rect 22468 39992 22520 40044
rect 1860 39967 1912 39976
rect 1860 39933 1869 39967
rect 1869 39933 1903 39967
rect 1903 39933 1912 39967
rect 1860 39924 1912 39933
rect 7932 39924 7984 39976
rect 27436 39924 27488 39976
rect 27804 39924 27856 39976
rect 29552 39924 29604 39976
rect 28816 39856 28868 39908
rect 32680 39992 32732 40044
rect 35716 39992 35768 40044
rect 34612 39967 34664 39976
rect 34612 39933 34621 39967
rect 34621 39933 34655 39967
rect 34655 39933 34664 39967
rect 34612 39924 34664 39933
rect 32220 39856 32272 39908
rect 36084 39924 36136 39976
rect 36544 39967 36596 39976
rect 35808 39856 35860 39908
rect 36544 39933 36553 39967
rect 36553 39933 36587 39967
rect 36587 39933 36596 39967
rect 36544 39924 36596 39933
rect 37280 39992 37332 40044
rect 38292 39992 38344 40044
rect 37740 39967 37792 39976
rect 36636 39899 36688 39908
rect 36636 39865 36645 39899
rect 36645 39865 36679 39899
rect 36679 39865 36688 39899
rect 36636 39856 36688 39865
rect 37740 39933 37749 39967
rect 37749 39933 37783 39967
rect 37783 39933 37792 39967
rect 37740 39924 37792 39933
rect 38108 39924 38160 39976
rect 8392 39831 8444 39840
rect 8392 39797 8401 39831
rect 8401 39797 8435 39831
rect 8435 39797 8444 39831
rect 8392 39788 8444 39797
rect 29552 39788 29604 39840
rect 31300 39788 31352 39840
rect 34888 39788 34940 39840
rect 38016 39856 38068 39908
rect 36912 39831 36964 39840
rect 36912 39797 36921 39831
rect 36921 39797 36955 39831
rect 36955 39797 36964 39831
rect 36912 39788 36964 39797
rect 37556 39788 37608 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 2688 39584 2740 39636
rect 18972 39584 19024 39636
rect 34888 39584 34940 39636
rect 35532 39584 35584 39636
rect 2136 39516 2188 39568
rect 10968 39516 11020 39568
rect 28908 39516 28960 39568
rect 29552 39516 29604 39568
rect 30196 39516 30248 39568
rect 30380 39559 30432 39568
rect 30380 39525 30414 39559
rect 30414 39525 30432 39559
rect 30380 39516 30432 39525
rect 31300 39516 31352 39568
rect 32312 39516 32364 39568
rect 32680 39516 32732 39568
rect 36084 39516 36136 39568
rect 1860 39491 1912 39500
rect 1860 39457 1869 39491
rect 1869 39457 1903 39491
rect 1903 39457 1912 39491
rect 1860 39448 1912 39457
rect 8208 39448 8260 39500
rect 17500 39448 17552 39500
rect 2044 39380 2096 39432
rect 9496 39380 9548 39432
rect 9220 39312 9272 39364
rect 16856 39380 16908 39432
rect 27804 39380 27856 39432
rect 34520 39448 34572 39500
rect 35532 39448 35584 39500
rect 35900 39448 35952 39500
rect 36268 39491 36320 39500
rect 36268 39457 36277 39491
rect 36277 39457 36311 39491
rect 36311 39457 36320 39491
rect 36268 39448 36320 39457
rect 36728 39584 36780 39636
rect 36544 39559 36596 39568
rect 36544 39525 36553 39559
rect 36553 39525 36587 39559
rect 36587 39525 36596 39559
rect 36544 39516 36596 39525
rect 36636 39491 36688 39500
rect 36636 39457 36645 39491
rect 36645 39457 36679 39491
rect 36679 39457 36688 39491
rect 36636 39448 36688 39457
rect 35256 39380 35308 39432
rect 12348 39312 12400 39364
rect 22560 39312 22612 39364
rect 23388 39312 23440 39364
rect 24032 39312 24084 39364
rect 31484 39355 31536 39364
rect 31484 39321 31493 39355
rect 31493 39321 31527 39355
rect 31527 39321 31536 39355
rect 31484 39312 31536 39321
rect 35992 39312 36044 39364
rect 36084 39312 36136 39364
rect 23296 39244 23348 39296
rect 28908 39244 28960 39296
rect 29552 39287 29604 39296
rect 29552 39253 29561 39287
rect 29561 39253 29595 39287
rect 29595 39253 29604 39287
rect 29552 39244 29604 39253
rect 36268 39244 36320 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 22836 39040 22888 39092
rect 25412 39040 25464 39092
rect 30564 39040 30616 39092
rect 31484 39040 31536 39092
rect 32864 39040 32916 39092
rect 35532 39040 35584 39092
rect 35992 39040 36044 39092
rect 28080 38972 28132 39024
rect 35256 38972 35308 39024
rect 36084 38972 36136 39024
rect 6276 38904 6328 38956
rect 17684 38836 17736 38888
rect 21824 38879 21876 38888
rect 21824 38845 21831 38879
rect 21831 38845 21876 38879
rect 21824 38836 21876 38845
rect 23020 38879 23072 38888
rect 23020 38845 23029 38879
rect 23029 38845 23063 38879
rect 23063 38845 23072 38879
rect 23020 38836 23072 38845
rect 21916 38811 21968 38820
rect 21916 38777 21925 38811
rect 21925 38777 21959 38811
rect 21959 38777 21968 38811
rect 21916 38768 21968 38777
rect 23480 38904 23532 38956
rect 24032 38904 24084 38956
rect 36544 38904 36596 38956
rect 24308 38836 24360 38888
rect 25228 38879 25280 38888
rect 25228 38845 25237 38879
rect 25237 38845 25271 38879
rect 25271 38845 25280 38879
rect 25228 38836 25280 38845
rect 24400 38768 24452 38820
rect 25504 38836 25556 38888
rect 28632 38879 28684 38888
rect 28632 38845 28641 38879
rect 28641 38845 28675 38879
rect 28675 38845 28684 38879
rect 28632 38836 28684 38845
rect 29092 38836 29144 38888
rect 34796 38836 34848 38888
rect 37096 39040 37148 39092
rect 37280 38904 37332 38956
rect 34520 38768 34572 38820
rect 35256 38768 35308 38820
rect 35532 38768 35584 38820
rect 36636 38811 36688 38820
rect 36636 38777 36645 38811
rect 36645 38777 36679 38811
rect 36679 38777 36688 38811
rect 37464 38836 37516 38888
rect 38108 39040 38160 39092
rect 38016 38972 38068 39024
rect 37740 38811 37792 38820
rect 36636 38768 36688 38777
rect 37740 38777 37749 38811
rect 37749 38777 37783 38811
rect 37783 38777 37792 38811
rect 37740 38768 37792 38777
rect 24032 38700 24084 38752
rect 25320 38743 25372 38752
rect 25320 38709 25329 38743
rect 25329 38709 25363 38743
rect 25363 38709 25372 38743
rect 25320 38700 25372 38709
rect 25504 38700 25556 38752
rect 30380 38700 30432 38752
rect 31944 38700 31996 38752
rect 37096 38700 37148 38752
rect 37280 38700 37332 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 22100 38496 22152 38548
rect 22744 38496 22796 38548
rect 1860 38471 1912 38480
rect 1860 38437 1869 38471
rect 1869 38437 1903 38471
rect 1903 38437 1912 38471
rect 1860 38428 1912 38437
rect 2044 38471 2096 38480
rect 2044 38437 2053 38471
rect 2053 38437 2087 38471
rect 2087 38437 2096 38471
rect 2044 38428 2096 38437
rect 17776 38428 17828 38480
rect 22284 38428 22336 38480
rect 22008 38360 22060 38412
rect 23388 38496 23440 38548
rect 23480 38428 23532 38480
rect 25320 38428 25372 38480
rect 26424 38471 26476 38480
rect 26424 38437 26433 38471
rect 26433 38437 26467 38471
rect 26467 38437 26476 38471
rect 26424 38428 26476 38437
rect 22560 38403 22612 38412
rect 22560 38369 22569 38403
rect 22569 38369 22603 38403
rect 22603 38369 22612 38403
rect 22560 38360 22612 38369
rect 6368 38292 6420 38344
rect 22284 38292 22336 38344
rect 23204 38360 23256 38412
rect 23388 38360 23440 38412
rect 24492 38360 24544 38412
rect 25872 38360 25924 38412
rect 26516 38403 26568 38412
rect 26516 38369 26525 38403
rect 26525 38369 26559 38403
rect 26559 38369 26568 38403
rect 26516 38360 26568 38369
rect 27344 38428 27396 38480
rect 31484 38428 31536 38480
rect 34612 38496 34664 38548
rect 35624 38496 35676 38548
rect 23296 38292 23348 38344
rect 27896 38360 27948 38412
rect 28816 38360 28868 38412
rect 29276 38360 29328 38412
rect 29460 38360 29512 38412
rect 35348 38360 35400 38412
rect 35716 38360 35768 38412
rect 35992 38360 36044 38412
rect 36544 38360 36596 38412
rect 36728 38360 36780 38412
rect 36912 38360 36964 38412
rect 38016 38496 38068 38548
rect 1584 38224 1636 38276
rect 22744 38224 22796 38276
rect 23388 38224 23440 38276
rect 29184 38335 29236 38344
rect 29184 38301 29193 38335
rect 29193 38301 29227 38335
rect 29227 38301 29236 38335
rect 29184 38292 29236 38301
rect 35532 38292 35584 38344
rect 26332 38224 26384 38276
rect 29736 38224 29788 38276
rect 34612 38224 34664 38276
rect 34980 38224 35032 38276
rect 35992 38224 36044 38276
rect 37372 38292 37424 38344
rect 25228 38199 25280 38208
rect 25228 38165 25237 38199
rect 25237 38165 25271 38199
rect 25271 38165 25280 38199
rect 25228 38156 25280 38165
rect 25320 38156 25372 38208
rect 27160 38156 27212 38208
rect 27896 38156 27948 38208
rect 36636 38156 36688 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 2504 37952 2556 38004
rect 26608 37952 26660 38004
rect 26792 37995 26844 38004
rect 26792 37961 26801 37995
rect 26801 37961 26835 37995
rect 26835 37961 26844 37995
rect 26792 37952 26844 37961
rect 28448 37952 28500 38004
rect 2136 37884 2188 37936
rect 1676 37816 1728 37868
rect 21916 37884 21968 37936
rect 18052 37816 18104 37868
rect 21732 37791 21784 37800
rect 21732 37757 21741 37791
rect 21741 37757 21775 37791
rect 21775 37757 21784 37791
rect 21732 37748 21784 37757
rect 21916 37791 21968 37800
rect 21916 37757 21923 37791
rect 21923 37757 21968 37791
rect 21916 37748 21968 37757
rect 22284 37816 22336 37868
rect 24216 37884 24268 37936
rect 22376 37748 22428 37800
rect 22468 37748 22520 37800
rect 25320 37816 25372 37868
rect 23296 37791 23348 37800
rect 23296 37757 23310 37791
rect 23310 37757 23344 37791
rect 23344 37757 23348 37791
rect 23296 37748 23348 37757
rect 23480 37748 23532 37800
rect 24400 37748 24452 37800
rect 26332 37816 26384 37868
rect 26516 37791 26568 37800
rect 26516 37757 26525 37791
rect 26525 37757 26559 37791
rect 26559 37757 26568 37791
rect 26516 37748 26568 37757
rect 28632 37884 28684 37936
rect 28448 37816 28500 37868
rect 30380 37884 30432 37936
rect 28264 37748 28316 37800
rect 28632 37748 28684 37800
rect 29276 37816 29328 37868
rect 29920 37816 29972 37868
rect 30288 37816 30340 37868
rect 29092 37748 29144 37800
rect 29460 37748 29512 37800
rect 1860 37723 1912 37732
rect 1860 37689 1869 37723
rect 1869 37689 1903 37723
rect 1903 37689 1912 37723
rect 1860 37680 1912 37689
rect 22008 37723 22060 37732
rect 22008 37689 22017 37723
rect 22017 37689 22051 37723
rect 22051 37689 22060 37723
rect 22008 37680 22060 37689
rect 22284 37680 22336 37732
rect 22560 37612 22612 37664
rect 22836 37612 22888 37664
rect 23388 37680 23440 37732
rect 24860 37680 24912 37732
rect 26424 37723 26476 37732
rect 26424 37689 26433 37723
rect 26433 37689 26467 37723
rect 26467 37689 26476 37723
rect 26424 37680 26476 37689
rect 24216 37655 24268 37664
rect 24216 37621 24225 37655
rect 24225 37621 24259 37655
rect 24259 37621 24268 37655
rect 24216 37612 24268 37621
rect 24676 37612 24728 37664
rect 30288 37680 30340 37732
rect 28448 37612 28500 37664
rect 28908 37612 28960 37664
rect 30380 37612 30432 37664
rect 30840 37952 30892 38004
rect 36912 37952 36964 38004
rect 30656 37680 30708 37732
rect 35716 37884 35768 37936
rect 31484 37816 31536 37868
rect 36176 37791 36228 37800
rect 36176 37757 36185 37791
rect 36185 37757 36219 37791
rect 36219 37757 36228 37791
rect 36176 37748 36228 37757
rect 37096 37723 37148 37732
rect 37096 37689 37105 37723
rect 37105 37689 37139 37723
rect 37139 37689 37148 37723
rect 37096 37680 37148 37689
rect 38476 37816 38528 37868
rect 37740 37791 37792 37800
rect 37740 37757 37749 37791
rect 37749 37757 37783 37791
rect 37783 37757 37792 37791
rect 37740 37748 37792 37757
rect 38292 37748 38344 37800
rect 35164 37612 35216 37664
rect 35348 37612 35400 37664
rect 35532 37612 35584 37664
rect 35992 37612 36044 37664
rect 36176 37612 36228 37664
rect 37372 37612 37424 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 17868 37272 17920 37324
rect 24676 37408 24728 37460
rect 21548 37340 21600 37392
rect 22836 37272 22888 37324
rect 23388 37272 23440 37324
rect 21732 37204 21784 37256
rect 23572 37247 23624 37256
rect 20352 37136 20404 37188
rect 22560 37136 22612 37188
rect 23204 37136 23256 37188
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 24032 37340 24084 37392
rect 24308 37383 24360 37392
rect 24308 37349 24338 37383
rect 24338 37349 24360 37383
rect 24308 37340 24360 37349
rect 26424 37383 26476 37392
rect 26424 37349 26433 37383
rect 26433 37349 26467 37383
rect 26467 37349 26476 37383
rect 26424 37340 26476 37349
rect 28080 37408 28132 37460
rect 29460 37408 29512 37460
rect 30380 37408 30432 37460
rect 32312 37408 32364 37460
rect 35164 37408 35216 37460
rect 36360 37408 36412 37460
rect 23572 37068 23624 37120
rect 26608 37315 26660 37324
rect 26608 37281 26622 37315
rect 26622 37281 26656 37315
rect 26656 37281 26660 37315
rect 26608 37272 26660 37281
rect 26516 37204 26568 37256
rect 26884 37272 26936 37324
rect 28908 37272 28960 37324
rect 29092 37272 29144 37324
rect 29460 37272 29512 37324
rect 29828 37315 29880 37324
rect 29828 37281 29837 37315
rect 29837 37281 29871 37315
rect 29871 37281 29880 37315
rect 29828 37272 29880 37281
rect 30012 37272 30064 37324
rect 29736 37247 29788 37256
rect 29736 37213 29745 37247
rect 29745 37213 29779 37247
rect 29779 37213 29788 37247
rect 29736 37204 29788 37213
rect 30288 37340 30340 37392
rect 35532 37315 35584 37324
rect 35532 37281 35541 37315
rect 35541 37281 35575 37315
rect 35575 37281 35584 37315
rect 35532 37272 35584 37281
rect 36360 37315 36412 37324
rect 36360 37281 36369 37315
rect 36369 37281 36403 37315
rect 36403 37281 36412 37315
rect 36360 37272 36412 37281
rect 37372 37340 37424 37392
rect 26884 37136 26936 37188
rect 27712 37136 27764 37188
rect 31852 37204 31904 37256
rect 35624 37204 35676 37256
rect 38476 37272 38528 37324
rect 37740 37204 37792 37256
rect 35992 37136 36044 37188
rect 38752 37136 38804 37188
rect 27344 37068 27396 37120
rect 28264 37068 28316 37120
rect 29736 37068 29788 37120
rect 36912 37068 36964 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 1584 36907 1636 36916
rect 1584 36873 1593 36907
rect 1593 36873 1627 36907
rect 1627 36873 1636 36907
rect 1584 36864 1636 36873
rect 23480 36907 23532 36916
rect 23480 36873 23489 36907
rect 23489 36873 23523 36907
rect 23523 36873 23532 36907
rect 23480 36864 23532 36873
rect 23572 36864 23624 36916
rect 25228 36864 25280 36916
rect 26332 36864 26384 36916
rect 26608 36864 26660 36916
rect 26700 36864 26752 36916
rect 29460 36864 29512 36916
rect 31392 36864 31444 36916
rect 35900 36864 35952 36916
rect 36176 36864 36228 36916
rect 22560 36796 22612 36848
rect 7104 36728 7156 36780
rect 15936 36728 15988 36780
rect 21732 36728 21784 36780
rect 23480 36728 23532 36780
rect 1400 36703 1452 36712
rect 1400 36669 1409 36703
rect 1409 36669 1443 36703
rect 1443 36669 1452 36703
rect 1400 36660 1452 36669
rect 22468 36660 22520 36712
rect 23572 36660 23624 36712
rect 24400 36728 24452 36780
rect 8760 36524 8812 36576
rect 20168 36592 20220 36644
rect 23204 36592 23256 36644
rect 26240 36703 26292 36712
rect 26240 36669 26249 36703
rect 26249 36669 26283 36703
rect 26283 36669 26292 36703
rect 26240 36660 26292 36669
rect 26516 36703 26568 36712
rect 26516 36669 26525 36703
rect 26525 36669 26559 36703
rect 26559 36669 26568 36703
rect 26516 36660 26568 36669
rect 26608 36703 26660 36712
rect 26608 36669 26622 36703
rect 26622 36669 26656 36703
rect 26656 36669 26660 36703
rect 27988 36728 28040 36780
rect 29920 36728 29972 36780
rect 26608 36660 26660 36669
rect 26424 36635 26476 36644
rect 22284 36524 22336 36576
rect 23296 36524 23348 36576
rect 26424 36601 26433 36635
rect 26433 36601 26467 36635
rect 26467 36601 26476 36635
rect 26424 36592 26476 36601
rect 27988 36592 28040 36644
rect 29092 36660 29144 36712
rect 30012 36660 30064 36712
rect 36084 36660 36136 36712
rect 36360 36660 36412 36712
rect 36452 36660 36504 36712
rect 37004 36660 37056 36712
rect 37924 36703 37976 36712
rect 37924 36669 37933 36703
rect 37933 36669 37967 36703
rect 37967 36669 37976 36703
rect 37924 36660 37976 36669
rect 35624 36592 35676 36644
rect 37372 36592 37424 36644
rect 37740 36635 37792 36644
rect 26332 36524 26384 36576
rect 26700 36524 26752 36576
rect 27712 36524 27764 36576
rect 35992 36567 36044 36576
rect 35992 36533 36001 36567
rect 36001 36533 36035 36567
rect 36035 36533 36044 36567
rect 35992 36524 36044 36533
rect 36084 36524 36136 36576
rect 37740 36601 37749 36635
rect 37749 36601 37783 36635
rect 37783 36601 37792 36635
rect 37740 36592 37792 36601
rect 37832 36635 37884 36644
rect 37832 36601 37841 36635
rect 37841 36601 37875 36635
rect 37875 36601 37884 36635
rect 37832 36592 37884 36601
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 1676 36320 1728 36372
rect 1768 36320 1820 36372
rect 26608 36320 26660 36372
rect 27160 36320 27212 36372
rect 33048 36320 33100 36372
rect 34796 36363 34848 36372
rect 34796 36329 34805 36363
rect 34805 36329 34839 36363
rect 34839 36329 34848 36363
rect 34796 36320 34848 36329
rect 35900 36320 35952 36372
rect 2044 36252 2096 36304
rect 1400 36227 1452 36236
rect 1400 36193 1409 36227
rect 1409 36193 1443 36227
rect 1443 36193 1452 36227
rect 1400 36184 1452 36193
rect 21456 36227 21508 36236
rect 21456 36193 21465 36227
rect 21465 36193 21499 36227
rect 21499 36193 21508 36227
rect 21456 36184 21508 36193
rect 22836 36184 22888 36236
rect 24216 36184 24268 36236
rect 22284 36116 22336 36168
rect 22468 36116 22520 36168
rect 26332 36184 26384 36236
rect 26516 36227 26568 36236
rect 26516 36193 26525 36227
rect 26525 36193 26559 36227
rect 26559 36193 26568 36227
rect 26516 36184 26568 36193
rect 27344 36252 27396 36304
rect 31852 36252 31904 36304
rect 26976 36184 27028 36236
rect 34796 36184 34848 36236
rect 35440 36227 35492 36236
rect 35440 36193 35449 36227
rect 35449 36193 35483 36227
rect 35483 36193 35492 36227
rect 35440 36184 35492 36193
rect 35900 36227 35952 36236
rect 35900 36193 35909 36227
rect 35909 36193 35943 36227
rect 35943 36193 35952 36227
rect 35900 36184 35952 36193
rect 36820 36320 36872 36372
rect 38936 36320 38988 36372
rect 37464 36252 37516 36304
rect 27344 36116 27396 36168
rect 35808 36116 35860 36168
rect 36360 36227 36412 36236
rect 36360 36193 36374 36227
rect 36374 36193 36408 36227
rect 36408 36193 36412 36227
rect 36360 36184 36412 36193
rect 24676 36048 24728 36100
rect 23388 35980 23440 36032
rect 24400 35980 24452 36032
rect 27528 35980 27580 36032
rect 27804 35980 27856 36032
rect 30288 35980 30340 36032
rect 34520 35980 34572 36032
rect 34612 35980 34664 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 23204 35776 23256 35828
rect 26332 35776 26384 35828
rect 27160 35776 27212 35828
rect 27804 35776 27856 35828
rect 28724 35776 28776 35828
rect 33324 35776 33376 35828
rect 33968 35776 34020 35828
rect 35256 35776 35308 35828
rect 35900 35776 35952 35828
rect 37556 35776 37608 35828
rect 7840 35708 7892 35760
rect 14832 35708 14884 35760
rect 20536 35708 20588 35760
rect 22836 35640 22888 35692
rect 26792 35640 26844 35692
rect 31944 35640 31996 35692
rect 8392 35504 8444 35556
rect 15752 35504 15804 35556
rect 23572 35572 23624 35624
rect 26240 35572 26292 35624
rect 33232 35572 33284 35624
rect 34796 35615 34848 35624
rect 34796 35581 34805 35615
rect 34805 35581 34839 35615
rect 34839 35581 34848 35615
rect 34796 35572 34848 35581
rect 35532 35572 35584 35624
rect 35900 35615 35952 35624
rect 35900 35581 35909 35615
rect 35909 35581 35943 35615
rect 35943 35581 35952 35615
rect 35900 35572 35952 35581
rect 36452 35640 36504 35692
rect 36820 35640 36872 35692
rect 24308 35504 24360 35556
rect 26976 35504 27028 35556
rect 33324 35504 33376 35556
rect 35348 35504 35400 35556
rect 36360 35615 36412 35624
rect 36360 35581 36374 35615
rect 36374 35581 36408 35615
rect 36408 35581 36412 35615
rect 37280 35640 37332 35692
rect 36360 35572 36412 35581
rect 23480 35436 23532 35488
rect 26608 35436 26660 35488
rect 31576 35436 31628 35488
rect 33048 35436 33100 35488
rect 36820 35504 36872 35556
rect 37464 35547 37516 35556
rect 37464 35513 37473 35547
rect 37473 35513 37507 35547
rect 37507 35513 37516 35547
rect 37464 35504 37516 35513
rect 38752 35436 38804 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 2504 35232 2556 35284
rect 2412 35164 2464 35216
rect 4804 35164 4856 35216
rect 23204 35232 23256 35284
rect 26240 35232 26292 35284
rect 28632 35232 28684 35284
rect 31392 35232 31444 35284
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 23112 35164 23164 35216
rect 18604 35096 18656 35148
rect 22468 35096 22520 35148
rect 23388 35139 23440 35148
rect 23388 35105 23397 35139
rect 23397 35105 23431 35139
rect 23431 35105 23440 35139
rect 23388 35096 23440 35105
rect 20904 35028 20956 35080
rect 27528 35096 27580 35148
rect 28448 35096 28500 35148
rect 34612 35164 34664 35216
rect 35900 35164 35952 35216
rect 36365 35207 36417 35216
rect 36365 35173 36369 35207
rect 36369 35173 36403 35207
rect 36403 35173 36417 35207
rect 36365 35164 36417 35173
rect 34520 35096 34572 35148
rect 35624 35096 35676 35148
rect 36268 35139 36320 35148
rect 36268 35105 36275 35139
rect 36275 35105 36320 35139
rect 36268 35096 36320 35105
rect 36452 35139 36504 35148
rect 36452 35105 36461 35139
rect 36461 35105 36495 35139
rect 36495 35105 36504 35139
rect 36452 35096 36504 35105
rect 18512 34892 18564 34944
rect 25872 34960 25924 35012
rect 29920 35028 29972 35080
rect 30656 35028 30708 35080
rect 37280 35096 37332 35148
rect 29276 34892 29328 34944
rect 35532 34935 35584 34944
rect 35532 34901 35541 34935
rect 35541 34901 35575 34935
rect 35575 34901 35584 34935
rect 35532 34892 35584 34901
rect 35624 34892 35676 34944
rect 36636 34892 36688 34944
rect 37832 34892 37884 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 1768 34688 1820 34740
rect 20628 34552 20680 34604
rect 22560 34620 22612 34672
rect 24216 34620 24268 34672
rect 27988 34620 28040 34672
rect 29000 34620 29052 34672
rect 29828 34620 29880 34672
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 10692 34484 10744 34536
rect 11796 34484 11848 34536
rect 11888 34484 11940 34536
rect 17776 34484 17828 34536
rect 22284 34484 22336 34536
rect 22560 34484 22612 34536
rect 26516 34484 26568 34536
rect 25872 34348 25924 34400
rect 28724 34552 28776 34604
rect 27712 34484 27764 34536
rect 29460 34552 29512 34604
rect 36636 34620 36688 34672
rect 37556 34620 37608 34672
rect 34612 34527 34664 34536
rect 29092 34416 29144 34468
rect 34612 34493 34621 34527
rect 34621 34493 34655 34527
rect 34655 34493 34664 34527
rect 34612 34484 34664 34493
rect 35532 34484 35584 34536
rect 35624 34416 35676 34468
rect 36360 34527 36412 34536
rect 36360 34493 36369 34527
rect 36369 34493 36403 34527
rect 36403 34493 36412 34527
rect 36360 34484 36412 34493
rect 37648 34484 37700 34536
rect 37832 34527 37884 34536
rect 37832 34493 37841 34527
rect 37841 34493 37875 34527
rect 37875 34493 37884 34527
rect 37832 34484 37884 34493
rect 38568 34484 38620 34536
rect 36453 34459 36505 34468
rect 36453 34425 36461 34459
rect 36461 34425 36495 34459
rect 36495 34425 36505 34459
rect 37740 34459 37792 34468
rect 36453 34416 36505 34425
rect 37740 34425 37749 34459
rect 37749 34425 37783 34459
rect 37783 34425 37792 34459
rect 37740 34416 37792 34425
rect 27712 34348 27764 34400
rect 28632 34391 28684 34400
rect 28632 34357 28641 34391
rect 28641 34357 28675 34391
rect 28675 34357 28684 34391
rect 28632 34348 28684 34357
rect 28816 34348 28868 34400
rect 36728 34391 36780 34400
rect 36728 34357 36737 34391
rect 36737 34357 36771 34391
rect 36771 34357 36780 34391
rect 36728 34348 36780 34357
rect 38108 34391 38160 34400
rect 38108 34357 38117 34391
rect 38117 34357 38151 34391
rect 38151 34357 38160 34391
rect 38108 34348 38160 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 28448 34144 28500 34196
rect 28908 34144 28960 34196
rect 30012 34144 30064 34196
rect 30748 34144 30800 34196
rect 36728 34144 36780 34196
rect 37188 34187 37240 34196
rect 37188 34153 37197 34187
rect 37197 34153 37231 34187
rect 37231 34153 37240 34187
rect 37188 34144 37240 34153
rect 18328 34076 18380 34128
rect 35532 34076 35584 34128
rect 35900 34076 35952 34128
rect 36360 34119 36412 34128
rect 25412 34051 25464 34060
rect 25412 34017 25421 34051
rect 25421 34017 25455 34051
rect 25455 34017 25464 34051
rect 25412 34008 25464 34017
rect 26792 34008 26844 34060
rect 23112 33940 23164 33992
rect 24676 33940 24728 33992
rect 26608 33983 26660 33992
rect 26608 33949 26617 33983
rect 26617 33949 26651 33983
rect 26651 33949 26660 33983
rect 26608 33940 26660 33949
rect 26700 33983 26752 33992
rect 26700 33949 26709 33983
rect 26709 33949 26743 33983
rect 26743 33949 26752 33983
rect 26700 33940 26752 33949
rect 7840 33872 7892 33924
rect 18420 33872 18472 33924
rect 27068 33872 27120 33924
rect 2136 33804 2188 33856
rect 18052 33804 18104 33856
rect 24952 33804 25004 33856
rect 26608 33804 26660 33856
rect 27712 34008 27764 34060
rect 28080 34051 28132 34060
rect 28080 34017 28114 34051
rect 28114 34017 28132 34051
rect 28080 34008 28132 34017
rect 28448 34008 28500 34060
rect 29828 34051 29880 34060
rect 29828 34017 29837 34051
rect 29837 34017 29871 34051
rect 29871 34017 29880 34051
rect 29828 34008 29880 34017
rect 35624 34051 35676 34060
rect 35624 34017 35633 34051
rect 35633 34017 35667 34051
rect 35667 34017 35676 34051
rect 35624 34008 35676 34017
rect 36360 34085 36369 34119
rect 36369 34085 36403 34119
rect 36403 34085 36412 34119
rect 36360 34076 36412 34085
rect 36452 34051 36504 34060
rect 30196 33940 30248 33992
rect 30012 33872 30064 33924
rect 36452 34017 36461 34051
rect 36461 34017 36495 34051
rect 36495 34017 36504 34051
rect 36452 34008 36504 34017
rect 36728 34008 36780 34060
rect 37372 34051 37424 34060
rect 37372 34017 37381 34051
rect 37381 34017 37415 34051
rect 37415 34017 37424 34051
rect 37372 34008 37424 34017
rect 27712 33804 27764 33856
rect 29092 33804 29144 33856
rect 35716 33804 35768 33856
rect 36912 33872 36964 33924
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 25780 33643 25832 33652
rect 25780 33609 25789 33643
rect 25789 33609 25823 33643
rect 25823 33609 25832 33643
rect 25780 33600 25832 33609
rect 2044 33575 2096 33584
rect 2044 33541 2053 33575
rect 2053 33541 2087 33575
rect 2087 33541 2096 33575
rect 2044 33532 2096 33541
rect 18788 33532 18840 33584
rect 1860 33439 1912 33448
rect 1860 33405 1869 33439
rect 1869 33405 1903 33439
rect 1903 33405 1912 33439
rect 1860 33396 1912 33405
rect 1952 33396 2004 33448
rect 25780 33464 25832 33516
rect 27988 33532 28040 33584
rect 28448 33532 28500 33584
rect 29000 33464 29052 33516
rect 38200 33600 38252 33652
rect 35900 33532 35952 33584
rect 36176 33532 36228 33584
rect 39028 33532 39080 33584
rect 25872 33396 25924 33448
rect 10140 33260 10192 33312
rect 14464 33260 14516 33312
rect 25320 33260 25372 33312
rect 25504 33371 25556 33380
rect 25504 33337 25513 33371
rect 25513 33337 25547 33371
rect 25547 33337 25556 33371
rect 25504 33328 25556 33337
rect 26884 33396 26936 33448
rect 28356 33396 28408 33448
rect 26516 33328 26568 33380
rect 27068 33328 27120 33380
rect 28540 33328 28592 33380
rect 36084 33439 36136 33448
rect 36084 33405 36093 33439
rect 36093 33405 36127 33439
rect 36127 33405 36136 33439
rect 36084 33396 36136 33405
rect 36176 33439 36228 33448
rect 36176 33405 36186 33439
rect 36186 33405 36220 33439
rect 36220 33405 36228 33439
rect 36176 33396 36228 33405
rect 37464 33439 37516 33448
rect 37464 33405 37473 33439
rect 37473 33405 37507 33439
rect 37507 33405 37516 33439
rect 37464 33396 37516 33405
rect 38016 33396 38068 33448
rect 29092 33328 29144 33380
rect 36360 33371 36412 33380
rect 36360 33337 36369 33371
rect 36369 33337 36403 33371
rect 36403 33337 36412 33371
rect 36360 33328 36412 33337
rect 36452 33371 36504 33380
rect 36452 33337 36461 33371
rect 36461 33337 36495 33371
rect 36495 33337 36504 33371
rect 36452 33328 36504 33337
rect 26884 33260 26936 33312
rect 27620 33260 27672 33312
rect 29736 33260 29788 33312
rect 35624 33260 35676 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 1952 33056 2004 33108
rect 24676 33056 24728 33108
rect 1860 32988 1912 33040
rect 22836 32988 22888 33040
rect 26884 33056 26936 33108
rect 29184 33099 29236 33108
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 1584 32852 1636 32904
rect 24860 32920 24912 32972
rect 25320 32963 25372 32972
rect 25320 32929 25329 32963
rect 25329 32929 25363 32963
rect 25363 32929 25372 32963
rect 25320 32920 25372 32929
rect 26424 32963 26476 32972
rect 26424 32929 26433 32963
rect 26433 32929 26467 32963
rect 26467 32929 26476 32963
rect 26424 32920 26476 32929
rect 26516 32920 26568 32972
rect 26332 32852 26384 32904
rect 25504 32784 25556 32836
rect 25688 32827 25740 32836
rect 25688 32793 25697 32827
rect 25697 32793 25731 32827
rect 25731 32793 25740 32827
rect 25688 32784 25740 32793
rect 26332 32716 26384 32768
rect 29184 33065 29193 33099
rect 29193 33065 29227 33099
rect 29227 33065 29236 33099
rect 29184 33056 29236 33065
rect 27896 32988 27948 33040
rect 32864 33056 32916 33108
rect 33968 33056 34020 33108
rect 36544 33056 36596 33108
rect 36360 33031 36412 33040
rect 36360 32997 36369 33031
rect 36369 32997 36403 33031
rect 36403 32997 36412 33031
rect 36360 32988 36412 32997
rect 33968 32920 34020 32972
rect 34152 32920 34204 32972
rect 35440 32963 35492 32972
rect 35440 32929 35449 32963
rect 35449 32929 35483 32963
rect 35483 32929 35492 32963
rect 35440 32920 35492 32929
rect 36084 32963 36136 32972
rect 36084 32929 36093 32963
rect 36093 32929 36127 32963
rect 36127 32929 36136 32963
rect 36084 32920 36136 32929
rect 36452 32963 36504 32972
rect 36452 32929 36461 32963
rect 36461 32929 36495 32963
rect 36495 32929 36504 32963
rect 36452 32920 36504 32929
rect 36544 32963 36596 32972
rect 36544 32929 36558 32963
rect 36558 32929 36592 32963
rect 36592 32929 36596 32963
rect 37372 32963 37424 32972
rect 36544 32920 36596 32929
rect 37372 32929 37381 32963
rect 37381 32929 37415 32963
rect 37415 32929 37424 32963
rect 37372 32920 37424 32929
rect 37648 32852 37700 32904
rect 27712 32784 27764 32836
rect 26976 32716 27028 32768
rect 27988 32716 28040 32768
rect 29920 32784 29972 32836
rect 35256 32784 35308 32836
rect 29276 32716 29328 32768
rect 30656 32716 30708 32768
rect 36360 32716 36412 32768
rect 37188 32716 37240 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 24032 32444 24084 32496
rect 25228 32444 25280 32496
rect 25504 32444 25556 32496
rect 25688 32444 25740 32496
rect 4712 32308 4764 32360
rect 25320 32308 25372 32360
rect 26056 32512 26108 32564
rect 26976 32512 27028 32564
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 27712 32512 27764 32564
rect 28172 32555 28224 32564
rect 28172 32521 28181 32555
rect 28181 32521 28215 32555
rect 28215 32521 28224 32555
rect 28172 32512 28224 32521
rect 36452 32512 36504 32564
rect 36544 32512 36596 32564
rect 36728 32512 36780 32564
rect 22836 32240 22888 32292
rect 24308 32240 24360 32292
rect 25688 32283 25740 32292
rect 25688 32249 25697 32283
rect 25697 32249 25731 32283
rect 25731 32249 25740 32283
rect 25688 32240 25740 32249
rect 25320 32172 25372 32224
rect 27436 32376 27488 32428
rect 27896 32444 27948 32496
rect 31760 32376 31812 32428
rect 36544 32376 36596 32428
rect 39488 32444 39540 32496
rect 27988 32351 28040 32360
rect 27344 32172 27396 32224
rect 27988 32317 28002 32351
rect 28002 32317 28036 32351
rect 28036 32317 28040 32351
rect 27988 32308 28040 32317
rect 28264 32308 28316 32360
rect 28632 32308 28684 32360
rect 35900 32308 35952 32360
rect 36728 32308 36780 32360
rect 36912 32351 36964 32360
rect 36912 32317 36921 32351
rect 36921 32317 36955 32351
rect 36955 32317 36964 32351
rect 36912 32308 36964 32317
rect 38384 32376 38436 32428
rect 38936 32308 38988 32360
rect 27896 32283 27948 32292
rect 27896 32249 27905 32283
rect 27905 32249 27939 32283
rect 27939 32249 27948 32283
rect 27896 32240 27948 32249
rect 27988 32172 28040 32224
rect 28632 32172 28684 32224
rect 31576 32240 31628 32292
rect 37740 32283 37792 32292
rect 37740 32249 37749 32283
rect 37749 32249 37783 32283
rect 37783 32249 37792 32283
rect 37740 32240 37792 32249
rect 37832 32283 37884 32292
rect 37832 32249 37841 32283
rect 37841 32249 37875 32283
rect 37875 32249 37884 32283
rect 37832 32240 37884 32249
rect 37464 32172 37516 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 1584 32011 1636 32020
rect 1584 31977 1593 32011
rect 1593 31977 1627 32011
rect 1627 31977 1636 32011
rect 1584 31968 1636 31977
rect 2780 31900 2832 31952
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 15292 31900 15344 31952
rect 23388 31900 23440 31952
rect 24952 31900 25004 31952
rect 22100 31832 22152 31884
rect 22836 31832 22888 31884
rect 24676 31832 24728 31884
rect 24860 31628 24912 31680
rect 25688 31968 25740 32020
rect 26056 31968 26108 32020
rect 27528 31968 27580 32020
rect 27896 31968 27948 32020
rect 28356 32011 28408 32020
rect 25504 31900 25556 31952
rect 27436 31900 27488 31952
rect 28356 31977 28373 32011
rect 28373 31977 28407 32011
rect 28407 31977 28408 32011
rect 28356 31968 28408 31977
rect 30932 31968 30984 32020
rect 26056 31832 26108 31884
rect 25504 31764 25556 31816
rect 25044 31696 25096 31748
rect 26884 31832 26936 31884
rect 27804 31875 27856 31884
rect 27804 31841 27813 31875
rect 27813 31841 27847 31875
rect 27847 31841 27856 31875
rect 27804 31832 27856 31841
rect 27896 31832 27948 31884
rect 34152 31832 34204 31884
rect 34520 31832 34572 31884
rect 35532 31875 35584 31884
rect 35532 31841 35541 31875
rect 35541 31841 35575 31875
rect 35575 31841 35584 31875
rect 35532 31832 35584 31841
rect 36176 31875 36228 31884
rect 36176 31841 36185 31875
rect 36185 31841 36219 31875
rect 36219 31841 36228 31875
rect 36176 31832 36228 31841
rect 36452 31900 36504 31952
rect 37188 31968 37240 32020
rect 37832 31900 37884 31952
rect 33324 31764 33376 31816
rect 34336 31764 34388 31816
rect 36544 31832 36596 31884
rect 37188 31875 37240 31884
rect 37188 31841 37197 31875
rect 37197 31841 37231 31875
rect 37231 31841 37240 31875
rect 37188 31832 37240 31841
rect 38844 31764 38896 31816
rect 25228 31628 25280 31680
rect 26240 31696 26292 31748
rect 26976 31696 27028 31748
rect 27344 31696 27396 31748
rect 34152 31696 34204 31748
rect 34796 31696 34848 31748
rect 35900 31696 35952 31748
rect 36728 31696 36780 31748
rect 36544 31628 36596 31680
rect 37004 31628 37056 31680
rect 37372 31671 37424 31680
rect 37372 31637 37381 31671
rect 37381 31637 37415 31671
rect 37415 31637 37424 31671
rect 37372 31628 37424 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 1860 31424 1912 31476
rect 2044 31288 2096 31340
rect 23572 31288 23624 31340
rect 26884 31356 26936 31408
rect 26792 31288 26844 31340
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 21732 31152 21784 31204
rect 26884 31220 26936 31272
rect 27344 31288 27396 31340
rect 27712 31424 27764 31476
rect 28540 31424 28592 31476
rect 36452 31424 36504 31476
rect 37740 31424 37792 31476
rect 27896 31356 27948 31408
rect 31024 31356 31076 31408
rect 31116 31288 31168 31340
rect 27528 31263 27580 31272
rect 27528 31229 27531 31263
rect 27531 31229 27580 31263
rect 27528 31220 27580 31229
rect 27896 31220 27948 31272
rect 29828 31220 29880 31272
rect 25320 31195 25372 31204
rect 25320 31161 25329 31195
rect 25329 31161 25363 31195
rect 25363 31161 25372 31195
rect 25320 31152 25372 31161
rect 9312 31084 9364 31136
rect 20076 31084 20128 31136
rect 24952 31084 25004 31136
rect 25504 31084 25556 31136
rect 27344 31195 27396 31204
rect 27344 31161 27353 31195
rect 27353 31161 27387 31195
rect 27387 31161 27396 31195
rect 38660 31356 38712 31408
rect 36912 31263 36964 31272
rect 36912 31229 36921 31263
rect 36921 31229 36955 31263
rect 36955 31229 36964 31263
rect 36912 31220 36964 31229
rect 39120 31288 39172 31340
rect 37832 31263 37884 31272
rect 27344 31152 27396 31161
rect 37280 31152 37332 31204
rect 37832 31229 37841 31263
rect 37841 31229 37875 31263
rect 37875 31229 37884 31263
rect 37832 31220 37884 31229
rect 38016 31220 38068 31272
rect 37740 31195 37792 31204
rect 37740 31161 37749 31195
rect 37749 31161 37783 31195
rect 37783 31161 37792 31195
rect 37740 31152 37792 31161
rect 32496 31084 32548 31136
rect 37004 31084 37056 31136
rect 37188 31084 37240 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 24952 30880 25004 30932
rect 25044 30812 25096 30864
rect 25412 30812 25464 30864
rect 26608 30812 26660 30864
rect 25044 30676 25096 30728
rect 25872 30744 25924 30796
rect 27896 30880 27948 30932
rect 34060 30880 34112 30932
rect 36268 30880 36320 30932
rect 37280 30880 37332 30932
rect 34520 30812 34572 30864
rect 35256 30812 35308 30864
rect 35808 30744 35860 30796
rect 36728 30787 36780 30796
rect 36728 30753 36737 30787
rect 36737 30753 36771 30787
rect 36771 30753 36780 30787
rect 36728 30744 36780 30753
rect 23940 30608 23992 30660
rect 24676 30608 24728 30660
rect 26424 30608 26476 30660
rect 26608 30608 26660 30660
rect 26976 30608 27028 30660
rect 27896 30608 27948 30660
rect 34060 30608 34112 30660
rect 36360 30608 36412 30660
rect 26240 30540 26292 30592
rect 26700 30583 26752 30592
rect 26700 30549 26709 30583
rect 26709 30549 26743 30583
rect 26743 30549 26752 30583
rect 26700 30540 26752 30549
rect 26884 30540 26936 30592
rect 28632 30540 28684 30592
rect 35440 30540 35492 30592
rect 35716 30540 35768 30592
rect 35992 30540 36044 30592
rect 36176 30540 36228 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 2780 30336 2832 30388
rect 27344 30336 27396 30388
rect 33600 30336 33652 30388
rect 34612 30336 34664 30388
rect 4712 30268 4764 30320
rect 26424 30268 26476 30320
rect 1216 30200 1268 30252
rect 23388 30200 23440 30252
rect 23940 30200 23992 30252
rect 24400 30200 24452 30252
rect 26240 30200 26292 30252
rect 1400 30175 1452 30184
rect 1400 30141 1409 30175
rect 1409 30141 1443 30175
rect 1443 30141 1452 30175
rect 1400 30132 1452 30141
rect 25044 30132 25096 30184
rect 22376 30064 22428 30116
rect 23296 30064 23348 30116
rect 23388 30064 23440 30116
rect 25320 30064 25372 30116
rect 26332 30132 26384 30184
rect 28264 30132 28316 30184
rect 28356 30132 28408 30184
rect 34704 30200 34756 30252
rect 35992 30175 36044 30184
rect 35992 30141 36001 30175
rect 36001 30141 36035 30175
rect 36035 30141 36044 30175
rect 35992 30132 36044 30141
rect 19984 29996 20036 30048
rect 28448 29996 28500 30048
rect 28724 29996 28776 30048
rect 34980 30064 35032 30116
rect 36176 30132 36228 30184
rect 36360 30175 36412 30184
rect 36360 30141 36369 30175
rect 36369 30141 36403 30175
rect 36403 30141 36412 30175
rect 36360 30132 36412 30141
rect 37832 30175 37884 30184
rect 37832 30141 37841 30175
rect 37841 30141 37875 30175
rect 37875 30141 37884 30175
rect 37832 30132 37884 30141
rect 38200 30132 38252 30184
rect 37280 30064 37332 30116
rect 37740 30107 37792 30116
rect 37740 30073 37749 30107
rect 37749 30073 37783 30107
rect 37783 30073 37792 30107
rect 37740 30064 37792 30073
rect 36452 29996 36504 30048
rect 36728 29996 36780 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 19248 29792 19300 29844
rect 23940 29792 23992 29844
rect 36176 29792 36228 29844
rect 17592 29656 17644 29708
rect 18972 29699 19024 29708
rect 18972 29665 18979 29699
rect 18979 29665 19024 29699
rect 18972 29656 19024 29665
rect 1676 29588 1728 29640
rect 15292 29588 15344 29640
rect 18328 29588 18380 29640
rect 4896 29520 4948 29572
rect 18880 29452 18932 29504
rect 25228 29724 25280 29776
rect 26516 29724 26568 29776
rect 32956 29724 33008 29776
rect 20352 29656 20404 29708
rect 22928 29699 22980 29708
rect 22928 29665 22937 29699
rect 22937 29665 22971 29699
rect 22971 29665 22980 29699
rect 22928 29656 22980 29665
rect 24032 29656 24084 29708
rect 24216 29656 24268 29708
rect 26332 29656 26384 29708
rect 26884 29699 26936 29708
rect 21456 29588 21508 29640
rect 23572 29588 23624 29640
rect 26516 29631 26568 29640
rect 26516 29597 26525 29631
rect 26525 29597 26559 29631
rect 26559 29597 26568 29631
rect 26516 29588 26568 29597
rect 26884 29665 26893 29699
rect 26893 29665 26927 29699
rect 26927 29665 26936 29699
rect 26884 29656 26936 29665
rect 27528 29656 27580 29708
rect 30288 29656 30340 29708
rect 35808 29656 35860 29708
rect 36360 29767 36412 29776
rect 36360 29733 36369 29767
rect 36369 29733 36403 29767
rect 36403 29733 36412 29767
rect 38292 29792 38344 29844
rect 36360 29724 36412 29733
rect 37740 29724 37792 29776
rect 23112 29520 23164 29572
rect 25688 29563 25740 29572
rect 25688 29529 25697 29563
rect 25697 29529 25731 29563
rect 25731 29529 25740 29563
rect 25688 29520 25740 29529
rect 26976 29588 27028 29640
rect 29276 29588 29328 29640
rect 36268 29699 36320 29708
rect 36268 29665 36277 29699
rect 36277 29665 36311 29699
rect 36311 29665 36320 29699
rect 36268 29656 36320 29665
rect 36452 29699 36504 29708
rect 36452 29665 36466 29699
rect 36466 29665 36500 29699
rect 36500 29665 36504 29699
rect 37372 29699 37424 29708
rect 36452 29656 36504 29665
rect 37372 29665 37381 29699
rect 37381 29665 37415 29699
rect 37415 29665 37424 29699
rect 37372 29656 37424 29665
rect 37188 29588 37240 29640
rect 22928 29452 22980 29504
rect 23940 29452 23992 29504
rect 26240 29495 26292 29504
rect 26240 29461 26249 29495
rect 26249 29461 26283 29495
rect 26283 29461 26292 29495
rect 26240 29452 26292 29461
rect 31116 29520 31168 29572
rect 34612 29520 34664 29572
rect 34980 29520 35032 29572
rect 35440 29520 35492 29572
rect 32312 29452 32364 29504
rect 35992 29452 36044 29504
rect 38752 29452 38804 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 2688 29248 2740 29300
rect 18880 29248 18932 29300
rect 20260 29248 20312 29300
rect 1400 29087 1452 29096
rect 1400 29053 1409 29087
rect 1409 29053 1443 29087
rect 1443 29053 1452 29087
rect 1400 29044 1452 29053
rect 6552 28976 6604 29028
rect 17408 29044 17460 29096
rect 23940 29180 23992 29232
rect 18880 29087 18932 29096
rect 22560 29112 22612 29164
rect 23296 29112 23348 29164
rect 26516 29248 26568 29300
rect 26976 29248 27028 29300
rect 24308 29180 24360 29232
rect 27528 29180 27580 29232
rect 18880 29053 18894 29087
rect 18894 29053 18928 29087
rect 18928 29053 18932 29087
rect 18880 29044 18932 29053
rect 22468 29087 22520 29096
rect 22468 29053 22477 29087
rect 22477 29053 22511 29087
rect 22511 29053 22520 29087
rect 22468 29044 22520 29053
rect 23480 29044 23532 29096
rect 24584 29112 24636 29164
rect 26976 29112 27028 29164
rect 31852 29180 31904 29232
rect 35072 29180 35124 29232
rect 18328 28976 18380 29028
rect 19156 28976 19208 29028
rect 20720 28976 20772 29028
rect 24216 29087 24268 29096
rect 24216 29053 24225 29087
rect 24225 29053 24259 29087
rect 24259 29053 24268 29087
rect 24216 29044 24268 29053
rect 27528 29044 27580 29096
rect 25320 28976 25372 29028
rect 27068 28976 27120 29028
rect 27344 28976 27396 29028
rect 31208 29112 31260 29164
rect 34520 29112 34572 29164
rect 35164 29112 35216 29164
rect 28632 29044 28684 29096
rect 28356 28976 28408 29028
rect 22468 28908 22520 28960
rect 22836 28951 22888 28960
rect 22836 28917 22845 28951
rect 22845 28917 22879 28951
rect 22879 28917 22888 28951
rect 22836 28908 22888 28917
rect 24032 28908 24084 28960
rect 24216 28908 24268 28960
rect 27712 28908 27764 28960
rect 35992 29180 36044 29232
rect 37556 29248 37608 29300
rect 37924 29291 37976 29300
rect 37924 29257 37933 29291
rect 37933 29257 37967 29291
rect 37967 29257 37976 29291
rect 37924 29248 37976 29257
rect 37464 29180 37516 29232
rect 36176 29112 36228 29164
rect 35992 29087 36044 29096
rect 35992 29053 36002 29087
rect 36002 29053 36036 29087
rect 36036 29053 36044 29087
rect 35992 29044 36044 29053
rect 37464 29087 37516 29096
rect 37464 29053 37473 29087
rect 37473 29053 37507 29087
rect 37507 29053 37516 29087
rect 37464 29044 37516 29053
rect 38108 29087 38160 29096
rect 38108 29053 38117 29087
rect 38117 29053 38151 29087
rect 38151 29053 38160 29087
rect 38108 29044 38160 29053
rect 36176 29019 36228 29028
rect 36176 28985 36185 29019
rect 36185 28985 36219 29019
rect 36219 28985 36228 29019
rect 36176 28976 36228 28985
rect 36452 28976 36504 29028
rect 35808 28908 35860 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 1676 28611 1728 28620
rect 1676 28577 1685 28611
rect 1685 28577 1719 28611
rect 1719 28577 1728 28611
rect 1676 28568 1728 28577
rect 2964 28568 3016 28620
rect 18328 28636 18380 28688
rect 17224 28568 17276 28620
rect 19984 28704 20036 28756
rect 20168 28704 20220 28756
rect 19248 28636 19300 28688
rect 22376 28704 22428 28756
rect 22652 28704 22704 28756
rect 23020 28704 23072 28756
rect 23388 28704 23440 28756
rect 26332 28704 26384 28756
rect 27160 28704 27212 28756
rect 33048 28704 33100 28756
rect 35900 28704 35952 28756
rect 36728 28704 36780 28756
rect 37188 28704 37240 28756
rect 32312 28636 32364 28688
rect 35072 28636 35124 28688
rect 36084 28636 36136 28688
rect 36268 28679 36320 28688
rect 36268 28645 36277 28679
rect 36277 28645 36311 28679
rect 36311 28645 36320 28679
rect 36268 28636 36320 28645
rect 19800 28611 19852 28620
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 18604 28432 18656 28484
rect 19800 28577 19809 28611
rect 19809 28577 19843 28611
rect 19843 28577 19852 28611
rect 19800 28568 19852 28577
rect 19984 28611 20036 28620
rect 19984 28577 19991 28611
rect 19991 28577 20036 28611
rect 19984 28568 20036 28577
rect 22560 28611 22612 28620
rect 19616 28432 19668 28484
rect 22560 28577 22569 28611
rect 22569 28577 22603 28611
rect 22603 28577 22612 28611
rect 22560 28568 22612 28577
rect 22468 28500 22520 28552
rect 23112 28568 23164 28620
rect 25044 28568 25096 28620
rect 36176 28611 36228 28620
rect 25044 28432 25096 28484
rect 19156 28364 19208 28416
rect 20812 28364 20864 28416
rect 24216 28364 24268 28416
rect 27528 28432 27580 28484
rect 28264 28432 28316 28484
rect 31944 28432 31996 28484
rect 35164 28432 35216 28484
rect 36176 28577 36185 28611
rect 36185 28577 36219 28611
rect 36219 28577 36228 28611
rect 36176 28568 36228 28577
rect 37188 28611 37240 28620
rect 36636 28500 36688 28552
rect 37188 28577 37197 28611
rect 37197 28577 37231 28611
rect 37231 28577 37240 28611
rect 37188 28568 37240 28577
rect 37372 28500 37424 28552
rect 37004 28432 37056 28484
rect 26608 28407 26660 28416
rect 26608 28373 26617 28407
rect 26617 28373 26651 28407
rect 26651 28373 26660 28407
rect 26608 28364 26660 28373
rect 29000 28364 29052 28416
rect 35256 28364 35308 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 2320 28160 2372 28212
rect 6368 28160 6420 28212
rect 21640 28160 21692 28212
rect 22100 28160 22152 28212
rect 18052 28092 18104 28144
rect 18788 28024 18840 28076
rect 24400 28092 24452 28144
rect 27160 28135 27212 28144
rect 26148 28067 26200 28076
rect 16028 27956 16080 28008
rect 18328 27888 18380 27940
rect 19156 27888 19208 27940
rect 5816 27820 5868 27872
rect 19984 27888 20036 27940
rect 20536 27888 20588 27940
rect 20260 27820 20312 27872
rect 22560 27956 22612 28008
rect 26148 28033 26157 28067
rect 26157 28033 26191 28067
rect 26191 28033 26200 28067
rect 26148 28024 26200 28033
rect 27160 28101 27169 28135
rect 27169 28101 27203 28135
rect 27203 28101 27212 28135
rect 27160 28092 27212 28101
rect 21272 27931 21324 27940
rect 21272 27897 21306 27931
rect 21306 27897 21324 27931
rect 21272 27888 21324 27897
rect 21456 27888 21508 27940
rect 22468 27888 22520 27940
rect 21640 27820 21692 27872
rect 22376 27863 22428 27872
rect 22376 27829 22385 27863
rect 22385 27829 22419 27863
rect 22419 27829 22428 27863
rect 22376 27820 22428 27829
rect 23112 27931 23164 27940
rect 23112 27897 23146 27931
rect 23146 27897 23164 27931
rect 23112 27888 23164 27897
rect 24676 27888 24728 27940
rect 26332 27956 26384 28008
rect 26884 27956 26936 28008
rect 28264 28024 28316 28076
rect 27252 27999 27304 28008
rect 27252 27965 27261 27999
rect 27261 27965 27295 27999
rect 27295 27965 27304 27999
rect 27252 27956 27304 27965
rect 27528 27999 27580 28008
rect 27528 27965 27537 27999
rect 27537 27965 27571 27999
rect 27571 27965 27580 27999
rect 27528 27956 27580 27965
rect 35900 27999 35952 28008
rect 35900 27965 35909 27999
rect 35909 27965 35943 27999
rect 35943 27965 35952 27999
rect 35900 27956 35952 27965
rect 36268 27999 36320 28008
rect 25780 27863 25832 27872
rect 25780 27829 25789 27863
rect 25789 27829 25823 27863
rect 25823 27829 25832 27863
rect 25780 27820 25832 27829
rect 26148 27820 26200 27872
rect 26884 27863 26936 27872
rect 26884 27829 26893 27863
rect 26893 27829 26927 27863
rect 26927 27829 26936 27863
rect 26884 27820 26936 27829
rect 27712 27888 27764 27940
rect 32680 27820 32732 27872
rect 36268 27965 36277 27999
rect 36277 27965 36311 27999
rect 36311 27965 36320 27999
rect 36268 27956 36320 27965
rect 36728 28160 36780 28212
rect 38476 28160 38528 28212
rect 36452 28092 36504 28144
rect 37464 27999 37516 28008
rect 37464 27965 37473 27999
rect 37473 27965 37507 27999
rect 37507 27965 37516 27999
rect 37464 27956 37516 27965
rect 37924 27999 37976 28008
rect 37924 27965 37933 27999
rect 37933 27965 37967 27999
rect 37967 27965 37976 27999
rect 37924 27956 37976 27965
rect 36176 27931 36228 27940
rect 36176 27897 36185 27931
rect 36185 27897 36219 27931
rect 36219 27897 36228 27931
rect 36176 27888 36228 27897
rect 37004 27820 37056 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 2964 27616 3016 27668
rect 18328 27616 18380 27668
rect 19248 27616 19300 27668
rect 20076 27616 20128 27668
rect 1860 27591 1912 27600
rect 1860 27557 1869 27591
rect 1869 27557 1903 27591
rect 1903 27557 1912 27591
rect 1860 27548 1912 27557
rect 2044 27591 2096 27600
rect 2044 27557 2053 27591
rect 2053 27557 2087 27591
rect 2087 27557 2096 27591
rect 2044 27548 2096 27557
rect 2780 27548 2832 27600
rect 10232 27548 10284 27600
rect 15292 27548 15344 27600
rect 20904 27616 20956 27668
rect 22376 27616 22428 27668
rect 20628 27548 20680 27600
rect 27068 27616 27120 27668
rect 27712 27616 27764 27668
rect 31668 27616 31720 27668
rect 36268 27616 36320 27668
rect 22652 27548 22704 27600
rect 24216 27548 24268 27600
rect 24492 27548 24544 27600
rect 2228 27480 2280 27532
rect 6276 27480 6328 27532
rect 8116 27480 8168 27532
rect 14924 27480 14976 27532
rect 20812 27480 20864 27532
rect 22100 27480 22152 27532
rect 25964 27523 26016 27532
rect 19984 27412 20036 27464
rect 20260 27455 20312 27464
rect 20260 27421 20269 27455
rect 20269 27421 20303 27455
rect 20303 27421 20312 27455
rect 20260 27412 20312 27421
rect 21640 27412 21692 27464
rect 24584 27412 24636 27464
rect 25964 27489 25973 27523
rect 25973 27489 26007 27523
rect 26007 27489 26016 27523
rect 25964 27480 26016 27489
rect 26148 27548 26200 27600
rect 31024 27548 31076 27600
rect 26332 27480 26384 27532
rect 26148 27412 26200 27464
rect 35900 27480 35952 27532
rect 36360 27480 36412 27532
rect 26884 27412 26936 27464
rect 27068 27412 27120 27464
rect 2136 27276 2188 27328
rect 2412 27276 2464 27328
rect 19616 27319 19668 27328
rect 19616 27285 19625 27319
rect 19625 27285 19659 27319
rect 19659 27285 19668 27319
rect 19616 27276 19668 27285
rect 23572 27344 23624 27396
rect 33968 27344 34020 27396
rect 21456 27276 21508 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 22468 27276 22520 27328
rect 22836 27276 22888 27328
rect 23940 27319 23992 27328
rect 23940 27285 23949 27319
rect 23949 27285 23983 27319
rect 23983 27285 23992 27319
rect 23940 27276 23992 27285
rect 24124 27276 24176 27328
rect 24676 27319 24728 27328
rect 24676 27285 24685 27319
rect 24685 27285 24719 27319
rect 24719 27285 24728 27319
rect 24676 27276 24728 27285
rect 25044 27319 25096 27328
rect 25044 27285 25053 27319
rect 25053 27285 25087 27319
rect 25087 27285 25096 27319
rect 25044 27276 25096 27285
rect 25320 27276 25372 27328
rect 26148 27276 26200 27328
rect 26884 27319 26936 27328
rect 26884 27285 26893 27319
rect 26893 27285 26927 27319
rect 26927 27285 26936 27319
rect 26884 27276 26936 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 21548 27072 21600 27124
rect 22928 27072 22980 27124
rect 25228 27072 25280 27124
rect 25872 27072 25924 27124
rect 36084 27072 36136 27124
rect 37832 27072 37884 27124
rect 2688 27004 2740 27056
rect 19984 26979 20036 26988
rect 19984 26945 19993 26979
rect 19993 26945 20027 26979
rect 20027 26945 20036 26979
rect 19984 26936 20036 26945
rect 21456 27004 21508 27056
rect 21732 27004 21784 27056
rect 23480 27004 23532 27056
rect 25596 26979 25648 26988
rect 20812 26868 20864 26920
rect 21824 26911 21876 26920
rect 21824 26877 21833 26911
rect 21833 26877 21867 26911
rect 21867 26877 21876 26911
rect 21824 26868 21876 26877
rect 22100 26911 22152 26920
rect 22100 26877 22134 26911
rect 22134 26877 22152 26911
rect 22100 26868 22152 26877
rect 22376 26868 22428 26920
rect 1860 26843 1912 26852
rect 1860 26809 1869 26843
rect 1869 26809 1903 26843
rect 1903 26809 1912 26843
rect 1860 26800 1912 26809
rect 20076 26800 20128 26852
rect 24676 26868 24728 26920
rect 25596 26945 25605 26979
rect 25605 26945 25639 26979
rect 25639 26945 25648 26979
rect 25596 26936 25648 26945
rect 30748 26936 30800 26988
rect 34612 26936 34664 26988
rect 35532 26936 35584 26988
rect 26884 26868 26936 26920
rect 37280 26911 37332 26920
rect 37280 26877 37289 26911
rect 37289 26877 37323 26911
rect 37323 26877 37332 26911
rect 37280 26868 37332 26877
rect 37924 26911 37976 26920
rect 37924 26877 37933 26911
rect 37933 26877 37967 26911
rect 37967 26877 37976 26911
rect 37924 26868 37976 26877
rect 24952 26800 25004 26852
rect 25320 26800 25372 26852
rect 25964 26800 26016 26852
rect 34152 26800 34204 26852
rect 35348 26800 35400 26852
rect 35532 26800 35584 26852
rect 21272 26732 21324 26784
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 25228 26775 25280 26784
rect 25228 26741 25237 26775
rect 25237 26741 25271 26775
rect 25271 26741 25280 26775
rect 25228 26732 25280 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 20076 26571 20128 26580
rect 20076 26537 20085 26571
rect 20085 26537 20119 26571
rect 20119 26537 20128 26571
rect 20076 26528 20128 26537
rect 24124 26528 24176 26580
rect 18604 26460 18656 26512
rect 20260 26460 20312 26512
rect 21640 26460 21692 26512
rect 25780 26460 25832 26512
rect 7932 26392 7984 26444
rect 20904 26324 20956 26376
rect 21824 26392 21876 26444
rect 22744 26392 22796 26444
rect 24400 26392 24452 26444
rect 22192 26324 22244 26376
rect 22560 26324 22612 26376
rect 22652 26256 22704 26308
rect 18880 26188 18932 26240
rect 19984 26188 20036 26240
rect 21272 26188 21324 26240
rect 26240 26392 26292 26444
rect 25044 26324 25096 26376
rect 26516 26299 26568 26308
rect 26516 26265 26525 26299
rect 26525 26265 26559 26299
rect 26559 26265 26568 26299
rect 26516 26256 26568 26265
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 2320 25916 2372 25968
rect 22652 25984 22704 26036
rect 24124 25984 24176 26036
rect 24308 25984 24360 26036
rect 1860 25823 1912 25832
rect 1860 25789 1869 25823
rect 1869 25789 1903 25823
rect 1903 25789 1912 25823
rect 1860 25780 1912 25789
rect 4804 25644 4856 25696
rect 14740 25780 14792 25832
rect 20812 25848 20864 25900
rect 21640 25780 21692 25832
rect 22560 25780 22612 25832
rect 26792 25984 26844 26036
rect 27344 25984 27396 26036
rect 36544 25984 36596 26036
rect 27528 25916 27580 25968
rect 33232 25916 33284 25968
rect 25044 25848 25096 25900
rect 25504 25823 25556 25832
rect 18236 25712 18288 25764
rect 18420 25755 18472 25764
rect 18420 25721 18429 25755
rect 18429 25721 18463 25755
rect 18463 25721 18472 25755
rect 18420 25712 18472 25721
rect 22192 25712 22244 25764
rect 25504 25789 25538 25823
rect 25538 25789 25556 25823
rect 25504 25780 25556 25789
rect 27528 25780 27580 25832
rect 27896 25780 27948 25832
rect 37280 25823 37332 25832
rect 37280 25789 37289 25823
rect 37289 25789 37323 25823
rect 37323 25789 37332 25823
rect 37280 25780 37332 25789
rect 37924 25823 37976 25832
rect 37924 25789 37933 25823
rect 37933 25789 37967 25823
rect 37967 25789 37976 25823
rect 37924 25780 37976 25789
rect 26976 25712 27028 25764
rect 23204 25644 23256 25696
rect 24124 25644 24176 25696
rect 28816 25644 28868 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 2044 25415 2096 25424
rect 2044 25381 2053 25415
rect 2053 25381 2087 25415
rect 2087 25381 2096 25415
rect 2044 25372 2096 25381
rect 1860 25347 1912 25356
rect 1860 25313 1869 25347
rect 1869 25313 1903 25347
rect 1903 25313 1912 25347
rect 1860 25304 1912 25313
rect 17776 25304 17828 25356
rect 18236 25415 18288 25424
rect 18236 25381 18245 25415
rect 18245 25381 18279 25415
rect 18279 25381 18288 25415
rect 18236 25372 18288 25381
rect 22192 25440 22244 25492
rect 18144 25347 18196 25356
rect 18144 25313 18153 25347
rect 18153 25313 18187 25347
rect 18187 25313 18196 25347
rect 18144 25304 18196 25313
rect 5632 25236 5684 25288
rect 18880 25304 18932 25356
rect 23296 25440 23348 25492
rect 23572 25372 23624 25424
rect 20812 25304 20864 25356
rect 21364 25347 21416 25356
rect 21364 25313 21373 25347
rect 21373 25313 21407 25347
rect 21407 25313 21416 25347
rect 21364 25304 21416 25313
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 20076 25168 20128 25220
rect 9404 25100 9456 25152
rect 20168 25100 20220 25152
rect 20904 25100 20956 25152
rect 24492 25440 24544 25492
rect 25044 25440 25096 25492
rect 31392 25440 31444 25492
rect 37648 25440 37700 25492
rect 24400 25372 24452 25424
rect 25136 25347 25188 25356
rect 25136 25313 25145 25347
rect 25145 25313 25179 25347
rect 25179 25313 25188 25347
rect 25136 25304 25188 25313
rect 26056 25347 26108 25356
rect 26056 25313 26065 25347
rect 26065 25313 26099 25347
rect 26099 25313 26108 25347
rect 26056 25304 26108 25313
rect 25964 25236 26016 25288
rect 26884 25304 26936 25356
rect 36820 25304 36872 25356
rect 37188 25347 37240 25356
rect 37188 25313 37197 25347
rect 37197 25313 37231 25347
rect 37231 25313 37240 25347
rect 37188 25304 37240 25313
rect 27712 25236 27764 25288
rect 35256 25236 35308 25288
rect 35440 25236 35492 25288
rect 24492 25168 24544 25220
rect 25044 25211 25096 25220
rect 24124 25100 24176 25152
rect 25044 25177 25053 25211
rect 25053 25177 25087 25211
rect 25087 25177 25096 25211
rect 25044 25168 25096 25177
rect 25136 25168 25188 25220
rect 34612 25168 34664 25220
rect 36728 25100 36780 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 16580 24896 16632 24948
rect 20904 24896 20956 24948
rect 1584 24828 1636 24880
rect 4896 24828 4948 24880
rect 15844 24760 15896 24812
rect 17224 24760 17276 24812
rect 23572 24896 23624 24948
rect 11796 24692 11848 24744
rect 17316 24735 17368 24744
rect 17316 24701 17330 24735
rect 17330 24701 17364 24735
rect 17364 24701 17368 24735
rect 17316 24692 17368 24701
rect 18420 24735 18472 24744
rect 18420 24701 18434 24735
rect 18434 24701 18468 24735
rect 18468 24701 18472 24735
rect 18420 24692 18472 24701
rect 19248 24692 19300 24744
rect 21272 24828 21324 24880
rect 22192 24760 22244 24812
rect 24032 24803 24084 24812
rect 24032 24769 24050 24803
rect 24050 24769 24084 24803
rect 24032 24760 24084 24769
rect 25044 24760 25096 24812
rect 28632 24828 28684 24880
rect 32036 24828 32088 24880
rect 21272 24692 21324 24744
rect 21548 24692 21600 24744
rect 22008 24692 22060 24744
rect 22284 24692 22336 24744
rect 17132 24667 17184 24676
rect 17132 24633 17141 24667
rect 17141 24633 17175 24667
rect 17175 24633 17184 24667
rect 17132 24624 17184 24633
rect 5724 24556 5776 24608
rect 17316 24556 17368 24608
rect 17408 24556 17460 24608
rect 17684 24624 17736 24676
rect 18144 24624 18196 24676
rect 18328 24667 18380 24676
rect 18328 24633 18337 24667
rect 18337 24633 18371 24667
rect 18371 24633 18380 24667
rect 18328 24624 18380 24633
rect 18512 24624 18564 24676
rect 20076 24667 20128 24676
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 20076 24633 20085 24667
rect 20085 24633 20119 24667
rect 20119 24633 20128 24667
rect 20076 24624 20128 24633
rect 21824 24624 21876 24676
rect 23848 24735 23900 24744
rect 23848 24701 23857 24735
rect 23857 24701 23891 24735
rect 23891 24701 23900 24735
rect 23848 24692 23900 24701
rect 25412 24735 25464 24744
rect 25412 24701 25421 24735
rect 25421 24701 25455 24735
rect 25455 24701 25464 24735
rect 25412 24692 25464 24701
rect 22744 24599 22796 24608
rect 22744 24565 22753 24599
rect 22753 24565 22787 24599
rect 22787 24565 22796 24599
rect 22744 24556 22796 24565
rect 23388 24556 23440 24608
rect 25780 24692 25832 24744
rect 30012 24760 30064 24812
rect 26884 24692 26936 24744
rect 37924 24735 37976 24744
rect 37924 24701 37933 24735
rect 37933 24701 37967 24735
rect 37967 24701 37976 24735
rect 37924 24692 37976 24701
rect 31300 24556 31352 24608
rect 38568 24556 38620 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 5540 24352 5592 24404
rect 18420 24352 18472 24404
rect 19248 24352 19300 24404
rect 23112 24352 23164 24404
rect 25780 24352 25832 24404
rect 29460 24352 29512 24404
rect 1860 24327 1912 24336
rect 1860 24293 1869 24327
rect 1869 24293 1903 24327
rect 1903 24293 1912 24327
rect 1860 24284 1912 24293
rect 2136 24284 2188 24336
rect 16672 24284 16724 24336
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18328 24284 18380 24336
rect 21640 24284 21692 24336
rect 23204 24284 23256 24336
rect 17684 24216 17736 24268
rect 2964 24148 3016 24200
rect 19984 24216 20036 24268
rect 20168 24216 20220 24268
rect 21456 24259 21508 24268
rect 21456 24225 21465 24259
rect 21465 24225 21499 24259
rect 21499 24225 21508 24259
rect 21456 24216 21508 24225
rect 24676 24259 24728 24268
rect 24676 24225 24685 24259
rect 24685 24225 24719 24259
rect 24719 24225 24728 24259
rect 24676 24216 24728 24225
rect 27252 24216 27304 24268
rect 1676 24080 1728 24132
rect 6552 24080 6604 24132
rect 21364 24148 21416 24200
rect 21548 24148 21600 24200
rect 22008 24148 22060 24200
rect 22744 24148 22796 24200
rect 24032 24148 24084 24200
rect 24308 24148 24360 24200
rect 37188 24259 37240 24268
rect 37188 24225 37197 24259
rect 37197 24225 37231 24259
rect 37231 24225 37240 24259
rect 37188 24216 37240 24225
rect 37556 24148 37608 24200
rect 17132 24080 17184 24132
rect 17684 24080 17736 24132
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 18420 24012 18472 24064
rect 19616 24012 19668 24064
rect 22560 24080 22612 24132
rect 27436 24080 27488 24132
rect 36636 24080 36688 24132
rect 22008 24012 22060 24064
rect 23572 24012 23624 24064
rect 31208 24012 31260 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 10508 23808 10560 23860
rect 18052 23808 18104 23860
rect 18144 23808 18196 23860
rect 27160 23808 27212 23860
rect 37372 23808 37424 23860
rect 38936 23808 38988 23860
rect 2228 23740 2280 23792
rect 19156 23740 19208 23792
rect 22100 23740 22152 23792
rect 25412 23740 25464 23792
rect 18604 23672 18656 23724
rect 28540 23672 28592 23724
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 18512 23647 18564 23656
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 19156 23604 19208 23656
rect 19800 23604 19852 23656
rect 19984 23647 20036 23656
rect 19984 23613 19993 23647
rect 19993 23613 20027 23647
rect 20027 23613 20036 23647
rect 19984 23604 20036 23613
rect 20720 23604 20772 23656
rect 20904 23604 20956 23656
rect 21456 23604 21508 23656
rect 21732 23604 21784 23656
rect 24676 23604 24728 23656
rect 37464 23647 37516 23656
rect 37464 23613 37473 23647
rect 37473 23613 37507 23647
rect 37507 23613 37516 23647
rect 37464 23604 37516 23613
rect 38108 23647 38160 23656
rect 38108 23613 38117 23647
rect 38117 23613 38151 23647
rect 38151 23613 38160 23647
rect 38108 23604 38160 23613
rect 17408 23536 17460 23588
rect 27528 23536 27580 23588
rect 20904 23468 20956 23520
rect 21456 23468 21508 23520
rect 23848 23468 23900 23520
rect 24308 23468 24360 23520
rect 25044 23468 25096 23520
rect 31944 23468 31996 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 13544 23264 13596 23316
rect 16120 23264 16172 23316
rect 17684 23307 17736 23316
rect 17684 23273 17693 23307
rect 17693 23273 17727 23307
rect 17727 23273 17736 23307
rect 17684 23264 17736 23273
rect 18328 23307 18380 23316
rect 18328 23273 18337 23307
rect 18337 23273 18371 23307
rect 18371 23273 18380 23307
rect 18328 23264 18380 23273
rect 19984 23264 20036 23316
rect 20628 23264 20680 23316
rect 20812 23264 20864 23316
rect 22008 23264 22060 23316
rect 23848 23264 23900 23316
rect 24400 23264 24452 23316
rect 27896 23264 27948 23316
rect 28908 23264 28960 23316
rect 34152 23264 34204 23316
rect 15936 23196 15988 23248
rect 16580 23196 16632 23248
rect 17500 23171 17552 23180
rect 17500 23137 17509 23171
rect 17509 23137 17543 23171
rect 17543 23137 17552 23171
rect 17500 23128 17552 23137
rect 18236 23128 18288 23180
rect 18512 23128 18564 23180
rect 20076 23128 20128 23180
rect 20812 23128 20864 23180
rect 21824 23128 21876 23180
rect 24124 23196 24176 23248
rect 25504 23196 25556 23248
rect 28540 23196 28592 23248
rect 27068 23128 27120 23180
rect 37188 23171 37240 23180
rect 37188 23137 37197 23171
rect 37197 23137 37231 23171
rect 37231 23137 37240 23171
rect 37188 23128 37240 23137
rect 9956 23060 10008 23112
rect 13176 23060 13228 23112
rect 18144 22992 18196 23044
rect 18512 22992 18564 23044
rect 20168 23060 20220 23112
rect 21456 23060 21508 23112
rect 22560 23103 22612 23112
rect 22560 23069 22569 23103
rect 22569 23069 22603 23103
rect 22603 23069 22612 23103
rect 22560 23060 22612 23069
rect 20628 22924 20680 22976
rect 22100 22924 22152 22976
rect 24584 22924 24636 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 18052 22652 18104 22704
rect 18880 22720 18932 22772
rect 22376 22720 22428 22772
rect 23112 22720 23164 22772
rect 18604 22695 18656 22704
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 13268 22516 13320 22568
rect 18144 22559 18196 22568
rect 18144 22525 18151 22559
rect 18151 22525 18196 22559
rect 18144 22516 18196 22525
rect 18604 22661 18613 22695
rect 18613 22661 18647 22695
rect 18647 22661 18656 22695
rect 18604 22652 18656 22661
rect 19156 22584 19208 22636
rect 23940 22720 23992 22772
rect 37740 22720 37792 22772
rect 38016 22720 38068 22772
rect 34520 22652 34572 22704
rect 1768 22448 1820 22500
rect 5816 22448 5868 22500
rect 7564 22448 7616 22500
rect 21456 22516 21508 22568
rect 23388 22516 23440 22568
rect 23572 22423 23624 22432
rect 23572 22389 23581 22423
rect 23581 22389 23615 22423
rect 23615 22389 23624 22423
rect 23572 22380 23624 22389
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 24400 22516 24452 22568
rect 37280 22559 37332 22568
rect 37280 22525 37289 22559
rect 37289 22525 37323 22559
rect 37323 22525 37332 22559
rect 37280 22516 37332 22525
rect 37924 22559 37976 22568
rect 37924 22525 37933 22559
rect 37933 22525 37967 22559
rect 37967 22525 37976 22559
rect 37924 22516 37976 22525
rect 34060 22448 34112 22500
rect 34612 22448 34664 22500
rect 24032 22380 24084 22432
rect 24216 22380 24268 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 14648 22176 14700 22228
rect 18604 22176 18656 22228
rect 23204 22176 23256 22228
rect 23848 22176 23900 22228
rect 24492 22176 24544 22228
rect 18880 22151 18932 22160
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 17776 22083 17828 22092
rect 17776 22049 17785 22083
rect 17785 22049 17819 22083
rect 17819 22049 17828 22083
rect 18880 22117 18889 22151
rect 18889 22117 18923 22151
rect 18923 22117 18932 22151
rect 18880 22108 18932 22117
rect 19156 22108 19208 22160
rect 17776 22040 17828 22049
rect 3608 21972 3660 22024
rect 17132 21972 17184 22024
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 1676 21904 1728 21956
rect 17960 21836 18012 21888
rect 18236 21836 18288 21888
rect 18880 21972 18932 22024
rect 20720 22108 20772 22160
rect 24400 22108 24452 22160
rect 20168 22083 20220 22092
rect 20168 22049 20177 22083
rect 20177 22049 20211 22083
rect 20211 22049 20220 22083
rect 20168 22040 20220 22049
rect 21364 22040 21416 22092
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 24676 22083 24728 22092
rect 24676 22049 24685 22083
rect 24685 22049 24719 22083
rect 24719 22049 24728 22083
rect 24676 22040 24728 22049
rect 24952 22015 25004 22024
rect 21456 21836 21508 21888
rect 21732 21836 21784 21888
rect 23204 21836 23256 21888
rect 23480 21836 23532 21888
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 24952 21981 24961 22015
rect 24961 21981 24995 22015
rect 24995 21981 25004 22015
rect 24952 21972 25004 21981
rect 37188 22083 37240 22092
rect 37188 22049 37197 22083
rect 37197 22049 37231 22083
rect 37231 22049 37240 22083
rect 37188 22040 37240 22049
rect 30472 21972 30524 22024
rect 35256 21904 35308 21956
rect 25228 21836 25280 21888
rect 28540 21836 28592 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 16856 21632 16908 21684
rect 10600 21564 10652 21616
rect 1676 21428 1728 21480
rect 5632 21428 5684 21480
rect 14832 21428 14884 21480
rect 16948 21471 17000 21480
rect 16948 21437 16955 21471
rect 16955 21437 17000 21471
rect 16948 21428 17000 21437
rect 17132 21471 17184 21480
rect 17132 21437 17141 21471
rect 17141 21437 17175 21471
rect 17175 21437 17184 21471
rect 17132 21428 17184 21437
rect 17408 21632 17460 21684
rect 18512 21675 18564 21684
rect 18052 21564 18104 21616
rect 18512 21641 18521 21675
rect 18521 21641 18555 21675
rect 18555 21641 18564 21675
rect 18512 21632 18564 21641
rect 18604 21632 18656 21684
rect 18880 21564 18932 21616
rect 21732 21632 21784 21684
rect 22284 21632 22336 21684
rect 35992 21632 36044 21684
rect 37096 21564 37148 21616
rect 20168 21496 20220 21548
rect 20628 21496 20680 21548
rect 22560 21496 22612 21548
rect 1584 21360 1636 21412
rect 14464 21360 14516 21412
rect 17040 21403 17092 21412
rect 17040 21369 17049 21403
rect 17049 21369 17083 21403
rect 17083 21369 17092 21403
rect 17040 21360 17092 21369
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 18328 21471 18380 21480
rect 18328 21437 18342 21471
rect 18342 21437 18376 21471
rect 18376 21437 18380 21471
rect 18328 21428 18380 21437
rect 18788 21428 18840 21480
rect 18512 21360 18564 21412
rect 19156 21360 19208 21412
rect 19984 21292 20036 21344
rect 22192 21428 22244 21480
rect 23848 21428 23900 21480
rect 37280 21471 37332 21480
rect 37280 21437 37289 21471
rect 37289 21437 37323 21471
rect 37323 21437 37332 21471
rect 37280 21428 37332 21437
rect 37924 21471 37976 21480
rect 37924 21437 37933 21471
rect 37933 21437 37967 21471
rect 37967 21437 37976 21471
rect 37924 21428 37976 21437
rect 21548 21360 21600 21412
rect 25964 21360 26016 21412
rect 32680 21360 32732 21412
rect 33416 21360 33468 21412
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 2688 21088 2740 21140
rect 17408 21088 17460 21140
rect 22100 21088 22152 21140
rect 22560 21088 22612 21140
rect 28172 21088 28224 21140
rect 17040 21020 17092 21072
rect 18052 21063 18104 21072
rect 18052 21029 18061 21063
rect 18061 21029 18095 21063
rect 18095 21029 18104 21063
rect 18052 21020 18104 21029
rect 18512 21020 18564 21072
rect 20812 21063 20864 21072
rect 20812 21029 20821 21063
rect 20821 21029 20855 21063
rect 20855 21029 20864 21063
rect 20812 21020 20864 21029
rect 23756 21020 23808 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 15292 20952 15344 21004
rect 17868 20995 17920 21004
rect 17868 20961 17878 20995
rect 17878 20961 17912 20995
rect 17912 20961 17920 20995
rect 17868 20952 17920 20961
rect 18236 20995 18288 21004
rect 18236 20961 18250 20995
rect 18250 20961 18284 20995
rect 18284 20961 18288 20995
rect 18236 20952 18288 20961
rect 6460 20884 6512 20936
rect 18328 20884 18380 20936
rect 22560 20952 22612 21004
rect 23480 20995 23532 21004
rect 23480 20961 23489 20995
rect 23489 20961 23523 20995
rect 23523 20961 23532 20995
rect 23480 20952 23532 20961
rect 24124 21020 24176 21072
rect 24400 21020 24452 21072
rect 24584 20995 24636 21004
rect 24584 20961 24593 20995
rect 24593 20961 24627 20995
rect 24627 20961 24636 20995
rect 24584 20952 24636 20961
rect 24768 20995 24820 21004
rect 24768 20961 24777 20995
rect 24777 20961 24811 20995
rect 24811 20961 24820 20995
rect 24768 20952 24820 20961
rect 21824 20884 21876 20936
rect 23848 20884 23900 20936
rect 19984 20816 20036 20868
rect 20628 20816 20680 20868
rect 17132 20748 17184 20800
rect 21364 20748 21416 20800
rect 24400 20791 24452 20800
rect 24400 20757 24409 20791
rect 24409 20757 24443 20791
rect 24443 20757 24452 20791
rect 24400 20748 24452 20757
rect 36452 20884 36504 20936
rect 35808 20748 35860 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 20536 20544 20588 20596
rect 23204 20544 23256 20596
rect 36820 20544 36872 20596
rect 18052 20476 18104 20528
rect 22836 20476 22888 20528
rect 35440 20476 35492 20528
rect 13452 20408 13504 20460
rect 16856 20408 16908 20460
rect 29644 20408 29696 20460
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 22560 20340 22612 20392
rect 21548 20272 21600 20324
rect 24124 20340 24176 20392
rect 37280 20383 37332 20392
rect 37280 20349 37289 20383
rect 37289 20349 37323 20383
rect 37323 20349 37332 20383
rect 37280 20340 37332 20349
rect 37924 20383 37976 20392
rect 37924 20349 37933 20383
rect 37933 20349 37967 20383
rect 37967 20349 37976 20383
rect 37924 20340 37976 20349
rect 16764 20204 16816 20256
rect 18236 20204 18288 20256
rect 20720 20204 20772 20256
rect 26240 20204 26292 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 7748 20000 7800 20052
rect 16580 20000 16632 20052
rect 1860 19932 1912 19984
rect 16764 19932 16816 19984
rect 6276 19796 6328 19848
rect 13176 19864 13228 19916
rect 17500 19932 17552 19984
rect 16488 19728 16540 19780
rect 17960 19932 18012 19984
rect 19524 19932 19576 19984
rect 20352 19932 20404 19984
rect 27804 19932 27856 19984
rect 36544 19932 36596 19984
rect 20352 19796 20404 19848
rect 19340 19728 19392 19780
rect 20536 19728 20588 19780
rect 16764 19660 16816 19712
rect 17500 19660 17552 19712
rect 28264 19660 28316 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 1584 19320 1636 19372
rect 5540 19320 5592 19372
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 1492 19252 1544 19304
rect 2964 19252 3016 19304
rect 16212 19295 16264 19304
rect 16764 19456 16816 19508
rect 18604 19456 18656 19508
rect 21732 19456 21784 19508
rect 16488 19388 16540 19440
rect 17316 19388 17368 19440
rect 16212 19261 16249 19295
rect 16249 19261 16264 19295
rect 16212 19252 16264 19261
rect 8944 19184 8996 19236
rect 1768 19116 1820 19168
rect 8668 19116 8720 19168
rect 13452 19116 13504 19168
rect 16028 19159 16080 19168
rect 16028 19125 16037 19159
rect 16037 19125 16071 19159
rect 16071 19125 16080 19159
rect 16028 19116 16080 19125
rect 17592 19388 17644 19440
rect 17224 19116 17276 19168
rect 17868 19252 17920 19304
rect 19432 19252 19484 19304
rect 19984 19295 20036 19304
rect 19984 19261 19993 19295
rect 19993 19261 20027 19295
rect 20027 19261 20036 19295
rect 19984 19252 20036 19261
rect 23572 19252 23624 19304
rect 26884 19252 26936 19304
rect 32772 19252 32824 19304
rect 37280 19295 37332 19304
rect 37280 19261 37289 19295
rect 37289 19261 37323 19295
rect 37323 19261 37332 19295
rect 37280 19252 37332 19261
rect 37924 19295 37976 19304
rect 37924 19261 37933 19295
rect 37933 19261 37967 19295
rect 37967 19261 37976 19295
rect 37924 19252 37976 19261
rect 18236 19184 18288 19236
rect 19248 19184 19300 19236
rect 24492 19184 24544 19236
rect 36912 19184 36964 19236
rect 17500 19116 17552 19168
rect 19984 19116 20036 19168
rect 20812 19116 20864 19168
rect 23296 19159 23348 19168
rect 23296 19125 23305 19159
rect 23305 19125 23339 19159
rect 23339 19125 23348 19159
rect 23296 19116 23348 19125
rect 31392 19116 31444 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 4804 18912 4856 18964
rect 16212 18912 16264 18964
rect 17868 18912 17920 18964
rect 18420 18912 18472 18964
rect 14464 18844 14516 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 15752 18819 15804 18828
rect 15752 18785 15761 18819
rect 15761 18785 15795 18819
rect 15795 18785 15804 18819
rect 15752 18776 15804 18785
rect 16028 18819 16080 18828
rect 16028 18785 16037 18819
rect 16037 18785 16071 18819
rect 16071 18785 16080 18819
rect 16028 18776 16080 18785
rect 16488 18776 16540 18828
rect 16856 18776 16908 18828
rect 17592 18819 17644 18828
rect 16764 18708 16816 18760
rect 17224 18708 17276 18760
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 18236 18844 18288 18896
rect 18604 18844 18656 18896
rect 19248 18912 19300 18964
rect 20628 18912 20680 18964
rect 20812 18912 20864 18964
rect 24952 18912 25004 18964
rect 37004 18912 37056 18964
rect 19984 18844 20036 18896
rect 25136 18844 25188 18896
rect 28172 18844 28224 18896
rect 29184 18844 29236 18896
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 17960 18708 18012 18760
rect 18328 18708 18380 18760
rect 18604 18708 18656 18760
rect 19432 18776 19484 18828
rect 20720 18776 20772 18828
rect 37188 18819 37240 18828
rect 37188 18785 37197 18819
rect 37197 18785 37231 18819
rect 37231 18785 37240 18819
rect 37188 18776 37240 18785
rect 19524 18640 19576 18692
rect 21640 18708 21692 18760
rect 27988 18708 28040 18760
rect 37004 18708 37056 18760
rect 21456 18640 21508 18692
rect 37648 18640 37700 18692
rect 21548 18572 21600 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 13268 18368 13320 18420
rect 17960 18368 18012 18420
rect 19340 18368 19392 18420
rect 20720 18368 20772 18420
rect 21548 18368 21600 18420
rect 23848 18368 23900 18420
rect 38200 18368 38252 18420
rect 4804 18232 4856 18284
rect 16580 18207 16632 18216
rect 16580 18173 16589 18207
rect 16589 18173 16623 18207
rect 16623 18173 16632 18207
rect 16580 18164 16632 18173
rect 16764 18207 16816 18216
rect 16764 18173 16771 18207
rect 16771 18173 16816 18207
rect 16764 18164 16816 18173
rect 17592 18300 17644 18352
rect 18236 18232 18288 18284
rect 19432 18232 19484 18284
rect 17776 18164 17828 18216
rect 18880 18207 18932 18216
rect 18880 18173 18889 18207
rect 18889 18173 18923 18207
rect 18923 18173 18932 18207
rect 18880 18164 18932 18173
rect 24400 18164 24452 18216
rect 21548 18028 21600 18080
rect 26056 18164 26108 18216
rect 37924 18207 37976 18216
rect 37924 18173 37933 18207
rect 37933 18173 37967 18207
rect 37967 18173 37976 18207
rect 37924 18164 37976 18173
rect 25412 18096 25464 18148
rect 28080 18096 28132 18148
rect 25320 18028 25372 18080
rect 27712 18028 27764 18080
rect 34428 18028 34480 18080
rect 36084 18028 36136 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 1676 17824 1728 17876
rect 7472 17824 7524 17876
rect 8392 17824 8444 17876
rect 17592 17799 17644 17808
rect 17592 17765 17601 17799
rect 17601 17765 17635 17799
rect 17635 17765 17644 17799
rect 17592 17756 17644 17765
rect 18328 17824 18380 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 1676 17688 1728 17740
rect 5724 17688 5776 17740
rect 11704 17688 11756 17740
rect 18236 17688 18288 17740
rect 19432 17688 19484 17740
rect 21364 17688 21416 17740
rect 22928 17756 22980 17808
rect 25964 17756 26016 17808
rect 28264 17824 28316 17876
rect 29092 17824 29144 17876
rect 32864 17824 32916 17876
rect 37464 17756 37516 17808
rect 24308 17688 24360 17740
rect 29644 17688 29696 17740
rect 33692 17688 33744 17740
rect 37188 17731 37240 17740
rect 37188 17697 37197 17731
rect 37197 17697 37231 17731
rect 37231 17697 37240 17731
rect 37188 17688 37240 17697
rect 17592 17620 17644 17672
rect 18420 17552 18472 17604
rect 9128 17484 9180 17536
rect 17316 17484 17368 17536
rect 18880 17484 18932 17536
rect 21732 17552 21784 17604
rect 21364 17484 21416 17536
rect 21824 17484 21876 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 14372 17280 14424 17332
rect 17592 17280 17644 17332
rect 21272 17323 21324 17332
rect 21272 17289 21281 17323
rect 21281 17289 21315 17323
rect 21315 17289 21324 17323
rect 21272 17280 21324 17289
rect 8300 17212 8352 17264
rect 16580 17212 16632 17264
rect 16764 17212 16816 17264
rect 2044 17144 2096 17196
rect 4804 17144 4856 17196
rect 17500 17144 17552 17196
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 20904 17076 20956 17128
rect 23388 17144 23440 17196
rect 21732 17119 21784 17128
rect 21732 17085 21767 17119
rect 21767 17085 21784 17119
rect 21732 17076 21784 17085
rect 19340 17008 19392 17060
rect 22468 17008 22520 17060
rect 23020 17008 23072 17060
rect 36728 17280 36780 17332
rect 34336 17212 34388 17264
rect 37096 17144 37148 17196
rect 37280 17119 37332 17128
rect 37280 17085 37289 17119
rect 37289 17085 37323 17119
rect 37323 17085 37332 17119
rect 37280 17076 37332 17085
rect 37924 17119 37976 17128
rect 37924 17085 37933 17119
rect 37933 17085 37967 17119
rect 37967 17085 37976 17119
rect 37924 17076 37976 17085
rect 37372 17008 37424 17060
rect 20904 16940 20956 16992
rect 21456 16940 21508 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 13452 16736 13504 16788
rect 18604 16736 18656 16788
rect 20076 16736 20128 16788
rect 21364 16736 21416 16788
rect 22928 16736 22980 16788
rect 28356 16736 28408 16788
rect 37004 16736 37056 16788
rect 5816 16668 5868 16720
rect 9404 16668 9456 16720
rect 24308 16600 24360 16652
rect 28448 16600 28500 16652
rect 37188 16643 37240 16652
rect 37188 16609 37197 16643
rect 37197 16609 37231 16643
rect 37231 16609 37240 16643
rect 37188 16600 37240 16609
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 1492 16192 1544 16244
rect 22008 16192 22060 16244
rect 24032 16124 24084 16176
rect 35532 16192 35584 16244
rect 32220 16124 32272 16176
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 16580 16031 16632 16040
rect 16580 15997 16589 16031
rect 16589 15997 16623 16031
rect 16623 15997 16632 16031
rect 16580 15988 16632 15997
rect 37832 16056 37884 16108
rect 1768 15920 1820 15972
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 17132 15920 17184 15972
rect 35256 15988 35308 16040
rect 37280 16031 37332 16040
rect 37280 15997 37289 16031
rect 37289 15997 37323 16031
rect 37323 15997 37332 16031
rect 37280 15988 37332 15997
rect 37924 16031 37976 16040
rect 37924 15997 37933 16031
rect 37933 15997 37967 16031
rect 37967 15997 37976 16031
rect 37924 15988 37976 15997
rect 18420 15920 18472 15972
rect 36176 15920 36228 15972
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 1676 15648 1728 15700
rect 8208 15648 8260 15700
rect 12348 15580 12400 15632
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 14924 15512 14976 15564
rect 15844 15555 15896 15564
rect 15844 15521 15854 15555
rect 15854 15521 15888 15555
rect 15888 15521 15896 15555
rect 15844 15512 15896 15521
rect 17132 15580 17184 15632
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 17500 15555 17552 15564
rect 17500 15521 17507 15555
rect 17507 15521 17552 15555
rect 17500 15512 17552 15521
rect 17592 15555 17644 15564
rect 17592 15521 17601 15555
rect 17601 15521 17635 15555
rect 17635 15521 17644 15555
rect 24676 15648 24728 15700
rect 36544 15648 36596 15700
rect 17592 15512 17644 15521
rect 37188 15555 37240 15564
rect 37188 15521 37197 15555
rect 37197 15521 37231 15555
rect 37231 15521 37240 15555
rect 37188 15512 37240 15521
rect 16856 15444 16908 15496
rect 24584 15376 24636 15428
rect 16856 15308 16908 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 8392 14968 8444 15020
rect 17684 15036 17736 15088
rect 22560 15104 22612 15156
rect 35624 15104 35676 15156
rect 23480 15036 23532 15088
rect 35716 15036 35768 15088
rect 14556 14900 14608 14952
rect 16580 14943 16632 14952
rect 16580 14909 16590 14943
rect 16590 14909 16624 14943
rect 16624 14909 16632 14943
rect 16764 14943 16816 14952
rect 16580 14900 16632 14909
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 17040 14900 17092 14952
rect 17684 14943 17736 14952
rect 17684 14909 17694 14943
rect 17694 14909 17728 14943
rect 17728 14909 17736 14943
rect 19156 14968 19208 15020
rect 24952 14968 25004 15020
rect 17684 14900 17736 14909
rect 18052 14943 18104 14952
rect 18052 14909 18066 14943
rect 18066 14909 18100 14943
rect 18100 14909 18104 14943
rect 37280 14943 37332 14952
rect 18052 14900 18104 14909
rect 37280 14909 37289 14943
rect 37289 14909 37323 14943
rect 37323 14909 37332 14943
rect 37280 14900 37332 14909
rect 37924 14943 37976 14952
rect 37924 14909 37933 14943
rect 37933 14909 37967 14943
rect 37967 14909 37976 14943
rect 37924 14900 37976 14909
rect 3516 14764 3568 14816
rect 17132 14832 17184 14884
rect 17040 14764 17092 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 7564 14560 7616 14612
rect 19984 14560 20036 14612
rect 37280 14560 37332 14612
rect 16028 14492 16080 14544
rect 38016 14492 38068 14544
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 16580 14424 16632 14476
rect 24860 14424 24912 14476
rect 25872 14424 25924 14476
rect 6368 14356 6420 14408
rect 18052 14356 18104 14408
rect 34520 14220 34572 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 3608 14016 3660 14068
rect 32496 14016 32548 14068
rect 25964 13948 26016 14000
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 37188 13855 37240 13864
rect 37188 13821 37197 13855
rect 37197 13821 37231 13855
rect 37231 13821 37240 13855
rect 37188 13812 37240 13821
rect 37924 13855 37976 13864
rect 37924 13821 37933 13855
rect 37933 13821 37967 13855
rect 37967 13821 37976 13855
rect 37924 13812 37976 13821
rect 15292 13744 15344 13796
rect 16396 13744 16448 13796
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 21824 13472 21876 13524
rect 26332 13472 26384 13524
rect 37188 13379 37240 13388
rect 37188 13345 37197 13379
rect 37197 13345 37231 13379
rect 37231 13345 37240 13379
rect 37188 13336 37240 13345
rect 10416 13268 10468 13320
rect 19340 13268 19392 13320
rect 17868 13200 17920 13252
rect 36912 13200 36964 13252
rect 1768 13132 1820 13184
rect 14372 13132 14424 13184
rect 21916 13132 21968 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 6460 12928 6512 12980
rect 29736 12928 29788 12980
rect 20720 12792 20772 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 20628 12724 20680 12776
rect 16396 12656 16448 12708
rect 21732 12699 21784 12708
rect 21732 12665 21741 12699
rect 21741 12665 21775 12699
rect 21775 12665 21784 12699
rect 21732 12656 21784 12665
rect 37924 12699 37976 12708
rect 37924 12665 37933 12699
rect 37933 12665 37967 12699
rect 37967 12665 37976 12699
rect 37924 12656 37976 12665
rect 20536 12588 20588 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 1860 12384 1912 12436
rect 36636 12384 36688 12436
rect 19892 12316 19944 12368
rect 20536 12316 20588 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 37188 12291 37240 12300
rect 37188 12257 37197 12291
rect 37197 12257 37231 12291
rect 37231 12257 37240 12291
rect 37188 12248 37240 12257
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 10232 11840 10284 11892
rect 20812 11840 20864 11892
rect 31116 11840 31168 11892
rect 17500 11772 17552 11824
rect 36268 11772 36320 11824
rect 4068 11704 4120 11756
rect 10508 11704 10560 11756
rect 16120 11704 16172 11756
rect 36728 11704 36780 11756
rect 37188 11679 37240 11688
rect 37188 11645 37197 11679
rect 37197 11645 37231 11679
rect 37231 11645 37240 11679
rect 37188 11636 37240 11645
rect 37924 11611 37976 11620
rect 37924 11577 37933 11611
rect 37933 11577 37967 11611
rect 37967 11577 37976 11611
rect 37924 11568 37976 11577
rect 18972 11500 19024 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 37188 11203 37240 11212
rect 37188 11169 37197 11203
rect 37197 11169 37231 11203
rect 37231 11169 37240 11203
rect 37188 11160 37240 11169
rect 17132 11092 17184 11144
rect 19892 11092 19944 11144
rect 20260 11092 20312 11144
rect 10600 11024 10652 11076
rect 12900 11024 12952 11076
rect 18788 11024 18840 11076
rect 21732 11024 21784 11076
rect 25964 11024 26016 11076
rect 2228 10956 2280 11008
rect 8208 10956 8260 11008
rect 16672 10956 16724 11008
rect 24768 10956 24820 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 14832 10548 14884 10600
rect 23112 10548 23164 10600
rect 17224 10480 17276 10532
rect 37740 10480 37792 10532
rect 37924 10523 37976 10532
rect 37924 10489 37933 10523
rect 37933 10489 37967 10523
rect 37967 10489 37976 10523
rect 37924 10480 37976 10489
rect 9404 10412 9456 10464
rect 20076 10412 20128 10464
rect 23204 10412 23256 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 37188 10115 37240 10124
rect 37188 10081 37197 10115
rect 37197 10081 37231 10115
rect 37231 10081 37240 10115
rect 37188 10072 37240 10081
rect 16212 9868 16264 9920
rect 24952 9868 25004 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 22928 9664 22980 9716
rect 26700 9664 26752 9716
rect 18236 9596 18288 9648
rect 23296 9596 23348 9648
rect 37556 9596 37608 9648
rect 37832 9596 37884 9648
rect 16948 9528 17000 9580
rect 23112 9528 23164 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 37188 9503 37240 9512
rect 37188 9469 37197 9503
rect 37197 9469 37231 9503
rect 37231 9469 37240 9503
rect 37188 9460 37240 9469
rect 37924 9435 37976 9444
rect 37924 9401 37933 9435
rect 37933 9401 37967 9435
rect 37967 9401 37976 9435
rect 37924 9392 37976 9401
rect 13268 9324 13320 9376
rect 17684 9324 17736 9376
rect 26884 9324 26936 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 15844 9120 15896 9172
rect 6920 8916 6972 8968
rect 21548 8916 21600 8968
rect 25872 9120 25924 9172
rect 31208 9120 31260 9172
rect 23388 9095 23440 9104
rect 23388 9061 23397 9095
rect 23397 9061 23431 9095
rect 23431 9061 23440 9095
rect 23388 9052 23440 9061
rect 26884 9052 26936 9104
rect 37556 9052 37608 9104
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 23020 9027 23072 9036
rect 23020 8993 23029 9027
rect 23029 8993 23063 9027
rect 23063 8993 23072 9027
rect 23020 8984 23072 8993
rect 25596 8984 25648 9036
rect 37188 9027 37240 9036
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 37832 8916 37884 8968
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 10784 8372 10836 8424
rect 19156 8372 19208 8424
rect 24768 8372 24820 8424
rect 13452 8304 13504 8356
rect 37924 8347 37976 8356
rect 37924 8313 37933 8347
rect 37933 8313 37967 8347
rect 37967 8313 37976 8347
rect 37924 8304 37976 8313
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 2044 8032 2096 8084
rect 2320 8032 2372 8084
rect 6276 8032 6328 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 37188 7939 37240 7948
rect 37188 7905 37197 7939
rect 37197 7905 37231 7939
rect 37231 7905 37240 7939
rect 37188 7896 37240 7905
rect 1584 7828 1636 7880
rect 12348 7828 12400 7880
rect 15016 7828 15068 7880
rect 23940 7828 23992 7880
rect 10968 7760 11020 7812
rect 23204 7760 23256 7812
rect 24860 7760 24912 7812
rect 36452 7760 36504 7812
rect 17408 7692 17460 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 20628 7488 20680 7540
rect 22468 7488 22520 7540
rect 26608 7488 26660 7540
rect 37648 7488 37700 7540
rect 16856 7327 16908 7336
rect 16856 7293 16865 7327
rect 16865 7293 16899 7327
rect 16899 7293 16908 7327
rect 16856 7284 16908 7293
rect 37188 7327 37240 7336
rect 37188 7293 37197 7327
rect 37197 7293 37231 7327
rect 37231 7293 37240 7327
rect 37188 7284 37240 7293
rect 37924 7259 37976 7268
rect 37924 7225 37933 7259
rect 37933 7225 37967 7259
rect 37967 7225 37976 7259
rect 37924 7216 37976 7225
rect 23296 7148 23348 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 20076 6944 20128 6996
rect 26516 6944 26568 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 13084 6808 13136 6860
rect 17316 6808 17368 6860
rect 35256 6808 35308 6860
rect 36544 6808 36596 6860
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 37280 6808 37332 6860
rect 15200 6740 15252 6792
rect 21272 6740 21324 6792
rect 1768 6672 1820 6724
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 1676 6400 1728 6452
rect 37096 6400 37148 6452
rect 18880 6332 18932 6384
rect 27344 6332 27396 6384
rect 36912 6332 36964 6384
rect 2504 6264 2556 6316
rect 14464 6264 14516 6316
rect 14924 6264 14976 6316
rect 22284 6264 22336 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 20352 6196 20404 6248
rect 5080 6128 5132 6180
rect 20168 6128 20220 6180
rect 36360 6128 36412 6180
rect 37004 6128 37056 6180
rect 37096 6128 37148 6180
rect 37924 6171 37976 6180
rect 37924 6137 37933 6171
rect 37933 6137 37967 6171
rect 37967 6137 37976 6171
rect 37924 6128 37976 6137
rect 37280 6060 37332 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 3516 5856 3568 5908
rect 28356 5788 28408 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 2136 5720 2188 5772
rect 30564 5720 30616 5772
rect 37188 5763 37240 5772
rect 37188 5729 37197 5763
rect 37197 5729 37231 5763
rect 37231 5729 37240 5763
rect 37188 5720 37240 5729
rect 4988 5652 5040 5704
rect 5540 5652 5592 5704
rect 23112 5584 23164 5636
rect 4896 5516 4948 5568
rect 13360 5516 13412 5568
rect 15752 5516 15804 5568
rect 17408 5516 17460 5568
rect 24216 5516 24268 5568
rect 35624 5516 35676 5568
rect 36084 5516 36136 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 6368 5312 6420 5364
rect 28908 5312 28960 5364
rect 29552 5312 29604 5364
rect 36544 5355 36596 5364
rect 36544 5321 36553 5355
rect 36553 5321 36587 5355
rect 36587 5321 36596 5355
rect 36544 5312 36596 5321
rect 37740 5312 37792 5364
rect 37372 5287 37424 5296
rect 37372 5253 37381 5287
rect 37381 5253 37415 5287
rect 37415 5253 37424 5287
rect 37372 5244 37424 5253
rect 34612 5176 34664 5228
rect 35532 5176 35584 5228
rect 1308 5108 1360 5160
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 31300 5108 31352 5160
rect 36912 5108 36964 5160
rect 37188 5151 37240 5160
rect 37188 5117 37197 5151
rect 37197 5117 37231 5151
rect 37231 5117 37240 5151
rect 37188 5108 37240 5117
rect 6184 5040 6236 5092
rect 12440 5040 12492 5092
rect 31760 5040 31812 5092
rect 34612 5083 34664 5092
rect 34612 5049 34621 5083
rect 34621 5049 34655 5083
rect 34655 5049 34664 5083
rect 34612 5040 34664 5049
rect 36636 5040 36688 5092
rect 37924 5083 37976 5092
rect 37924 5049 37933 5083
rect 37933 5049 37967 5083
rect 37967 5049 37976 5083
rect 37924 5040 37976 5049
rect 11704 4972 11756 5024
rect 22192 4972 22244 5024
rect 33600 4972 33652 5024
rect 38936 4972 38988 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 9588 4768 9640 4820
rect 20904 4768 20956 4820
rect 36268 4768 36320 4820
rect 25964 4700 26016 4752
rect 34520 4700 34572 4752
rect 36176 4700 36228 4752
rect 37464 4700 37516 4752
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 22284 4632 22336 4684
rect 22652 4564 22704 4616
rect 25136 4632 25188 4684
rect 26608 4632 26660 4684
rect 30196 4632 30248 4684
rect 31024 4632 31076 4684
rect 33232 4632 33284 4684
rect 35808 4632 35860 4684
rect 36544 4632 36596 4684
rect 37188 4675 37240 4684
rect 37188 4641 37197 4675
rect 37197 4641 37231 4675
rect 37231 4641 37240 4675
rect 37188 4632 37240 4641
rect 36268 4564 36320 4616
rect 33324 4496 33376 4548
rect 1124 4428 1176 4480
rect 2044 4428 2096 4480
rect 2964 4428 3016 4480
rect 8944 4428 8996 4480
rect 20720 4428 20772 4480
rect 22560 4471 22612 4480
rect 22560 4437 22569 4471
rect 22569 4437 22603 4471
rect 22603 4437 22612 4471
rect 22560 4428 22612 4437
rect 25228 4471 25280 4480
rect 25228 4437 25237 4471
rect 25237 4437 25271 4471
rect 25271 4437 25280 4471
rect 25228 4428 25280 4437
rect 26240 4428 26292 4480
rect 29736 4428 29788 4480
rect 31392 4471 31444 4480
rect 31392 4437 31401 4471
rect 31401 4437 31435 4471
rect 31435 4437 31444 4471
rect 31392 4428 31444 4437
rect 35440 4428 35492 4480
rect 36176 4428 36228 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 1952 4088 2004 4140
rect 21180 4224 21232 4276
rect 22376 4224 22428 4276
rect 25228 4224 25280 4276
rect 32496 4224 32548 4276
rect 20720 4156 20772 4208
rect 23940 4199 23992 4208
rect 2044 4020 2096 4072
rect 2596 4063 2648 4072
rect 2596 4029 2605 4063
rect 2605 4029 2639 4063
rect 2639 4029 2648 4063
rect 2596 4020 2648 4029
rect 14740 4088 14792 4140
rect 23940 4165 23949 4199
rect 23949 4165 23983 4199
rect 23983 4165 23992 4199
rect 23940 4156 23992 4165
rect 28540 4199 28592 4208
rect 28540 4165 28549 4199
rect 28549 4165 28583 4199
rect 28583 4165 28592 4199
rect 28540 4156 28592 4165
rect 33048 4156 33100 4208
rect 1492 3952 1544 4004
rect 3608 3952 3660 4004
rect 4804 3952 4856 4004
rect 5908 4020 5960 4072
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 8944 3952 8996 4004
rect 940 3884 992 3936
rect 4896 3884 4948 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 10600 3884 10652 3936
rect 11428 3884 11480 3936
rect 15016 4063 15068 4072
rect 15016 4029 15025 4063
rect 15025 4029 15059 4063
rect 15059 4029 15068 4063
rect 15936 4063 15988 4072
rect 15016 4020 15068 4029
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 17868 4020 17920 4072
rect 19432 4020 19484 4072
rect 20536 4020 20588 4072
rect 21364 4020 21416 4072
rect 23296 4063 23348 4072
rect 15384 3952 15436 4004
rect 23296 4029 23305 4063
rect 23305 4029 23339 4063
rect 23339 4029 23348 4063
rect 23296 4020 23348 4029
rect 23112 3952 23164 4004
rect 24860 4020 24912 4072
rect 25780 4020 25832 4072
rect 30288 4088 30340 4140
rect 30380 4088 30432 4140
rect 34336 4156 34388 4208
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15844 3884 15896 3936
rect 17592 3884 17644 3936
rect 17960 3884 18012 3936
rect 20628 3927 20680 3936
rect 20628 3893 20637 3927
rect 20637 3893 20671 3927
rect 20671 3893 20680 3927
rect 20628 3884 20680 3893
rect 22100 3884 22152 3936
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 23388 3884 23440 3936
rect 27160 3952 27212 4004
rect 27436 4020 27488 4072
rect 28356 4020 28408 4072
rect 29276 4020 29328 4072
rect 28540 3952 28592 4004
rect 30564 4020 30616 4072
rect 30840 4063 30892 4072
rect 30840 4029 30849 4063
rect 30849 4029 30883 4063
rect 30883 4029 30892 4063
rect 30840 4020 30892 4029
rect 32496 4063 32548 4072
rect 32496 4029 32505 4063
rect 32505 4029 32539 4063
rect 32539 4029 32548 4063
rect 32496 4020 32548 4029
rect 25228 3927 25280 3936
rect 25228 3893 25237 3927
rect 25237 3893 25271 3927
rect 25271 3893 25280 3927
rect 25228 3884 25280 3893
rect 26516 3884 26568 3936
rect 27344 3927 27396 3936
rect 27344 3893 27353 3927
rect 27353 3893 27387 3927
rect 27387 3893 27396 3927
rect 27344 3884 27396 3893
rect 27896 3927 27948 3936
rect 27896 3893 27905 3927
rect 27905 3893 27939 3927
rect 27939 3893 27948 3927
rect 27896 3884 27948 3893
rect 27988 3884 28040 3936
rect 30472 3952 30524 4004
rect 29552 3884 29604 3936
rect 30748 3884 30800 3936
rect 31576 3884 31628 3936
rect 33232 4020 33284 4072
rect 36360 4088 36412 4140
rect 36452 4088 36504 4140
rect 37556 4088 37608 4140
rect 37832 4088 37884 4140
rect 34520 4063 34572 4072
rect 34520 4029 34529 4063
rect 34529 4029 34563 4063
rect 34563 4029 34572 4063
rect 34520 4020 34572 4029
rect 33324 3952 33376 4004
rect 33600 3952 33652 4004
rect 36268 4020 36320 4072
rect 39488 4020 39540 4072
rect 36452 3995 36504 4004
rect 36452 3961 36461 3995
rect 36461 3961 36495 3995
rect 36495 3961 36504 3995
rect 36452 3952 36504 3961
rect 36820 3952 36872 4004
rect 38108 3952 38160 4004
rect 33232 3927 33284 3936
rect 33232 3893 33241 3927
rect 33241 3893 33275 3927
rect 33275 3893 33284 3927
rect 33232 3884 33284 3893
rect 34612 3884 34664 3936
rect 35348 3884 35400 3936
rect 36912 3884 36964 3936
rect 37464 3884 37516 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 2320 3680 2372 3732
rect 2412 3680 2464 3732
rect 3424 3723 3476 3732
rect 3056 3612 3108 3664
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 8760 3723 8812 3732
rect 4068 3655 4120 3664
rect 4068 3621 4077 3655
rect 4077 3621 4111 3655
rect 4111 3621 4120 3655
rect 4068 3612 4120 3621
rect 6920 3655 6972 3664
rect 6920 3621 6929 3655
rect 6929 3621 6963 3655
rect 6963 3621 6972 3655
rect 6920 3612 6972 3621
rect 2964 3476 3016 3528
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 5356 3544 5408 3596
rect 7380 3544 7432 3596
rect 3332 3476 3384 3528
rect 8760 3689 8769 3723
rect 8769 3689 8803 3723
rect 8803 3689 8812 3723
rect 8760 3680 8812 3689
rect 11060 3723 11112 3732
rect 11060 3689 11069 3723
rect 11069 3689 11103 3723
rect 11103 3689 11112 3723
rect 11060 3680 11112 3689
rect 12256 3723 12308 3732
rect 12256 3689 12265 3723
rect 12265 3689 12299 3723
rect 12299 3689 12308 3723
rect 12256 3680 12308 3689
rect 16304 3723 16356 3732
rect 16304 3689 16313 3723
rect 16313 3689 16347 3723
rect 16347 3689 16356 3723
rect 16304 3680 16356 3689
rect 9404 3655 9456 3664
rect 9404 3621 9413 3655
rect 9413 3621 9447 3655
rect 9447 3621 9456 3655
rect 9404 3612 9456 3621
rect 10232 3612 10284 3664
rect 12900 3655 12952 3664
rect 12900 3621 12909 3655
rect 12909 3621 12943 3655
rect 12943 3621 12952 3655
rect 12900 3612 12952 3621
rect 14004 3612 14056 3664
rect 14556 3612 14608 3664
rect 19984 3680 20036 3732
rect 20444 3680 20496 3732
rect 17408 3655 17460 3664
rect 17408 3621 17417 3655
rect 17417 3621 17451 3655
rect 17451 3621 17460 3655
rect 17408 3612 17460 3621
rect 18144 3655 18196 3664
rect 18144 3621 18153 3655
rect 18153 3621 18187 3655
rect 18187 3621 18196 3655
rect 18144 3612 18196 3621
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 11060 3544 11112 3596
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 16028 3544 16080 3596
rect 16396 3544 16448 3596
rect 15384 3476 15436 3528
rect 18880 3587 18932 3596
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 23296 3680 23348 3732
rect 22192 3612 22244 3664
rect 26148 3680 26200 3732
rect 26792 3680 26844 3732
rect 33508 3723 33560 3732
rect 24308 3612 24360 3664
rect 24400 3612 24452 3664
rect 25412 3655 25464 3664
rect 22928 3587 22980 3596
rect 18788 3476 18840 3528
rect 16856 3408 16908 3460
rect 16948 3408 17000 3460
rect 22192 3476 22244 3528
rect 22928 3553 22937 3587
rect 22937 3553 22971 3587
rect 22971 3553 22980 3587
rect 22928 3544 22980 3553
rect 23756 3544 23808 3596
rect 24032 3544 24084 3596
rect 25412 3621 25421 3655
rect 25421 3621 25455 3655
rect 25455 3621 25464 3655
rect 25412 3612 25464 3621
rect 27988 3612 28040 3664
rect 28264 3612 28316 3664
rect 28908 3655 28960 3664
rect 28908 3621 28917 3655
rect 28917 3621 28951 3655
rect 28951 3621 28960 3655
rect 28908 3612 28960 3621
rect 26056 3587 26108 3596
rect 26056 3553 26065 3587
rect 26065 3553 26099 3587
rect 26099 3553 26108 3587
rect 26056 3544 26108 3553
rect 26148 3544 26200 3596
rect 30380 3612 30432 3664
rect 30472 3655 30524 3664
rect 30472 3621 30481 3655
rect 30481 3621 30515 3655
rect 30515 3621 30524 3655
rect 30472 3612 30524 3621
rect 30656 3612 30708 3664
rect 29552 3587 29604 3596
rect 29552 3553 29561 3587
rect 29561 3553 29595 3587
rect 29595 3553 29604 3587
rect 29552 3544 29604 3553
rect 29736 3544 29788 3596
rect 30564 3544 30616 3596
rect 33508 3689 33517 3723
rect 33517 3689 33551 3723
rect 33551 3689 33560 3723
rect 33508 3680 33560 3689
rect 34244 3723 34296 3732
rect 34244 3689 34253 3723
rect 34253 3689 34287 3723
rect 34287 3689 34296 3723
rect 34244 3680 34296 3689
rect 34796 3680 34848 3732
rect 35900 3723 35952 3732
rect 35900 3689 35909 3723
rect 35909 3689 35943 3723
rect 35943 3689 35952 3723
rect 35900 3680 35952 3689
rect 36728 3680 36780 3732
rect 31484 3612 31536 3664
rect 34336 3612 34388 3664
rect 34612 3612 34664 3664
rect 36912 3612 36964 3664
rect 33324 3587 33376 3596
rect 33324 3553 33333 3587
rect 33333 3553 33367 3587
rect 33367 3553 33376 3587
rect 33324 3544 33376 3553
rect 33968 3544 34020 3596
rect 34244 3544 34296 3596
rect 35716 3587 35768 3596
rect 35716 3553 35725 3587
rect 35725 3553 35759 3587
rect 35759 3553 35768 3587
rect 35716 3544 35768 3553
rect 37188 3587 37240 3596
rect 37188 3553 37197 3587
rect 37197 3553 37231 3587
rect 37231 3553 37240 3587
rect 37188 3544 37240 3553
rect 23388 3476 23440 3528
rect 33048 3476 33100 3528
rect 33232 3476 33284 3528
rect 39212 3476 39264 3528
rect 3240 3340 3292 3392
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 6828 3340 6880 3392
rect 8852 3340 8904 3392
rect 9680 3340 9732 3392
rect 12348 3340 12400 3392
rect 14096 3340 14148 3392
rect 16672 3340 16724 3392
rect 17684 3340 17736 3392
rect 18512 3340 18564 3392
rect 19524 3383 19576 3392
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 19984 3340 20036 3392
rect 27344 3408 27396 3460
rect 22836 3340 22888 3392
rect 23756 3340 23808 3392
rect 24492 3383 24544 3392
rect 24492 3349 24501 3383
rect 24501 3349 24535 3383
rect 24535 3349 24544 3383
rect 24492 3340 24544 3349
rect 25504 3383 25556 3392
rect 25504 3349 25513 3383
rect 25513 3349 25547 3383
rect 25547 3349 25556 3383
rect 25504 3340 25556 3349
rect 25872 3340 25924 3392
rect 26792 3340 26844 3392
rect 28080 3340 28132 3392
rect 29000 3383 29052 3392
rect 29000 3349 29009 3383
rect 29009 3349 29043 3383
rect 29043 3349 29052 3383
rect 29000 3340 29052 3349
rect 31392 3408 31444 3460
rect 36268 3408 36320 3460
rect 30288 3340 30340 3392
rect 34428 3340 34480 3392
rect 36176 3340 36228 3392
rect 38660 3340 38712 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 2504 3136 2556 3188
rect 4620 3136 4672 3188
rect 7840 3179 7892 3188
rect 7840 3145 7849 3179
rect 7849 3145 7883 3179
rect 7883 3145 7892 3179
rect 7840 3136 7892 3145
rect 8944 3136 8996 3188
rect 11152 3136 11204 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 18696 3179 18748 3188
rect 18696 3145 18705 3179
rect 18705 3145 18739 3179
rect 18739 3145 18748 3179
rect 18696 3136 18748 3145
rect 20996 3179 21048 3188
rect 20996 3145 21005 3179
rect 21005 3145 21039 3179
rect 21039 3145 21048 3179
rect 20996 3136 21048 3145
rect 24492 3136 24544 3188
rect 664 3068 716 3120
rect 4252 3068 4304 3120
rect 5172 3068 5224 3120
rect 16948 3068 17000 3120
rect 20628 3068 20680 3120
rect 22100 3068 22152 3120
rect 23848 3068 23900 3120
rect 26148 3136 26200 3188
rect 27896 3136 27948 3188
rect 29368 3136 29420 3188
rect 29920 3136 29972 3188
rect 30564 3136 30616 3188
rect 25228 3068 25280 3120
rect 26792 3111 26844 3120
rect 26792 3077 26801 3111
rect 26801 3077 26835 3111
rect 26835 3077 26844 3111
rect 26792 3068 26844 3077
rect 27160 3068 27212 3120
rect 31668 3136 31720 3188
rect 32404 3179 32456 3188
rect 32404 3145 32413 3179
rect 32413 3145 32447 3179
rect 32447 3145 32456 3179
rect 32404 3136 32456 3145
rect 33140 3179 33192 3188
rect 33140 3145 33149 3179
rect 33149 3145 33183 3179
rect 33183 3145 33192 3179
rect 33140 3136 33192 3145
rect 33876 3179 33928 3188
rect 33876 3145 33885 3179
rect 33885 3145 33919 3179
rect 33919 3145 33928 3179
rect 33876 3136 33928 3145
rect 37832 3136 37884 3188
rect 38016 3179 38068 3188
rect 38016 3145 38025 3179
rect 38025 3145 38059 3179
rect 38059 3145 38068 3179
rect 38016 3136 38068 3145
rect 35624 3068 35676 3120
rect 112 3000 164 3052
rect 1216 3000 1268 3052
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 13728 3000 13780 3052
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 19524 3000 19576 3052
rect 22376 3000 22428 3052
rect 2964 2932 3016 2984
rect 4160 2932 4212 2984
rect 5080 2975 5132 2984
rect 5080 2941 5089 2975
rect 5089 2941 5123 2975
rect 5123 2941 5132 2975
rect 5080 2932 5132 2941
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 6460 2975 6512 2984
rect 6460 2941 6469 2975
rect 6469 2941 6503 2975
rect 6503 2941 6512 2975
rect 6460 2932 6512 2941
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 8208 2932 8260 2984
rect 9404 2932 9456 2984
rect 10876 2975 10928 2984
rect 10876 2941 10885 2975
rect 10885 2941 10919 2975
rect 10919 2941 10928 2975
rect 10876 2932 10928 2941
rect 11796 2975 11848 2984
rect 11796 2941 11805 2975
rect 11805 2941 11839 2975
rect 11839 2941 11848 2975
rect 11796 2932 11848 2941
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 14740 2932 14792 2984
rect 15568 2975 15620 2984
rect 2780 2864 2832 2916
rect 7932 2864 7984 2916
rect 9588 2907 9640 2916
rect 4620 2796 4672 2848
rect 5632 2796 5684 2848
rect 9588 2873 9597 2907
rect 9597 2873 9631 2907
rect 9631 2873 9640 2907
rect 9588 2864 9640 2873
rect 14556 2864 14608 2916
rect 14832 2907 14884 2916
rect 14832 2873 14841 2907
rect 14841 2873 14875 2907
rect 14875 2873 14884 2907
rect 14832 2864 14884 2873
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 17040 2932 17092 2984
rect 17960 2932 18012 2984
rect 18144 2932 18196 2984
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 20812 2975 20864 2984
rect 20812 2941 20821 2975
rect 20821 2941 20855 2975
rect 20855 2941 20864 2975
rect 20812 2932 20864 2941
rect 21824 2932 21876 2984
rect 20260 2864 20312 2916
rect 22100 2864 22152 2916
rect 22376 2907 22428 2916
rect 22376 2873 22385 2907
rect 22385 2873 22419 2907
rect 22419 2873 22428 2907
rect 22376 2864 22428 2873
rect 22560 3000 22612 3052
rect 26516 3043 26568 3052
rect 23940 2932 23992 2984
rect 25320 2975 25372 2984
rect 25320 2941 25329 2975
rect 25329 2941 25363 2975
rect 25363 2941 25372 2975
rect 25320 2932 25372 2941
rect 26240 2932 26292 2984
rect 26516 3009 26525 3043
rect 26525 3009 26559 3043
rect 26559 3009 26568 3043
rect 26516 3000 26568 3009
rect 31484 3000 31536 3052
rect 35992 3043 36044 3052
rect 27528 2932 27580 2984
rect 28172 2975 28224 2984
rect 28172 2941 28181 2975
rect 28181 2941 28215 2975
rect 28215 2941 28224 2975
rect 28172 2932 28224 2941
rect 29552 2932 29604 2984
rect 32220 2975 32272 2984
rect 26332 2864 26384 2916
rect 13176 2796 13228 2848
rect 17776 2796 17828 2848
rect 19340 2796 19392 2848
rect 21088 2796 21140 2848
rect 22008 2796 22060 2848
rect 22928 2796 22980 2848
rect 24584 2796 24636 2848
rect 25596 2796 25648 2848
rect 30472 2864 30524 2916
rect 31116 2864 31168 2916
rect 32220 2941 32229 2975
rect 32229 2941 32263 2975
rect 32263 2941 32272 2975
rect 32220 2932 32272 2941
rect 32496 2932 32548 2984
rect 33048 2932 33100 2984
rect 34428 2975 34480 2984
rect 34428 2941 34437 2975
rect 34437 2941 34471 2975
rect 34471 2941 34480 2975
rect 34428 2932 34480 2941
rect 35256 2932 35308 2984
rect 35992 3009 36001 3043
rect 36001 3009 36035 3043
rect 36035 3009 36044 3043
rect 35992 3000 36044 3009
rect 37280 3000 37332 3052
rect 38016 3000 38068 3052
rect 37740 2932 37792 2984
rect 35348 2864 35400 2916
rect 36728 2864 36780 2916
rect 37924 2907 37976 2916
rect 37924 2873 37933 2907
rect 37933 2873 37967 2907
rect 37967 2873 37976 2907
rect 37924 2864 37976 2873
rect 28264 2839 28316 2848
rect 28264 2805 28273 2839
rect 28273 2805 28307 2839
rect 28307 2805 28316 2839
rect 28264 2796 28316 2805
rect 28448 2796 28500 2848
rect 37832 2796 37884 2848
rect 39764 2796 39816 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 4252 2592 4304 2644
rect 5540 2592 5592 2644
rect 2872 2524 2924 2576
rect 4712 2524 4764 2576
rect 5264 2567 5316 2576
rect 5264 2533 5273 2567
rect 5273 2533 5307 2567
rect 5307 2533 5316 2567
rect 5264 2524 5316 2533
rect 7196 2567 7248 2576
rect 7196 2533 7205 2567
rect 7205 2533 7239 2567
rect 7239 2533 7248 2567
rect 7196 2524 7248 2533
rect 388 2456 440 2508
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3884 2456 3936 2508
rect 6184 2456 6236 2508
rect 8668 2592 8720 2644
rect 20996 2592 21048 2644
rect 22100 2592 22152 2644
rect 29828 2592 29880 2644
rect 32128 2635 32180 2644
rect 32128 2601 32137 2635
rect 32137 2601 32171 2635
rect 32171 2601 32180 2635
rect 32128 2592 32180 2601
rect 33784 2635 33836 2644
rect 33784 2601 33793 2635
rect 33793 2601 33827 2635
rect 33827 2601 33836 2635
rect 33784 2592 33836 2601
rect 35532 2592 35584 2644
rect 10140 2524 10192 2576
rect 12440 2524 12492 2576
rect 13912 2524 13964 2576
rect 15292 2524 15344 2576
rect 17132 2524 17184 2576
rect 17408 2524 17460 2576
rect 19064 2524 19116 2576
rect 23664 2524 23716 2576
rect 25688 2524 25740 2576
rect 32680 2524 32732 2576
rect 34704 2524 34756 2576
rect 9128 2456 9180 2508
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 10324 2456 10376 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 14372 2456 14424 2508
rect 17316 2456 17368 2508
rect 19892 2456 19944 2508
rect 21640 2456 21692 2508
rect 23480 2499 23532 2508
rect 23480 2465 23489 2499
rect 23489 2465 23523 2499
rect 23523 2465 23532 2499
rect 23480 2456 23532 2465
rect 24308 2456 24360 2508
rect 26976 2499 27028 2508
rect 26976 2465 26985 2499
rect 26985 2465 27019 2499
rect 27019 2465 27028 2499
rect 26976 2456 27028 2465
rect 27804 2456 27856 2508
rect 28724 2456 28776 2508
rect 30472 2456 30524 2508
rect 31944 2499 31996 2508
rect 31944 2465 31953 2499
rect 31953 2465 31987 2499
rect 31987 2465 31996 2499
rect 31944 2456 31996 2465
rect 32772 2456 32824 2508
rect 34796 2499 34848 2508
rect 34796 2465 34805 2499
rect 34805 2465 34839 2499
rect 34839 2465 34848 2499
rect 34796 2456 34848 2465
rect 36544 2499 36596 2508
rect 36544 2465 36553 2499
rect 36553 2465 36587 2499
rect 36587 2465 36596 2499
rect 36544 2456 36596 2465
rect 38292 2456 38344 2508
rect 15292 2388 15344 2440
rect 19064 2388 19116 2440
rect 19156 2388 19208 2440
rect 28540 2388 28592 2440
rect 29644 2388 29696 2440
rect 32588 2388 32640 2440
rect 7840 2320 7892 2372
rect 21272 2320 21324 2372
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 27252 1436 27304 1488
rect 28264 1436 28316 1488
<< metal2 >>
rect 110 119200 166 120800
rect 294 119200 350 120800
rect 478 119200 534 120800
rect 662 119200 718 120800
rect 938 119200 994 120800
rect 1122 119200 1178 120800
rect 1306 119200 1362 120800
rect 1582 119200 1638 120800
rect 1766 119200 1822 120800
rect 1950 119200 2006 120800
rect 2226 119200 2282 120800
rect 2410 119200 2466 120800
rect 2594 119200 2650 120800
rect 2778 119200 2834 120800
rect 3054 119200 3110 120800
rect 3238 119200 3294 120800
rect 3330 119504 3386 119513
rect 3330 119439 3386 119448
rect 124 117298 152 119200
rect 308 117434 336 119200
rect 296 117428 348 117434
rect 296 117370 348 117376
rect 112 117292 164 117298
rect 112 117234 164 117240
rect 492 115734 520 119200
rect 676 117230 704 119200
rect 664 117224 716 117230
rect 664 117166 716 117172
rect 952 117094 980 119200
rect 1136 117366 1164 119200
rect 1124 117360 1176 117366
rect 1124 117302 1176 117308
rect 940 117088 992 117094
rect 940 117030 992 117036
rect 1320 116890 1348 119200
rect 1308 116884 1360 116890
rect 1308 116826 1360 116832
rect 1398 116240 1454 116249
rect 1398 116175 1454 116184
rect 480 115728 532 115734
rect 480 115670 532 115676
rect 1412 115258 1440 116175
rect 1596 115598 1624 119200
rect 1676 115796 1728 115802
rect 1676 115738 1728 115744
rect 1584 115592 1636 115598
rect 1584 115534 1636 115540
rect 1400 115252 1452 115258
rect 1400 115194 1452 115200
rect 1688 112946 1716 115738
rect 1780 113490 1808 119200
rect 1860 117156 1912 117162
rect 1860 117098 1912 117104
rect 1872 116278 1900 117098
rect 1964 116906 1992 119200
rect 1964 116878 2176 116906
rect 2148 116822 2176 116878
rect 2136 116816 2188 116822
rect 2136 116758 2188 116764
rect 2240 116346 2268 119200
rect 2228 116340 2280 116346
rect 2228 116282 2280 116288
rect 1860 116272 1912 116278
rect 1860 116214 1912 116220
rect 2320 116068 2372 116074
rect 2320 116010 2372 116016
rect 1952 115456 2004 115462
rect 1950 115424 1952 115433
rect 2004 115424 2006 115433
rect 1950 115359 2006 115368
rect 1860 114980 1912 114986
rect 1860 114922 1912 114928
rect 1768 113484 1820 113490
rect 1768 113426 1820 113432
rect 1872 113174 1900 114922
rect 2042 114608 2098 114617
rect 2042 114543 2098 114552
rect 2056 114510 2084 114543
rect 2044 114504 2096 114510
rect 2044 114446 2096 114452
rect 2136 113892 2188 113898
rect 2136 113834 2188 113840
rect 1952 113824 2004 113830
rect 1950 113792 1952 113801
rect 2004 113792 2006 113801
rect 1950 113727 2006 113736
rect 1780 113146 1900 113174
rect 1676 112940 1728 112946
rect 1676 112882 1728 112888
rect 1398 111344 1454 111353
rect 1398 111279 1400 111288
rect 1452 111279 1454 111288
rect 1400 111250 1452 111256
rect 1780 107794 1808 113146
rect 1858 112976 1914 112985
rect 1858 112911 1914 112920
rect 1872 112878 1900 112911
rect 1860 112872 1912 112878
rect 1860 112814 1912 112820
rect 1952 112192 2004 112198
rect 1950 112160 1952 112169
rect 2004 112160 2006 112169
rect 1950 112095 2006 112104
rect 1952 110560 2004 110566
rect 1950 110528 1952 110537
rect 2004 110528 2006 110537
rect 1950 110463 2006 110472
rect 2044 109608 2096 109614
rect 2042 109576 2044 109585
rect 2096 109576 2098 109585
rect 2042 109511 2098 109520
rect 1950 108760 2006 108769
rect 1950 108695 1952 108704
rect 2004 108695 2006 108704
rect 1952 108666 2004 108672
rect 2042 107944 2098 107953
rect 2042 107879 2044 107888
rect 2096 107879 2098 107888
rect 2044 107850 2096 107856
rect 1780 107766 2084 107794
rect 1950 107128 2006 107137
rect 1950 107063 1952 107072
rect 2004 107063 2006 107072
rect 1952 107034 2004 107040
rect 1768 106344 1820 106350
rect 1766 106312 1768 106321
rect 1820 106312 1822 106321
rect 1766 106247 1822 106256
rect 1398 105496 1454 105505
rect 1398 105431 1454 105440
rect 1412 105262 1440 105431
rect 1400 105256 1452 105262
rect 1400 105198 1452 105204
rect 1860 104780 1912 104786
rect 1860 104722 1912 104728
rect 1872 104689 1900 104722
rect 1858 104680 1914 104689
rect 1858 104615 1914 104624
rect 1858 103864 1914 103873
rect 1858 103799 1914 103808
rect 1872 103766 1900 103799
rect 1860 103760 1912 103766
rect 1860 103702 1912 103708
rect 2056 103222 2084 107766
rect 2044 103216 2096 103222
rect 2044 103158 2096 103164
rect 1858 103048 1914 103057
rect 1858 102983 1860 102992
rect 1912 102983 1914 102992
rect 1860 102954 1912 102960
rect 1858 102232 1914 102241
rect 1858 102167 1914 102176
rect 1872 101998 1900 102167
rect 1860 101992 1912 101998
rect 1860 101934 1912 101940
rect 2044 101924 2096 101930
rect 2044 101866 2096 101872
rect 1860 101516 1912 101522
rect 1860 101458 1912 101464
rect 1872 101425 1900 101458
rect 1858 101416 1914 101425
rect 1858 101351 1914 101360
rect 1858 100600 1914 100609
rect 1858 100535 1914 100544
rect 1872 100502 1900 100535
rect 1860 100496 1912 100502
rect 1860 100438 1912 100444
rect 1860 99748 1912 99754
rect 1860 99690 1912 99696
rect 1872 99657 1900 99690
rect 1858 99648 1914 99657
rect 1858 99583 1914 99592
rect 1858 98832 1914 98841
rect 1858 98767 1914 98776
rect 1872 98734 1900 98767
rect 1860 98728 1912 98734
rect 1860 98670 1912 98676
rect 1860 98252 1912 98258
rect 1860 98194 1912 98200
rect 1872 98025 1900 98194
rect 1858 98016 1914 98025
rect 1858 97951 1914 97960
rect 1858 97200 1914 97209
rect 1858 97135 1860 97144
rect 1912 97135 1914 97144
rect 1860 97106 1912 97112
rect 1860 96484 1912 96490
rect 1860 96426 1912 96432
rect 1872 96393 1900 96426
rect 1858 96384 1914 96393
rect 1858 96319 1914 96328
rect 1952 95872 2004 95878
rect 1952 95814 2004 95820
rect 1964 95674 1992 95814
rect 1952 95668 2004 95674
rect 1952 95610 2004 95616
rect 1858 95568 1914 95577
rect 1858 95503 1914 95512
rect 1872 95470 1900 95503
rect 1860 95464 1912 95470
rect 1860 95406 1912 95412
rect 1860 94988 1912 94994
rect 1860 94930 1912 94936
rect 1872 94761 1900 94930
rect 1858 94752 1914 94761
rect 1858 94687 1914 94696
rect 1858 93936 1914 93945
rect 1858 93871 1860 93880
rect 1912 93871 1914 93880
rect 1860 93842 1912 93848
rect 2056 93294 2084 101866
rect 2148 101658 2176 113834
rect 2332 113490 2360 116010
rect 2424 115802 2452 119200
rect 2608 116890 2636 119200
rect 2596 116884 2648 116890
rect 2596 116826 2648 116832
rect 2596 116748 2648 116754
rect 2596 116690 2648 116696
rect 2412 115796 2464 115802
rect 2412 115738 2464 115744
rect 2504 115660 2556 115666
rect 2504 115602 2556 115608
rect 2412 114572 2464 114578
rect 2412 114514 2464 114520
rect 2320 113484 2372 113490
rect 2320 113426 2372 113432
rect 2228 110628 2280 110634
rect 2228 110570 2280 110576
rect 2136 101652 2188 101658
rect 2136 101594 2188 101600
rect 2240 98394 2268 110570
rect 2424 101454 2452 114514
rect 2516 109070 2544 115602
rect 2608 114170 2636 116690
rect 2792 116346 2820 119200
rect 2962 117872 3018 117881
rect 2962 117807 3018 117816
rect 2870 117056 2926 117065
rect 2870 116991 2926 117000
rect 2780 116340 2832 116346
rect 2780 116282 2832 116288
rect 2884 115190 2912 116991
rect 2976 115734 3004 117807
rect 3068 116362 3096 119200
rect 3146 118688 3202 118697
rect 3146 118623 3202 118632
rect 3160 116498 3188 118623
rect 3252 116822 3280 119200
rect 3240 116816 3292 116822
rect 3240 116758 3292 116764
rect 3160 116470 3280 116498
rect 3068 116334 3188 116362
rect 3056 116068 3108 116074
rect 3056 116010 3108 116016
rect 2964 115728 3016 115734
rect 2964 115670 3016 115676
rect 2872 115184 2924 115190
rect 2872 115126 2924 115132
rect 2688 115048 2740 115054
rect 2688 114990 2740 114996
rect 2596 114164 2648 114170
rect 2596 114106 2648 114112
rect 2504 109064 2556 109070
rect 2504 109006 2556 109012
rect 2700 102746 2728 114990
rect 3068 113490 3096 116010
rect 3160 113490 3188 116334
rect 3252 114510 3280 116470
rect 3240 114504 3292 114510
rect 3240 114446 3292 114452
rect 3344 114374 3372 119439
rect 3422 119200 3478 120800
rect 3698 119200 3754 120800
rect 3882 119200 3938 120800
rect 4066 119200 4122 120800
rect 4342 119200 4398 120800
rect 4526 119200 4582 120800
rect 4710 119200 4766 120800
rect 4894 119200 4950 120800
rect 5170 119200 5226 120800
rect 5354 119200 5410 120800
rect 5538 119200 5594 120800
rect 5814 119200 5870 120800
rect 5998 119200 6054 120800
rect 6182 119200 6238 120800
rect 6458 119200 6514 120800
rect 6642 119200 6698 120800
rect 6826 119200 6882 120800
rect 7010 119200 7066 120800
rect 7286 119200 7342 120800
rect 7470 119200 7526 120800
rect 7654 119200 7710 120800
rect 7930 119200 7986 120800
rect 8114 119200 8170 120800
rect 8298 119200 8354 120800
rect 8574 119200 8630 120800
rect 8758 119200 8814 120800
rect 8942 119200 8998 120800
rect 9126 119200 9182 120800
rect 9402 119200 9458 120800
rect 9586 119200 9642 120800
rect 9770 119200 9826 120800
rect 10046 119200 10102 120800
rect 10230 119200 10286 120800
rect 10414 119200 10470 120800
rect 10690 119200 10746 120800
rect 10874 119200 10930 120800
rect 11058 119200 11114 120800
rect 11242 119200 11298 120800
rect 11518 119200 11574 120800
rect 11702 119200 11758 120800
rect 11886 119200 11942 120800
rect 12162 119200 12218 120800
rect 12346 119200 12402 120800
rect 12530 119200 12586 120800
rect 12806 119200 12862 120800
rect 12990 119200 13046 120800
rect 13174 119200 13230 120800
rect 13450 119200 13506 120800
rect 13634 119200 13690 120800
rect 13818 119200 13874 120800
rect 14002 119200 14058 120800
rect 14278 119200 14334 120800
rect 14462 119200 14518 120800
rect 14646 119200 14702 120800
rect 14922 119200 14978 120800
rect 15106 119200 15162 120800
rect 15290 119200 15346 120800
rect 15566 119200 15622 120800
rect 15750 119200 15806 120800
rect 15934 119200 15990 120800
rect 16118 119200 16174 120800
rect 16394 119200 16450 120800
rect 16578 119200 16634 120800
rect 16762 119200 16818 120800
rect 17038 119200 17094 120800
rect 17222 119200 17278 120800
rect 17406 119200 17462 120800
rect 17682 119200 17738 120800
rect 17866 119200 17922 120800
rect 18050 119200 18106 120800
rect 18234 119200 18290 120800
rect 18510 119200 18566 120800
rect 18694 119200 18750 120800
rect 18878 119200 18934 120800
rect 19154 119200 19210 120800
rect 19338 119200 19394 120800
rect 19522 119200 19578 120800
rect 19798 119200 19854 120800
rect 19982 119200 20038 120800
rect 20166 119200 20222 120800
rect 20350 119200 20406 120800
rect 20626 119200 20682 120800
rect 20810 119200 20866 120800
rect 20994 119200 21050 120800
rect 21270 119200 21326 120800
rect 21454 119200 21510 120800
rect 21638 119200 21694 120800
rect 21914 119200 21970 120800
rect 22098 119200 22154 120800
rect 22282 119200 22338 120800
rect 22466 119200 22522 120800
rect 22742 119200 22798 120800
rect 22926 119200 22982 120800
rect 23110 119200 23166 120800
rect 23386 119200 23442 120800
rect 23570 119200 23626 120800
rect 23754 119200 23810 120800
rect 24030 119200 24086 120800
rect 24214 119200 24270 120800
rect 24398 119200 24454 120800
rect 24582 119200 24638 120800
rect 24858 119200 24914 120800
rect 25042 119200 25098 120800
rect 25226 119200 25282 120800
rect 25502 119200 25558 120800
rect 25686 119200 25742 120800
rect 25870 119200 25926 120800
rect 26146 119200 26202 120800
rect 26330 119200 26386 120800
rect 26514 119200 26570 120800
rect 26790 119200 26846 120800
rect 26974 119200 27030 120800
rect 27158 119200 27214 120800
rect 27342 119200 27398 120800
rect 27618 119200 27674 120800
rect 27802 119200 27858 120800
rect 27986 119200 28042 120800
rect 28262 119200 28318 120800
rect 28446 119200 28502 120800
rect 28630 119200 28686 120800
rect 28906 119200 28962 120800
rect 29090 119200 29146 120800
rect 29274 119200 29330 120800
rect 29458 119200 29514 120800
rect 29734 119200 29790 120800
rect 29918 119200 29974 120800
rect 30102 119200 30158 120800
rect 30378 119200 30434 120800
rect 30562 119200 30618 120800
rect 30746 119200 30802 120800
rect 31022 119200 31078 120800
rect 31206 119200 31262 120800
rect 31390 119200 31446 120800
rect 31574 119200 31630 120800
rect 31850 119200 31906 120800
rect 32034 119200 32090 120800
rect 32218 119200 32274 120800
rect 32494 119200 32550 120800
rect 32678 119200 32734 120800
rect 32862 119200 32918 120800
rect 33138 119200 33194 120800
rect 33322 119200 33378 120800
rect 33506 119200 33562 120800
rect 33690 119200 33746 120800
rect 33966 119200 34022 120800
rect 34150 119200 34206 120800
rect 34334 119200 34390 120800
rect 34610 119200 34666 120800
rect 34794 119200 34850 120800
rect 34978 119200 35034 120800
rect 35254 119200 35310 120800
rect 35438 119200 35494 120800
rect 35622 119200 35678 120800
rect 35806 119200 35862 120800
rect 36082 119200 36138 120800
rect 36266 119200 36322 120800
rect 36358 119640 36414 119649
rect 36358 119575 36414 119584
rect 3436 116634 3464 119200
rect 3608 117156 3660 117162
rect 3608 117098 3660 117104
rect 3436 116606 3556 116634
rect 3424 116544 3476 116550
rect 3424 116486 3476 116492
rect 3436 115802 3464 116486
rect 3528 115802 3556 116606
rect 3620 116210 3648 117098
rect 3608 116204 3660 116210
rect 3608 116146 3660 116152
rect 3424 115796 3476 115802
rect 3424 115738 3476 115744
rect 3516 115796 3568 115802
rect 3516 115738 3568 115744
rect 3608 115660 3660 115666
rect 3608 115602 3660 115608
rect 3516 114640 3568 114646
rect 3516 114582 3568 114588
rect 3332 114368 3384 114374
rect 3332 114310 3384 114316
rect 3056 113484 3108 113490
rect 3056 113426 3108 113432
rect 3148 113484 3200 113490
rect 3148 113426 3200 113432
rect 3424 109064 3476 109070
rect 3424 109006 3476 109012
rect 2688 102740 2740 102746
rect 2688 102682 2740 102688
rect 2412 101448 2464 101454
rect 2412 101390 2464 101396
rect 3436 99142 3464 109006
rect 3528 103290 3556 114582
rect 3620 114102 3648 115602
rect 3712 114730 3740 119200
rect 3792 116748 3844 116754
rect 3792 116690 3844 116696
rect 3804 114866 3832 116690
rect 3896 116686 3924 119200
rect 4080 116906 4108 119200
rect 4356 117706 4384 119200
rect 4540 117722 4568 119200
rect 4344 117700 4396 117706
rect 4540 117694 4660 117722
rect 4344 117642 4396 117648
rect 4220 117532 4516 117552
rect 4276 117530 4300 117532
rect 4356 117530 4380 117532
rect 4436 117530 4460 117532
rect 4298 117478 4300 117530
rect 4362 117478 4374 117530
rect 4436 117478 4438 117530
rect 4276 117476 4300 117478
rect 4356 117476 4380 117478
rect 4436 117476 4460 117478
rect 4220 117456 4516 117476
rect 3988 116878 4108 116906
rect 3884 116680 3936 116686
rect 3884 116622 3936 116628
rect 3988 115734 4016 116878
rect 4068 116748 4120 116754
rect 4068 116690 4120 116696
rect 3976 115728 4028 115734
rect 3976 115670 4028 115676
rect 4080 115258 4108 116690
rect 4220 116444 4516 116464
rect 4276 116442 4300 116444
rect 4356 116442 4380 116444
rect 4436 116442 4460 116444
rect 4298 116390 4300 116442
rect 4362 116390 4374 116442
rect 4436 116390 4438 116442
rect 4276 116388 4300 116390
rect 4356 116388 4380 116390
rect 4436 116388 4460 116390
rect 4220 116368 4516 116388
rect 4632 116346 4660 117694
rect 4620 116340 4672 116346
rect 4620 116282 4672 116288
rect 4528 116204 4580 116210
rect 4528 116146 4580 116152
rect 4540 115530 4568 116146
rect 4724 115802 4752 119200
rect 4908 117858 4936 119200
rect 4908 117830 5028 117858
rect 4896 117700 4948 117706
rect 4896 117642 4948 117648
rect 4804 116748 4856 116754
rect 4804 116690 4856 116696
rect 4712 115796 4764 115802
rect 4712 115738 4764 115744
rect 4620 115660 4672 115666
rect 4620 115602 4672 115608
rect 4528 115524 4580 115530
rect 4528 115466 4580 115472
rect 4220 115356 4516 115376
rect 4276 115354 4300 115356
rect 4356 115354 4380 115356
rect 4436 115354 4460 115356
rect 4298 115302 4300 115354
rect 4362 115302 4374 115354
rect 4436 115302 4438 115354
rect 4276 115300 4300 115302
rect 4356 115300 4380 115302
rect 4436 115300 4460 115302
rect 4220 115280 4516 115300
rect 4068 115252 4120 115258
rect 4068 115194 4120 115200
rect 3804 114838 3924 114866
rect 3712 114702 3832 114730
rect 3700 114572 3752 114578
rect 3700 114514 3752 114520
rect 3608 114096 3660 114102
rect 3608 114038 3660 114044
rect 3516 103284 3568 103290
rect 3516 103226 3568 103232
rect 3424 99136 3476 99142
rect 3424 99078 3476 99084
rect 3516 98660 3568 98666
rect 3516 98602 3568 98608
rect 2228 98388 2280 98394
rect 2228 98330 2280 98336
rect 2044 93288 2096 93294
rect 2044 93230 2096 93236
rect 1860 93220 1912 93226
rect 1860 93162 1912 93168
rect 1872 93129 1900 93162
rect 1858 93120 1914 93129
rect 1858 93055 1914 93064
rect 1858 92304 1914 92313
rect 1858 92239 1914 92248
rect 1872 92206 1900 92239
rect 1860 92200 1912 92206
rect 1860 92142 1912 92148
rect 1860 91724 1912 91730
rect 1860 91666 1912 91672
rect 1872 91497 1900 91666
rect 1952 91520 2004 91526
rect 1858 91488 1914 91497
rect 1952 91462 2004 91468
rect 1858 91423 1914 91432
rect 1964 91322 1992 91462
rect 1952 91316 2004 91322
rect 1952 91258 2004 91264
rect 1858 90672 1914 90681
rect 1858 90607 1860 90616
rect 1912 90607 1914 90616
rect 1860 90578 1912 90584
rect 1952 90432 2004 90438
rect 1952 90374 2004 90380
rect 1964 90234 1992 90374
rect 1952 90228 2004 90234
rect 1952 90170 2004 90176
rect 1858 89720 1914 89729
rect 1858 89655 1914 89664
rect 1872 89622 1900 89655
rect 1860 89616 1912 89622
rect 1860 89558 1912 89564
rect 3424 89412 3476 89418
rect 3424 89354 3476 89360
rect 1858 88904 1914 88913
rect 1858 88839 1860 88848
rect 1912 88839 1914 88848
rect 1860 88810 1912 88816
rect 1858 88088 1914 88097
rect 1858 88023 1914 88032
rect 1872 87854 1900 88023
rect 1860 87848 1912 87854
rect 1860 87790 1912 87796
rect 1860 87372 1912 87378
rect 1860 87314 1912 87320
rect 1872 87281 1900 87314
rect 1858 87272 1914 87281
rect 1858 87207 1914 87216
rect 1952 87168 2004 87174
rect 1952 87110 2004 87116
rect 1858 86456 1914 86465
rect 1858 86391 1914 86400
rect 1872 86358 1900 86391
rect 1860 86352 1912 86358
rect 1860 86294 1912 86300
rect 1860 85672 1912 85678
rect 1858 85640 1860 85649
rect 1912 85640 1914 85649
rect 1858 85575 1914 85584
rect 1858 84824 1914 84833
rect 1858 84759 1914 84768
rect 1872 84590 1900 84759
rect 1860 84584 1912 84590
rect 1860 84526 1912 84532
rect 1860 84108 1912 84114
rect 1860 84050 1912 84056
rect 1872 84017 1900 84050
rect 1858 84008 1914 84017
rect 1858 83943 1914 83952
rect 1398 83192 1454 83201
rect 1398 83127 1454 83136
rect 1412 83026 1440 83127
rect 1400 83020 1452 83026
rect 1400 82962 1452 82968
rect 1964 82482 1992 87110
rect 2044 86148 2096 86154
rect 2044 86090 2096 86096
rect 2056 82550 2084 86090
rect 2688 85604 2740 85610
rect 2688 85546 2740 85552
rect 2596 84516 2648 84522
rect 2596 84458 2648 84464
rect 2044 82544 2096 82550
rect 2044 82486 2096 82492
rect 1952 82476 2004 82482
rect 1952 82418 2004 82424
rect 1858 82376 1914 82385
rect 1858 82311 1860 82320
rect 1912 82311 1914 82320
rect 1860 82282 1912 82288
rect 1858 81560 1914 81569
rect 1858 81495 1914 81504
rect 1872 81326 1900 81495
rect 1860 81320 1912 81326
rect 1860 81262 1912 81268
rect 2044 81252 2096 81258
rect 2044 81194 2096 81200
rect 1400 80844 1452 80850
rect 1400 80786 1452 80792
rect 1412 80753 1440 80786
rect 1398 80744 1454 80753
rect 1398 80679 1454 80688
rect 1398 79792 1454 79801
rect 1398 79727 1400 79736
rect 1452 79727 1454 79736
rect 1400 79698 1452 79704
rect 2056 79694 2084 81194
rect 2608 80238 2636 84458
rect 2700 80918 2728 85546
rect 3436 83638 3464 89354
rect 3528 88942 3556 98602
rect 3516 88936 3568 88942
rect 3516 88878 3568 88884
rect 3516 87780 3568 87786
rect 3516 87722 3568 87728
rect 3424 83632 3476 83638
rect 3424 83574 3476 83580
rect 3528 83094 3556 87722
rect 3516 83088 3568 83094
rect 3516 83030 3568 83036
rect 2688 80912 2740 80918
rect 2688 80854 2740 80860
rect 2688 80640 2740 80646
rect 2688 80582 2740 80588
rect 2596 80232 2648 80238
rect 2596 80174 2648 80180
rect 2044 79688 2096 79694
rect 2044 79630 2096 79636
rect 1584 79552 1636 79558
rect 1584 79494 1636 79500
rect 1596 78538 1624 79494
rect 2700 79218 2728 80582
rect 2688 79212 2740 79218
rect 2688 79154 2740 79160
rect 1860 79076 1912 79082
rect 1860 79018 1912 79024
rect 2044 79076 2096 79082
rect 2044 79018 2096 79024
rect 1872 78985 1900 79018
rect 1858 78976 1914 78985
rect 1858 78911 1914 78920
rect 1584 78532 1636 78538
rect 1584 78474 1636 78480
rect 1858 78160 1914 78169
rect 1858 78095 1914 78104
rect 1872 78062 1900 78095
rect 1860 78056 1912 78062
rect 1860 77998 1912 78004
rect 1952 77920 2004 77926
rect 1952 77862 2004 77868
rect 1400 77580 1452 77586
rect 1400 77522 1452 77528
rect 1412 77353 1440 77522
rect 1398 77344 1454 77353
rect 1398 77279 1454 77288
rect 1398 76528 1454 76537
rect 1398 76463 1400 76472
rect 1452 76463 1454 76472
rect 1400 76434 1452 76440
rect 1860 75812 1912 75818
rect 1860 75754 1912 75760
rect 1872 75721 1900 75754
rect 1858 75712 1914 75721
rect 1858 75647 1914 75656
rect 1858 74896 1914 74905
rect 1858 74831 1914 74840
rect 1872 74798 1900 74831
rect 1860 74792 1912 74798
rect 1860 74734 1912 74740
rect 1860 74316 1912 74322
rect 1860 74258 1912 74264
rect 1872 74089 1900 74258
rect 1858 74080 1914 74089
rect 1858 74015 1914 74024
rect 1858 73264 1914 73273
rect 1858 73199 1860 73208
rect 1912 73199 1914 73208
rect 1860 73170 1912 73176
rect 1860 72548 1912 72554
rect 1860 72490 1912 72496
rect 1872 72457 1900 72490
rect 1858 72448 1914 72457
rect 1858 72383 1914 72392
rect 1858 71632 1914 71641
rect 1858 71567 1914 71576
rect 1872 71534 1900 71567
rect 1860 71528 1912 71534
rect 1860 71470 1912 71476
rect 1860 71052 1912 71058
rect 1860 70994 1912 71000
rect 1872 70825 1900 70994
rect 1858 70816 1914 70825
rect 1858 70751 1914 70760
rect 1860 69964 1912 69970
rect 1860 69906 1912 69912
rect 1872 69873 1900 69906
rect 1858 69864 1914 69873
rect 1858 69799 1914 69808
rect 1858 69048 1914 69057
rect 1858 68983 1914 68992
rect 1872 68950 1900 68983
rect 1860 68944 1912 68950
rect 1860 68886 1912 68892
rect 1860 68264 1912 68270
rect 1858 68232 1860 68241
rect 1912 68232 1914 68241
rect 1858 68167 1914 68176
rect 1398 67416 1454 67425
rect 1398 67351 1454 67360
rect 1412 67182 1440 67351
rect 1400 67176 1452 67182
rect 1400 67118 1452 67124
rect 1400 66700 1452 66706
rect 1400 66642 1452 66648
rect 1412 66609 1440 66642
rect 1398 66600 1454 66609
rect 1398 66535 1454 66544
rect 1398 65784 1454 65793
rect 1398 65719 1454 65728
rect 1412 65618 1440 65719
rect 1400 65612 1452 65618
rect 1400 65554 1452 65560
rect 1964 65550 1992 77862
rect 1952 65544 2004 65550
rect 1952 65486 2004 65492
rect 1676 65408 1728 65414
rect 1676 65350 1728 65356
rect 1400 65000 1452 65006
rect 1398 64968 1400 64977
rect 1452 64968 1454 64977
rect 1398 64903 1454 64912
rect 1398 64152 1454 64161
rect 1398 64087 1454 64096
rect 1412 63918 1440 64087
rect 1400 63912 1452 63918
rect 1400 63854 1452 63860
rect 1400 63436 1452 63442
rect 1400 63378 1452 63384
rect 1412 63345 1440 63378
rect 1398 63336 1454 63345
rect 1398 63271 1454 63280
rect 1398 62520 1454 62529
rect 1398 62455 1454 62464
rect 1412 62354 1440 62455
rect 1400 62348 1452 62354
rect 1400 62290 1452 62296
rect 1400 61736 1452 61742
rect 1398 61704 1400 61713
rect 1452 61704 1454 61713
rect 1398 61639 1454 61648
rect 1398 60888 1454 60897
rect 1398 60823 1454 60832
rect 1412 60654 1440 60823
rect 1400 60648 1452 60654
rect 1400 60590 1452 60596
rect 1400 60172 1452 60178
rect 1400 60114 1452 60120
rect 1412 59945 1440 60114
rect 1398 59936 1454 59945
rect 1398 59871 1454 59880
rect 1398 59120 1454 59129
rect 1398 59055 1400 59064
rect 1452 59055 1454 59064
rect 1400 59026 1452 59032
rect 1584 58880 1636 58886
rect 1584 58822 1636 58828
rect 1400 58472 1452 58478
rect 1400 58414 1452 58420
rect 1412 58313 1440 58414
rect 1398 58304 1454 58313
rect 1398 58239 1454 58248
rect 1398 57488 1454 57497
rect 1398 57423 1454 57432
rect 1412 57390 1440 57423
rect 1400 57384 1452 57390
rect 1400 57326 1452 57332
rect 1596 57050 1624 58822
rect 1584 57044 1636 57050
rect 1584 56986 1636 56992
rect 1400 56908 1452 56914
rect 1400 56850 1452 56856
rect 1412 56681 1440 56850
rect 1584 56704 1636 56710
rect 1398 56672 1454 56681
rect 1584 56646 1636 56652
rect 1398 56607 1454 56616
rect 1398 55856 1454 55865
rect 1398 55791 1400 55800
rect 1452 55791 1454 55800
rect 1400 55762 1452 55768
rect 1596 55758 1624 56646
rect 1584 55752 1636 55758
rect 1584 55694 1636 55700
rect 1400 55208 1452 55214
rect 1400 55150 1452 55156
rect 1412 55049 1440 55150
rect 1584 55072 1636 55078
rect 1398 55040 1454 55049
rect 1584 55014 1636 55020
rect 1398 54975 1454 54984
rect 1398 54224 1454 54233
rect 1398 54159 1454 54168
rect 1412 54126 1440 54159
rect 1400 54120 1452 54126
rect 1400 54062 1452 54068
rect 1400 53644 1452 53650
rect 1400 53586 1452 53592
rect 1412 53417 1440 53586
rect 1398 53408 1454 53417
rect 1398 53343 1454 53352
rect 1400 47592 1452 47598
rect 1398 47560 1400 47569
rect 1452 47560 1454 47569
rect 1398 47495 1454 47504
rect 1398 46744 1454 46753
rect 1398 46679 1454 46688
rect 1412 46578 1440 46679
rect 1400 46572 1452 46578
rect 1400 46514 1452 46520
rect 1596 40730 1624 55014
rect 1688 51066 1716 65350
rect 2056 58546 2084 79018
rect 3516 71460 3568 71466
rect 3516 71402 3568 71408
rect 3424 69828 3476 69834
rect 3424 69770 3476 69776
rect 2136 68740 2188 68746
rect 2136 68682 2188 68688
rect 2044 58540 2096 58546
rect 2044 58482 2096 58488
rect 1768 58336 1820 58342
rect 1768 58278 1820 58284
rect 1676 51060 1728 51066
rect 1676 51002 1728 51008
rect 1676 49700 1728 49706
rect 1676 49642 1728 49648
rect 1688 47666 1716 49642
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1780 44198 1808 58278
rect 1952 53984 2004 53990
rect 1952 53926 2004 53932
rect 1858 52592 1914 52601
rect 1858 52527 1860 52536
rect 1912 52527 1914 52536
rect 1860 52498 1912 52504
rect 1860 51876 1912 51882
rect 1860 51818 1912 51824
rect 1872 51785 1900 51818
rect 1858 51776 1914 51785
rect 1858 51711 1914 51720
rect 1858 50960 1914 50969
rect 1858 50895 1914 50904
rect 1872 50862 1900 50895
rect 1860 50856 1912 50862
rect 1860 50798 1912 50804
rect 1858 50008 1914 50017
rect 1858 49943 1914 49952
rect 1872 49774 1900 49943
rect 1860 49768 1912 49774
rect 1860 49710 1912 49716
rect 1860 49292 1912 49298
rect 1860 49234 1912 49240
rect 1872 49201 1900 49234
rect 1858 49192 1914 49201
rect 1858 49127 1914 49136
rect 1858 48376 1914 48385
rect 1858 48311 1914 48320
rect 1872 48278 1900 48311
rect 1860 48272 1912 48278
rect 1860 48214 1912 48220
rect 1860 46028 1912 46034
rect 1860 45970 1912 45976
rect 1872 45937 1900 45970
rect 1858 45928 1914 45937
rect 1858 45863 1914 45872
rect 1858 45112 1914 45121
rect 1858 45047 1914 45056
rect 1872 45014 1900 45047
rect 1860 45008 1912 45014
rect 1860 44950 1912 44956
rect 1860 44328 1912 44334
rect 1858 44296 1860 44305
rect 1912 44296 1914 44305
rect 1858 44231 1914 44240
rect 1768 44192 1820 44198
rect 1768 44134 1820 44140
rect 1964 43994 1992 53926
rect 2148 50368 2176 68682
rect 3148 68332 3200 68338
rect 3148 68274 3200 68280
rect 2228 66496 2280 66502
rect 2228 66438 2280 66444
rect 2240 55214 2268 66438
rect 2240 55186 2360 55214
rect 2148 50340 2268 50368
rect 2044 49224 2096 49230
rect 2044 49166 2096 49172
rect 2056 48278 2084 49166
rect 2044 48272 2096 48278
rect 2044 48214 2096 48220
rect 2044 47728 2096 47734
rect 2044 47670 2096 47676
rect 2056 46102 2084 47670
rect 2136 46504 2188 46510
rect 2136 46446 2188 46452
rect 2044 46096 2096 46102
rect 2044 46038 2096 46044
rect 2148 44470 2176 46446
rect 2240 44946 2268 50340
rect 2332 48278 2360 55186
rect 2872 54528 2924 54534
rect 2872 54470 2924 54476
rect 2320 48272 2372 48278
rect 2320 48214 2372 48220
rect 2596 47524 2648 47530
rect 2596 47466 2648 47472
rect 2320 46912 2372 46918
rect 2320 46854 2372 46860
rect 2332 45014 2360 46854
rect 2320 45008 2372 45014
rect 2320 44950 2372 44956
rect 2228 44940 2280 44946
rect 2228 44882 2280 44888
rect 2136 44464 2188 44470
rect 2136 44406 2188 44412
rect 1952 43988 2004 43994
rect 1952 43930 2004 43936
rect 1858 43480 1914 43489
rect 1858 43415 1914 43424
rect 2044 43444 2096 43450
rect 1872 43246 1900 43415
rect 2044 43386 2096 43392
rect 1860 43240 1912 43246
rect 1860 43182 1912 43188
rect 2056 42770 2084 43386
rect 2136 43240 2188 43246
rect 2136 43182 2188 43188
rect 1860 42764 1912 42770
rect 1860 42706 1912 42712
rect 2044 42764 2096 42770
rect 2044 42706 2096 42712
rect 1872 42673 1900 42706
rect 1858 42664 1914 42673
rect 1858 42599 1914 42608
rect 2044 42628 2096 42634
rect 2044 42570 2096 42576
rect 1858 41848 1914 41857
rect 1858 41783 1914 41792
rect 1872 41750 1900 41783
rect 1860 41744 1912 41750
rect 1860 41686 1912 41692
rect 1860 41064 1912 41070
rect 1858 41032 1860 41041
rect 1912 41032 1914 41041
rect 1858 40967 1914 40976
rect 1584 40724 1636 40730
rect 1584 40666 1636 40672
rect 1858 40080 1914 40089
rect 2056 40050 2084 42570
rect 2148 41206 2176 43182
rect 2136 41200 2188 41206
rect 2136 41142 2188 41148
rect 1858 40015 1914 40024
rect 2044 40044 2096 40050
rect 1872 39982 1900 40015
rect 2044 39986 2096 39992
rect 1860 39976 1912 39982
rect 1860 39918 1912 39924
rect 2136 39568 2188 39574
rect 2136 39510 2188 39516
rect 1860 39500 1912 39506
rect 1860 39442 1912 39448
rect 1872 39273 1900 39442
rect 2044 39432 2096 39438
rect 2044 39374 2096 39380
rect 1858 39264 1914 39273
rect 1858 39199 1914 39208
rect 2056 38486 2084 39374
rect 1860 38480 1912 38486
rect 1858 38448 1860 38457
rect 2044 38480 2096 38486
rect 1912 38448 1914 38457
rect 2044 38422 2096 38428
rect 1858 38383 1914 38392
rect 1584 38276 1636 38282
rect 1584 38218 1636 38224
rect 1596 36922 1624 38218
rect 2148 37942 2176 39510
rect 2504 38004 2556 38010
rect 2504 37946 2556 37952
rect 2136 37936 2188 37942
rect 2136 37878 2188 37884
rect 1676 37868 1728 37874
rect 1676 37810 1728 37816
rect 1584 36916 1636 36922
rect 1584 36858 1636 36864
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1412 36718 1440 36751
rect 1400 36712 1452 36718
rect 1400 36654 1452 36660
rect 1688 36378 1716 37810
rect 1860 37732 1912 37738
rect 1860 37674 1912 37680
rect 1872 37641 1900 37674
rect 1858 37632 1914 37641
rect 1858 37567 1914 37576
rect 1676 36372 1728 36378
rect 1676 36314 1728 36320
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1400 36236 1452 36242
rect 1400 36178 1452 36184
rect 1412 36009 1440 36178
rect 1398 36000 1454 36009
rect 1398 35935 1454 35944
rect 1398 35184 1454 35193
rect 1398 35119 1400 35128
rect 1452 35119 1454 35128
rect 1400 35090 1452 35096
rect 1780 34746 1808 36314
rect 2044 36304 2096 36310
rect 2044 36246 2096 36252
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 1412 34377 1440 34478
rect 1398 34368 1454 34377
rect 1398 34303 1454 34312
rect 2056 33590 2084 36246
rect 2516 35290 2544 37946
rect 2504 35284 2556 35290
rect 2504 35226 2556 35232
rect 2412 35216 2464 35222
rect 2412 35158 2464 35164
rect 2136 33856 2188 33862
rect 2136 33798 2188 33804
rect 2044 33584 2096 33590
rect 1858 33552 1914 33561
rect 2044 33526 2096 33532
rect 1858 33487 1914 33496
rect 1872 33454 1900 33487
rect 1860 33448 1912 33454
rect 1860 33390 1912 33396
rect 1952 33448 2004 33454
rect 1952 33390 2004 33396
rect 1964 33114 1992 33390
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1860 33040 1912 33046
rect 1860 32982 1912 32988
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1412 32745 1440 32914
rect 1584 32904 1636 32910
rect 1584 32846 1636 32852
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 1596 32026 1624 32846
rect 1584 32020 1636 32026
rect 1584 31962 1636 31968
rect 1398 31920 1454 31929
rect 1398 31855 1400 31864
rect 1452 31855 1454 31864
rect 1400 31826 1452 31832
rect 1872 31482 1900 32982
rect 1860 31476 1912 31482
rect 1860 31418 1912 31424
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1400 31272 1452 31278
rect 1400 31214 1452 31220
rect 1412 31113 1440 31214
rect 1398 31104 1454 31113
rect 1398 31039 1454 31048
rect 1216 30252 1268 30258
rect 1216 30194 1268 30200
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 664 3120 716 3126
rect 664 3062 716 3068
rect 112 3052 164 3058
rect 112 2994 164 3000
rect 124 800 152 2994
rect 388 2508 440 2514
rect 388 2450 440 2456
rect 400 800 428 2450
rect 676 800 704 3062
rect 952 800 980 3878
rect 1136 2258 1164 4422
rect 1228 3058 1256 30194
rect 1400 30184 1452 30190
rect 1398 30152 1400 30161
rect 1452 30152 1454 30161
rect 1398 30087 1454 30096
rect 1676 29640 1728 29646
rect 1676 29582 1728 29588
rect 1398 29336 1454 29345
rect 1398 29271 1454 29280
rect 1412 29102 1440 29271
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1688 28626 1716 29582
rect 1676 28620 1728 28626
rect 1676 28562 1728 28568
rect 1400 28552 1452 28558
rect 1398 28520 1400 28529
rect 1452 28520 1454 28529
rect 1398 28455 1454 28464
rect 1858 27704 1914 27713
rect 1858 27639 1914 27648
rect 1872 27606 1900 27639
rect 2056 27606 2084 31282
rect 1860 27600 1912 27606
rect 1860 27542 1912 27548
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 2148 27418 2176 33798
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 2056 27390 2176 27418
rect 1858 26888 1914 26897
rect 1858 26823 1860 26832
rect 1912 26823 1914 26832
rect 1860 26794 1912 26800
rect 1858 26072 1914 26081
rect 1858 26007 1914 26016
rect 1872 25838 1900 26007
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 2056 25430 2084 27390
rect 2136 27328 2188 27334
rect 2136 27270 2188 27276
rect 2044 25424 2096 25430
rect 2044 25366 2096 25372
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1872 25265 1900 25298
rect 1858 25256 1914 25265
rect 1858 25191 1914 25200
rect 1584 24880 1636 24886
rect 1584 24822 1636 24828
rect 1398 22808 1454 22817
rect 1596 22778 1624 24822
rect 1858 24440 1914 24449
rect 1858 24375 1914 24384
rect 1872 24342 1900 24375
rect 2148 24342 2176 27270
rect 1860 24336 1912 24342
rect 1860 24278 1912 24284
rect 2136 24336 2188 24342
rect 2136 24278 2188 24284
rect 1676 24132 1728 24138
rect 1676 24074 1728 24080
rect 1398 22743 1454 22752
rect 1584 22772 1636 22778
rect 1412 22574 1440 22743
rect 1584 22714 1636 22720
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1412 22001 1440 22034
rect 1398 21992 1454 22001
rect 1688 21962 1716 24074
rect 2240 23798 2268 27474
rect 2332 25974 2360 28154
rect 2424 27334 2452 35158
rect 2412 27328 2464 27334
rect 2412 27270 2464 27276
rect 2320 25968 2372 25974
rect 2320 25910 2372 25916
rect 2228 23792 2280 23798
rect 2228 23734 2280 23740
rect 1860 23656 1912 23662
rect 1858 23624 1860 23633
rect 1912 23624 1914 23633
rect 1858 23559 1914 23568
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 1398 21927 1454 21936
rect 1676 21956 1728 21962
rect 1676 21898 1728 21904
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1584 21412 1636 21418
rect 1584 21354 1636 21360
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1412 21010 1440 21111
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1596 20602 1624 21354
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1412 20233 1440 20334
rect 1398 20224 1454 20233
rect 1398 20159 1454 20168
rect 1398 19408 1454 19417
rect 1398 19343 1454 19352
rect 1584 19372 1636 19378
rect 1412 19310 1440 19343
rect 1584 19314 1636 19320
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18601 1440 18770
rect 1398 18592 1454 18601
rect 1398 18527 1454 18536
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1412 16969 1440 17070
rect 1398 16960 1454 16969
rect 1398 16895 1454 16904
rect 1504 16250 1532 19246
rect 1596 17338 1624 19314
rect 1688 17882 1716 21422
rect 1780 19174 1808 22442
rect 1860 19984 1912 19990
rect 1860 19926 1912 19932
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 1412 16046 1440 16079
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1688 15706 1716 17682
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 15337 1440 15506
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1398 14512 1454 14521
rect 1398 14447 1400 14456
rect 1452 14447 1454 14456
rect 1400 14418 1452 14424
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1780 13274 1808 15914
rect 1688 13246 1808 13274
rect 1398 12880 1454 12889
rect 1398 12815 1454 12824
rect 1412 12782 1440 12815
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 12073 1440 12242
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1398 11248 1454 11257
rect 1398 11183 1400 11192
rect 1452 11183 1454 11192
rect 1400 11154 1452 11160
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 1412 10130 1440 10231
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1400 9512 1452 9518
rect 1398 9480 1400 9489
rect 1452 9480 1454 9489
rect 1398 9415 1454 9424
rect 1398 8664 1454 8673
rect 1398 8599 1454 8608
rect 1412 8430 1440 8599
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1412 7857 1440 7890
rect 1584 7880 1636 7886
rect 1398 7848 1454 7857
rect 1584 7822 1636 7828
rect 1398 7783 1454 7792
rect 1398 7032 1454 7041
rect 1398 6967 1454 6976
rect 1412 6866 1440 6967
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1400 6248 1452 6254
rect 1398 6216 1400 6225
rect 1452 6216 1454 6225
rect 1398 6151 1454 6160
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1308 5160 1360 5166
rect 1308 5102 1360 5108
rect 1216 3052 1268 3058
rect 1216 2994 1268 3000
rect 1320 2961 1348 5102
rect 1412 4593 1440 5714
rect 1596 5370 1624 7822
rect 1688 6458 1716 13246
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 6730 1808 13126
rect 1872 12442 1900 19926
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2056 8090 2084 17138
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2042 5400 2098 5409
rect 1584 5364 1636 5370
rect 2042 5335 2098 5344
rect 1584 5306 1636 5312
rect 2056 5166 2084 5335
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1492 4004 1544 4010
rect 1492 3946 1544 3952
rect 1306 2952 1362 2961
rect 1306 2887 1362 2896
rect 1136 2230 1256 2258
rect 1228 800 1256 2230
rect 1504 800 1532 3946
rect 1964 2122 1992 4082
rect 2056 4078 2084 4422
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 1872 2094 1992 2122
rect 1872 800 1900 2094
rect 2148 800 2176 5714
rect 2240 5370 2268 10950
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2332 3738 2360 8026
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2424 800 2452 3674
rect 2516 3194 2544 6258
rect 2608 4078 2636 47466
rect 2780 46164 2832 46170
rect 2780 46106 2832 46112
rect 2792 45554 2820 46106
rect 2700 45526 2820 45554
rect 2700 43314 2728 45526
rect 2688 43308 2740 43314
rect 2688 43250 2740 43256
rect 2780 41812 2832 41818
rect 2780 41754 2832 41760
rect 2792 40066 2820 41754
rect 2700 40038 2820 40066
rect 2700 39642 2728 40038
rect 2688 39636 2740 39642
rect 2688 39578 2740 39584
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2792 30546 2820 31894
rect 2700 30518 2820 30546
rect 2700 29306 2728 30518
rect 2780 30388 2832 30394
rect 2780 30330 2832 30336
rect 2688 29300 2740 29306
rect 2688 29242 2740 29248
rect 2792 27690 2820 30330
rect 2700 27662 2820 27690
rect 2700 27062 2728 27662
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2688 27056 2740 27062
rect 2688 26998 2740 27004
rect 2792 23474 2820 27542
rect 2700 23446 2820 23474
rect 2700 21146 2728 23446
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2792 3777 2820 5102
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2700 800 2728 2450
rect 110 -800 166 800
rect 386 -800 442 800
rect 662 -800 718 800
rect 938 -800 994 800
rect 1214 -800 1270 800
rect 1490 -800 1546 800
rect 1858 -800 1914 800
rect 2134 -800 2190 800
rect 2410 -800 2466 800
rect 2686 -800 2742 800
rect 2792 513 2820 2858
rect 2884 2582 2912 54470
rect 2964 28620 3016 28626
rect 2964 28562 3016 28568
rect 2976 27674 3004 28562
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2976 19310 3004 24142
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2976 3534 3004 4422
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2976 800 3004 2926
rect 3068 1329 3096 3606
rect 3160 3058 3188 68274
rect 3436 53106 3464 69770
rect 3424 53100 3476 53106
rect 3424 53042 3476 53048
rect 3424 51400 3476 51406
rect 3424 51342 3476 51348
rect 3436 3738 3464 51342
rect 3528 45014 3556 71402
rect 3712 71058 3740 114514
rect 3804 112878 3832 114702
rect 3896 113830 3924 114838
rect 4220 114268 4516 114288
rect 4276 114266 4300 114268
rect 4356 114266 4380 114268
rect 4436 114266 4460 114268
rect 4298 114214 4300 114266
rect 4362 114214 4374 114266
rect 4436 114214 4438 114266
rect 4276 114212 4300 114214
rect 4356 114212 4380 114214
rect 4436 114212 4460 114214
rect 4220 114192 4516 114212
rect 4632 114170 4660 115602
rect 4712 115524 4764 115530
rect 4712 115466 4764 115472
rect 4620 114164 4672 114170
rect 4620 114106 4672 114112
rect 3884 113824 3936 113830
rect 3884 113766 3936 113772
rect 4724 113354 4752 115466
rect 4816 114510 4844 116690
rect 4804 114504 4856 114510
rect 4804 114446 4856 114452
rect 4712 113348 4764 113354
rect 4712 113290 4764 113296
rect 4220 113180 4516 113200
rect 4276 113178 4300 113180
rect 4356 113178 4380 113180
rect 4436 113178 4460 113180
rect 4298 113126 4300 113178
rect 4362 113126 4374 113178
rect 4436 113126 4438 113178
rect 4276 113124 4300 113126
rect 4356 113124 4380 113126
rect 4436 113124 4460 113126
rect 4220 113104 4516 113124
rect 4908 112878 4936 117642
rect 5000 114578 5028 117830
rect 5080 117156 5132 117162
rect 5080 117098 5132 117104
rect 5092 116006 5120 117098
rect 5184 116278 5212 119200
rect 5264 117088 5316 117094
rect 5264 117030 5316 117036
rect 5172 116272 5224 116278
rect 5172 116214 5224 116220
rect 5172 116136 5224 116142
rect 5172 116078 5224 116084
rect 5080 116000 5132 116006
rect 5080 115942 5132 115948
rect 5080 115660 5132 115666
rect 5080 115602 5132 115608
rect 4988 114572 5040 114578
rect 4988 114514 5040 114520
rect 5092 114374 5120 115602
rect 5080 114368 5132 114374
rect 5080 114310 5132 114316
rect 5184 113626 5212 116078
rect 5276 113626 5304 117030
rect 5368 115190 5396 119200
rect 5552 116872 5580 119200
rect 5552 116844 5764 116872
rect 5540 116748 5592 116754
rect 5540 116690 5592 116696
rect 5448 116068 5500 116074
rect 5448 116010 5500 116016
rect 5356 115184 5408 115190
rect 5356 115126 5408 115132
rect 5460 115122 5488 116010
rect 5552 115258 5580 116690
rect 5736 116226 5764 116844
rect 5828 116346 5856 119200
rect 5908 117088 5960 117094
rect 5908 117030 5960 117036
rect 5816 116340 5868 116346
rect 5816 116282 5868 116288
rect 5736 116198 5856 116226
rect 5724 116068 5776 116074
rect 5724 116010 5776 116016
rect 5632 116000 5684 116006
rect 5632 115942 5684 115948
rect 5540 115252 5592 115258
rect 5540 115194 5592 115200
rect 5644 115138 5672 115942
rect 5448 115116 5500 115122
rect 5448 115058 5500 115064
rect 5552 115110 5672 115138
rect 5552 115002 5580 115110
rect 5460 114974 5580 115002
rect 5632 114980 5684 114986
rect 5460 114102 5488 114974
rect 5632 114922 5684 114928
rect 5540 114572 5592 114578
rect 5540 114514 5592 114520
rect 5448 114096 5500 114102
rect 5448 114038 5500 114044
rect 5172 113620 5224 113626
rect 5172 113562 5224 113568
rect 5264 113620 5316 113626
rect 5264 113562 5316 113568
rect 5552 112878 5580 114514
rect 5644 114170 5672 114922
rect 5736 114510 5764 116010
rect 5724 114504 5776 114510
rect 5724 114446 5776 114452
rect 5632 114164 5684 114170
rect 5632 114106 5684 114112
rect 5828 112878 5856 116198
rect 5920 115598 5948 117030
rect 6012 116278 6040 119200
rect 6000 116272 6052 116278
rect 6000 116214 6052 116220
rect 5908 115592 5960 115598
rect 5908 115534 5960 115540
rect 6196 112962 6224 119200
rect 6472 116890 6500 119200
rect 6460 116884 6512 116890
rect 6460 116826 6512 116832
rect 6552 116612 6604 116618
rect 6552 116554 6604 116560
rect 6276 116068 6328 116074
rect 6276 116010 6328 116016
rect 6288 115258 6316 116010
rect 6276 115252 6328 115258
rect 6276 115194 6328 115200
rect 6276 115048 6328 115054
rect 6276 114990 6328 114996
rect 6288 113490 6316 114990
rect 6564 114578 6592 116554
rect 6656 116346 6684 119200
rect 6736 117156 6788 117162
rect 6736 117098 6788 117104
rect 6644 116340 6696 116346
rect 6644 116282 6696 116288
rect 6644 114708 6696 114714
rect 6644 114650 6696 114656
rect 6552 114572 6604 114578
rect 6552 114514 6604 114520
rect 6656 113558 6684 114650
rect 6644 113552 6696 113558
rect 6644 113494 6696 113500
rect 6276 113484 6328 113490
rect 6276 113426 6328 113432
rect 6748 113354 6776 117098
rect 6736 113348 6788 113354
rect 6736 113290 6788 113296
rect 6840 113014 6868 119200
rect 7024 116872 7052 119200
rect 7104 116884 7156 116890
rect 7024 116844 7104 116872
rect 7104 116826 7156 116832
rect 6920 116748 6972 116754
rect 6920 116690 6972 116696
rect 7012 116748 7064 116754
rect 7012 116690 7064 116696
rect 6932 115666 6960 116690
rect 6920 115660 6972 115666
rect 6920 115602 6972 115608
rect 7024 114510 7052 116690
rect 7300 115802 7328 119200
rect 7288 115796 7340 115802
rect 7288 115738 7340 115744
rect 7012 114504 7064 114510
rect 7012 114446 7064 114452
rect 7484 113558 7512 119200
rect 7668 116550 7696 119200
rect 7840 117224 7892 117230
rect 7840 117166 7892 117172
rect 7852 116822 7880 117166
rect 7840 116816 7892 116822
rect 7840 116758 7892 116764
rect 7656 116544 7708 116550
rect 7656 116486 7708 116492
rect 7564 116068 7616 116074
rect 7564 116010 7616 116016
rect 7748 116068 7800 116074
rect 7748 116010 7800 116016
rect 7576 114510 7604 116010
rect 7564 114504 7616 114510
rect 7564 114446 7616 114452
rect 7760 114170 7788 116010
rect 7944 115258 7972 119200
rect 8128 117314 8156 119200
rect 8128 117286 8248 117314
rect 8312 117298 8340 119200
rect 8116 117156 8168 117162
rect 8116 117098 8168 117104
rect 7932 115252 7984 115258
rect 7932 115194 7984 115200
rect 8024 114980 8076 114986
rect 8024 114922 8076 114928
rect 7748 114164 7800 114170
rect 7748 114106 7800 114112
rect 7472 113552 7524 113558
rect 7472 113494 7524 113500
rect 6828 113008 6880 113014
rect 6196 112934 6316 112962
rect 6828 112950 6880 112956
rect 6288 112878 6316 112934
rect 3792 112872 3844 112878
rect 3792 112814 3844 112820
rect 4896 112872 4948 112878
rect 4896 112814 4948 112820
rect 5540 112872 5592 112878
rect 5540 112814 5592 112820
rect 5816 112872 5868 112878
rect 5816 112814 5868 112820
rect 6276 112872 6328 112878
rect 6276 112814 6328 112820
rect 4220 112092 4516 112112
rect 4276 112090 4300 112092
rect 4356 112090 4380 112092
rect 4436 112090 4460 112092
rect 4298 112038 4300 112090
rect 4362 112038 4374 112090
rect 4436 112038 4438 112090
rect 4276 112036 4300 112038
rect 4356 112036 4380 112038
rect 4436 112036 4460 112038
rect 4220 112016 4516 112036
rect 7656 111240 7708 111246
rect 7656 111182 7708 111188
rect 4220 111004 4516 111024
rect 4276 111002 4300 111004
rect 4356 111002 4380 111004
rect 4436 111002 4460 111004
rect 4298 110950 4300 111002
rect 4362 110950 4374 111002
rect 4436 110950 4438 111002
rect 4276 110948 4300 110950
rect 4356 110948 4380 110950
rect 4436 110948 4460 110950
rect 4220 110928 4516 110948
rect 4220 109916 4516 109936
rect 4276 109914 4300 109916
rect 4356 109914 4380 109916
rect 4436 109914 4460 109916
rect 4298 109862 4300 109914
rect 4362 109862 4374 109914
rect 4436 109862 4438 109914
rect 4276 109860 4300 109862
rect 4356 109860 4380 109862
rect 4436 109860 4460 109862
rect 4220 109840 4516 109860
rect 5264 109744 5316 109750
rect 5264 109686 5316 109692
rect 4220 108828 4516 108848
rect 4276 108826 4300 108828
rect 4356 108826 4380 108828
rect 4436 108826 4460 108828
rect 4298 108774 4300 108826
rect 4362 108774 4374 108826
rect 4436 108774 4438 108826
rect 4276 108772 4300 108774
rect 4356 108772 4380 108774
rect 4436 108772 4460 108774
rect 4220 108752 4516 108772
rect 4220 107740 4516 107760
rect 4276 107738 4300 107740
rect 4356 107738 4380 107740
rect 4436 107738 4460 107740
rect 4298 107686 4300 107738
rect 4362 107686 4374 107738
rect 4436 107686 4438 107738
rect 4276 107684 4300 107686
rect 4356 107684 4380 107686
rect 4436 107684 4460 107686
rect 4220 107664 4516 107684
rect 4220 106652 4516 106672
rect 4276 106650 4300 106652
rect 4356 106650 4380 106652
rect 4436 106650 4460 106652
rect 4298 106598 4300 106650
rect 4362 106598 4374 106650
rect 4436 106598 4438 106650
rect 4276 106596 4300 106598
rect 4356 106596 4380 106598
rect 4436 106596 4460 106598
rect 4220 106576 4516 106596
rect 4220 105564 4516 105584
rect 4276 105562 4300 105564
rect 4356 105562 4380 105564
rect 4436 105562 4460 105564
rect 4298 105510 4300 105562
rect 4362 105510 4374 105562
rect 4436 105510 4438 105562
rect 4276 105508 4300 105510
rect 4356 105508 4380 105510
rect 4436 105508 4460 105510
rect 4220 105488 4516 105508
rect 4220 104476 4516 104496
rect 4276 104474 4300 104476
rect 4356 104474 4380 104476
rect 4436 104474 4460 104476
rect 4298 104422 4300 104474
rect 4362 104422 4374 104474
rect 4436 104422 4438 104474
rect 4276 104420 4300 104422
rect 4356 104420 4380 104422
rect 4436 104420 4460 104422
rect 4220 104400 4516 104420
rect 4220 103388 4516 103408
rect 4276 103386 4300 103388
rect 4356 103386 4380 103388
rect 4436 103386 4460 103388
rect 4298 103334 4300 103386
rect 4362 103334 4374 103386
rect 4436 103334 4438 103386
rect 4276 103332 4300 103334
rect 4356 103332 4380 103334
rect 4436 103332 4460 103334
rect 4220 103312 4516 103332
rect 4804 103012 4856 103018
rect 4804 102954 4856 102960
rect 4220 102300 4516 102320
rect 4276 102298 4300 102300
rect 4356 102298 4380 102300
rect 4436 102298 4460 102300
rect 4298 102246 4300 102298
rect 4362 102246 4374 102298
rect 4436 102246 4438 102298
rect 4276 102244 4300 102246
rect 4356 102244 4380 102246
rect 4436 102244 4460 102246
rect 4220 102224 4516 102244
rect 4068 101380 4120 101386
rect 4068 101322 4120 101328
rect 4080 95946 4108 101322
rect 4220 101212 4516 101232
rect 4276 101210 4300 101212
rect 4356 101210 4380 101212
rect 4436 101210 4460 101212
rect 4298 101158 4300 101210
rect 4362 101158 4374 101210
rect 4436 101158 4438 101210
rect 4276 101156 4300 101158
rect 4356 101156 4380 101158
rect 4436 101156 4460 101158
rect 4220 101136 4516 101156
rect 4220 100124 4516 100144
rect 4276 100122 4300 100124
rect 4356 100122 4380 100124
rect 4436 100122 4460 100124
rect 4298 100070 4300 100122
rect 4362 100070 4374 100122
rect 4436 100070 4438 100122
rect 4276 100068 4300 100070
rect 4356 100068 4380 100070
rect 4436 100068 4460 100070
rect 4220 100048 4516 100068
rect 4220 99036 4516 99056
rect 4276 99034 4300 99036
rect 4356 99034 4380 99036
rect 4436 99034 4460 99036
rect 4298 98982 4300 99034
rect 4362 98982 4374 99034
rect 4436 98982 4438 99034
rect 4276 98980 4300 98982
rect 4356 98980 4380 98982
rect 4436 98980 4460 98982
rect 4220 98960 4516 98980
rect 4220 97948 4516 97968
rect 4276 97946 4300 97948
rect 4356 97946 4380 97948
rect 4436 97946 4460 97948
rect 4298 97894 4300 97946
rect 4362 97894 4374 97946
rect 4436 97894 4438 97946
rect 4276 97892 4300 97894
rect 4356 97892 4380 97894
rect 4436 97892 4460 97894
rect 4220 97872 4516 97892
rect 4220 96860 4516 96880
rect 4276 96858 4300 96860
rect 4356 96858 4380 96860
rect 4436 96858 4460 96860
rect 4298 96806 4300 96858
rect 4362 96806 4374 96858
rect 4436 96806 4438 96858
rect 4276 96804 4300 96806
rect 4356 96804 4380 96806
rect 4436 96804 4460 96806
rect 4220 96784 4516 96804
rect 4068 95940 4120 95946
rect 4068 95882 4120 95888
rect 4220 95772 4516 95792
rect 4276 95770 4300 95772
rect 4356 95770 4380 95772
rect 4436 95770 4460 95772
rect 4298 95718 4300 95770
rect 4362 95718 4374 95770
rect 4436 95718 4438 95770
rect 4276 95716 4300 95718
rect 4356 95716 4380 95718
rect 4436 95716 4460 95718
rect 4220 95696 4516 95716
rect 4220 94684 4516 94704
rect 4276 94682 4300 94684
rect 4356 94682 4380 94684
rect 4436 94682 4460 94684
rect 4298 94630 4300 94682
rect 4362 94630 4374 94682
rect 4436 94630 4438 94682
rect 4276 94628 4300 94630
rect 4356 94628 4380 94630
rect 4436 94628 4460 94630
rect 4220 94608 4516 94628
rect 4220 93596 4516 93616
rect 4276 93594 4300 93596
rect 4356 93594 4380 93596
rect 4436 93594 4460 93596
rect 4298 93542 4300 93594
rect 4362 93542 4374 93594
rect 4436 93542 4438 93594
rect 4276 93540 4300 93542
rect 4356 93540 4380 93542
rect 4436 93540 4460 93542
rect 4220 93520 4516 93540
rect 4220 92508 4516 92528
rect 4276 92506 4300 92508
rect 4356 92506 4380 92508
rect 4436 92506 4460 92508
rect 4298 92454 4300 92506
rect 4362 92454 4374 92506
rect 4436 92454 4438 92506
rect 4276 92452 4300 92454
rect 4356 92452 4380 92454
rect 4436 92452 4460 92454
rect 4220 92432 4516 92452
rect 4220 91420 4516 91440
rect 4276 91418 4300 91420
rect 4356 91418 4380 91420
rect 4436 91418 4460 91420
rect 4298 91366 4300 91418
rect 4362 91366 4374 91418
rect 4436 91366 4438 91418
rect 4276 91364 4300 91366
rect 4356 91364 4380 91366
rect 4436 91364 4460 91366
rect 4220 91344 4516 91364
rect 4220 90332 4516 90352
rect 4276 90330 4300 90332
rect 4356 90330 4380 90332
rect 4436 90330 4460 90332
rect 4298 90278 4300 90330
rect 4362 90278 4374 90330
rect 4436 90278 4438 90330
rect 4276 90276 4300 90278
rect 4356 90276 4380 90278
rect 4436 90276 4460 90278
rect 4220 90256 4516 90276
rect 4220 89244 4516 89264
rect 4276 89242 4300 89244
rect 4356 89242 4380 89244
rect 4436 89242 4460 89244
rect 4298 89190 4300 89242
rect 4362 89190 4374 89242
rect 4436 89190 4438 89242
rect 4276 89188 4300 89190
rect 4356 89188 4380 89190
rect 4436 89188 4460 89190
rect 4220 89168 4516 89188
rect 4220 88156 4516 88176
rect 4276 88154 4300 88156
rect 4356 88154 4380 88156
rect 4436 88154 4460 88156
rect 4298 88102 4300 88154
rect 4362 88102 4374 88154
rect 4436 88102 4438 88154
rect 4276 88100 4300 88102
rect 4356 88100 4380 88102
rect 4436 88100 4460 88102
rect 4220 88080 4516 88100
rect 4220 87068 4516 87088
rect 4276 87066 4300 87068
rect 4356 87066 4380 87068
rect 4436 87066 4460 87068
rect 4298 87014 4300 87066
rect 4362 87014 4374 87066
rect 4436 87014 4438 87066
rect 4276 87012 4300 87014
rect 4356 87012 4380 87014
rect 4436 87012 4460 87014
rect 4220 86992 4516 87012
rect 4816 86970 4844 102954
rect 4988 98252 5040 98258
rect 4988 98194 5040 98200
rect 4804 86964 4856 86970
rect 4804 86906 4856 86912
rect 4220 85980 4516 86000
rect 4276 85978 4300 85980
rect 4356 85978 4380 85980
rect 4436 85978 4460 85980
rect 4298 85926 4300 85978
rect 4362 85926 4374 85978
rect 4436 85926 4438 85978
rect 4276 85924 4300 85926
rect 4356 85924 4380 85926
rect 4436 85924 4460 85926
rect 4220 85904 4516 85924
rect 4220 84892 4516 84912
rect 4276 84890 4300 84892
rect 4356 84890 4380 84892
rect 4436 84890 4460 84892
rect 4298 84838 4300 84890
rect 4362 84838 4374 84890
rect 4436 84838 4438 84890
rect 4276 84836 4300 84838
rect 4356 84836 4380 84838
rect 4436 84836 4460 84838
rect 4220 84816 4516 84836
rect 4068 83972 4120 83978
rect 4068 83914 4120 83920
rect 4080 80306 4108 83914
rect 4220 83804 4516 83824
rect 4276 83802 4300 83804
rect 4356 83802 4380 83804
rect 4436 83802 4460 83804
rect 4298 83750 4300 83802
rect 4362 83750 4374 83802
rect 4436 83750 4438 83802
rect 4276 83748 4300 83750
rect 4356 83748 4380 83750
rect 4436 83748 4460 83750
rect 4220 83728 4516 83748
rect 4220 82716 4516 82736
rect 4276 82714 4300 82716
rect 4356 82714 4380 82716
rect 4436 82714 4460 82716
rect 4298 82662 4300 82714
rect 4362 82662 4374 82714
rect 4436 82662 4438 82714
rect 4276 82660 4300 82662
rect 4356 82660 4380 82662
rect 4436 82660 4460 82662
rect 4220 82640 4516 82660
rect 4220 81628 4516 81648
rect 4276 81626 4300 81628
rect 4356 81626 4380 81628
rect 4436 81626 4460 81628
rect 4298 81574 4300 81626
rect 4362 81574 4374 81626
rect 4436 81574 4438 81626
rect 4276 81572 4300 81574
rect 4356 81572 4380 81574
rect 4436 81572 4460 81574
rect 4220 81552 4516 81572
rect 4220 80540 4516 80560
rect 4276 80538 4300 80540
rect 4356 80538 4380 80540
rect 4436 80538 4460 80540
rect 4298 80486 4300 80538
rect 4362 80486 4374 80538
rect 4436 80486 4438 80538
rect 4276 80484 4300 80486
rect 4356 80484 4380 80486
rect 4436 80484 4460 80486
rect 4220 80464 4516 80484
rect 4068 80300 4120 80306
rect 4068 80242 4120 80248
rect 4220 79452 4516 79472
rect 4276 79450 4300 79452
rect 4356 79450 4380 79452
rect 4436 79450 4460 79452
rect 4298 79398 4300 79450
rect 4362 79398 4374 79450
rect 4436 79398 4438 79450
rect 4276 79396 4300 79398
rect 4356 79396 4380 79398
rect 4436 79396 4460 79398
rect 4220 79376 4516 79396
rect 4220 78364 4516 78384
rect 4276 78362 4300 78364
rect 4356 78362 4380 78364
rect 4436 78362 4460 78364
rect 4298 78310 4300 78362
rect 4362 78310 4374 78362
rect 4436 78310 4438 78362
rect 4276 78308 4300 78310
rect 4356 78308 4380 78310
rect 4436 78308 4460 78310
rect 4220 78288 4516 78308
rect 4220 77276 4516 77296
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4298 77222 4300 77274
rect 4362 77222 4374 77274
rect 4436 77222 4438 77274
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4220 77200 4516 77220
rect 4220 76188 4516 76208
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4298 76134 4300 76186
rect 4362 76134 4374 76186
rect 4436 76134 4438 76186
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4220 76112 4516 76132
rect 4220 75100 4516 75120
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4298 75046 4300 75098
rect 4362 75046 4374 75098
rect 4436 75046 4438 75098
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4220 75024 4516 75044
rect 4220 74012 4516 74032
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4298 73958 4300 74010
rect 4362 73958 4374 74010
rect 4436 73958 4438 74010
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4220 73936 4516 73956
rect 4220 72924 4516 72944
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4298 72870 4300 72922
rect 4362 72870 4374 72922
rect 4436 72870 4438 72922
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4220 72848 4516 72868
rect 4804 72548 4856 72554
rect 4804 72490 4856 72496
rect 4220 71836 4516 71856
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4298 71782 4300 71834
rect 4362 71782 4374 71834
rect 4436 71782 4438 71834
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4220 71760 4516 71780
rect 3700 71052 3752 71058
rect 3700 70994 3752 71000
rect 4220 70748 4516 70768
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4298 70694 4300 70746
rect 4362 70694 4374 70746
rect 4436 70694 4438 70746
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4220 70672 4516 70692
rect 4220 69660 4516 69680
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4298 69606 4300 69658
rect 4362 69606 4374 69658
rect 4436 69606 4438 69658
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4220 69584 4516 69604
rect 4220 68572 4516 68592
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4298 68518 4300 68570
rect 4362 68518 4374 68570
rect 4436 68518 4438 68570
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4220 68496 4516 68516
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 4220 59868 4516 59888
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 3608 57248 3660 57254
rect 3608 57190 3660 57196
rect 3516 45008 3568 45014
rect 3516 44950 3568 44956
rect 3620 42158 3648 57190
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 4068 50856 4120 50862
rect 4068 50798 4120 50804
rect 4080 46578 4108 50798
rect 4620 50788 4672 50794
rect 4620 50730 4672 50736
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4068 46572 4120 46578
rect 4068 46514 4120 46520
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 3608 42152 3660 42158
rect 3608 42094 3660 42100
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 5914 3556 14758
rect 3620 14074 3648 21966
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3054 1320 3110 1329
rect 3054 1255 3110 1264
rect 3252 800 3280 3334
rect 3344 2145 3372 3470
rect 3330 2136 3386 2145
rect 3330 2071 3386 2080
rect 3620 800 3648 3946
rect 4080 3670 4108 11698
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4632 3194 4660 50730
rect 4816 47258 4844 72490
rect 4896 55616 4948 55622
rect 4896 55558 4948 55564
rect 4804 47252 4856 47258
rect 4804 47194 4856 47200
rect 4908 40662 4936 55558
rect 4896 40656 4948 40662
rect 4896 40598 4948 40604
rect 4804 35216 4856 35222
rect 4804 35158 4856 35164
rect 4712 32360 4764 32366
rect 4712 32302 4764 32308
rect 4724 30326 4752 32302
rect 4712 30320 4764 30326
rect 4712 30262 4764 30268
rect 4816 26234 4844 35158
rect 4896 29572 4948 29578
rect 4896 29514 4948 29520
rect 4724 26206 4844 26234
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3896 800 3924 2450
rect 4172 2394 4200 2926
rect 4264 2650 4292 3062
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4080 2366 4200 2394
rect 4080 1986 4108 2366
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4080 1958 4200 1986
rect 4172 800 4200 1958
rect 4632 1442 4660 2790
rect 4724 2582 4752 26206
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4816 18970 4844 25638
rect 4908 24886 4936 29514
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4816 17202 4844 18226
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5000 5710 5028 98194
rect 5080 57044 5132 57050
rect 5080 56986 5132 56992
rect 5092 41682 5120 56986
rect 5080 41676 5132 41682
rect 5080 41618 5132 41624
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 2122 4844 3946
rect 4908 3942 4936 5510
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4448 1414 4660 1442
rect 4724 2094 4844 2122
rect 4448 800 4476 1414
rect 4724 800 4752 2094
rect 5000 800 5028 3538
rect 5092 2990 5120 6122
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 3126 5212 3334
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5276 2582 5304 109686
rect 7564 108452 7616 108458
rect 7564 108394 7616 108400
rect 6184 103080 6236 103086
rect 6184 103022 6236 103028
rect 6828 103080 6880 103086
rect 6828 103022 6880 103028
rect 5724 101516 5776 101522
rect 5724 101458 5776 101464
rect 5736 100026 5764 101458
rect 5724 100020 5776 100026
rect 5724 99962 5776 99968
rect 5540 44192 5592 44198
rect 5540 44134 5592 44140
rect 5552 41750 5580 44134
rect 5540 41744 5592 41750
rect 5540 41686 5592 41692
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5552 19378 5580 24346
rect 5644 21486 5672 25230
rect 5724 24608 5776 24614
rect 5724 24550 5776 24556
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5736 17746 5764 24550
rect 5828 22506 5856 27814
rect 5816 22500 5868 22506
rect 5816 22442 5868 22448
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5368 800 5396 3538
rect 5552 2650 5580 5646
rect 5828 2990 5856 16662
rect 6196 5098 6224 103022
rect 6276 99748 6328 99754
rect 6276 99690 6328 99696
rect 6288 89554 6316 99690
rect 6840 97306 6868 103022
rect 7576 102474 7604 108394
rect 7564 102468 7616 102474
rect 7564 102410 7616 102416
rect 6828 97300 6880 97306
rect 6828 97242 6880 97248
rect 6276 89548 6328 89554
rect 6276 89490 6328 89496
rect 6276 73228 6328 73234
rect 6276 73170 6328 73176
rect 6288 46102 6316 73170
rect 6368 70916 6420 70922
rect 6368 70858 6420 70864
rect 6276 46096 6328 46102
rect 6276 46038 6328 46044
rect 6380 45082 6408 70858
rect 7564 63776 7616 63782
rect 7564 63718 7616 63724
rect 6552 60512 6604 60518
rect 6552 60454 6604 60460
rect 6460 55752 6512 55758
rect 6460 55694 6512 55700
rect 6368 45076 6420 45082
rect 6368 45018 6420 45024
rect 6472 41138 6500 55694
rect 6564 44402 6592 60454
rect 7288 59152 7340 59158
rect 7288 59094 7340 59100
rect 7012 57044 7064 57050
rect 7012 56986 7064 56992
rect 6736 55888 6788 55894
rect 6736 55830 6788 55836
rect 6552 44396 6604 44402
rect 6552 44338 6604 44344
rect 6460 41132 6512 41138
rect 6460 41074 6512 41080
rect 6276 38956 6328 38962
rect 6276 38898 6328 38904
rect 6288 27538 6316 38898
rect 6368 38344 6420 38350
rect 6368 38286 6420 38292
rect 6380 28218 6408 38286
rect 6552 29028 6604 29034
rect 6552 28970 6604 28976
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6276 27532 6328 27538
rect 6276 27474 6328 27480
rect 6564 24138 6592 28970
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6288 8090 6316 19790
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6380 5370 6408 14350
rect 6472 12986 6500 20878
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 800 5672 2790
rect 5920 800 5948 4014
rect 6748 3058 6776 55830
rect 7024 50998 7052 56986
rect 7012 50992 7064 50998
rect 7012 50934 7064 50940
rect 7300 50386 7328 59094
rect 7288 50380 7340 50386
rect 7288 50322 7340 50328
rect 7300 48686 7328 50322
rect 7472 50176 7524 50182
rect 7472 50118 7524 50124
rect 7288 48680 7340 48686
rect 7288 48622 7340 48628
rect 7300 47598 7328 48622
rect 7380 48544 7432 48550
rect 7380 48486 7432 48492
rect 7012 47592 7064 47598
rect 7012 47534 7064 47540
rect 7288 47592 7340 47598
rect 7288 47534 7340 47540
rect 7024 46510 7052 47534
rect 7288 47456 7340 47462
rect 7288 47398 7340 47404
rect 7012 46504 7064 46510
rect 7012 46446 7064 46452
rect 7196 46368 7248 46374
rect 7196 46310 7248 46316
rect 7208 42158 7236 46310
rect 7300 45422 7328 47398
rect 7392 45490 7420 48486
rect 7484 48142 7512 50118
rect 7472 48136 7524 48142
rect 7472 48078 7524 48084
rect 7484 47666 7512 48078
rect 7472 47660 7524 47666
rect 7472 47602 7524 47608
rect 7484 47054 7512 47602
rect 7576 47122 7604 63718
rect 7668 59158 7696 111182
rect 7748 106956 7800 106962
rect 7748 106898 7800 106904
rect 7760 102134 7788 106898
rect 7748 102128 7800 102134
rect 7748 102070 7800 102076
rect 7748 67040 7800 67046
rect 7748 66982 7800 66988
rect 7656 59152 7708 59158
rect 7656 59094 7708 59100
rect 7656 51536 7708 51542
rect 7656 51478 7708 51484
rect 7668 49706 7696 51478
rect 7760 49706 7788 66982
rect 8036 62830 8064 114922
rect 8128 113354 8156 117098
rect 8220 114578 8248 117286
rect 8300 117292 8352 117298
rect 8300 117234 8352 117240
rect 8392 117156 8444 117162
rect 8392 117098 8444 117104
rect 8404 115802 8432 117098
rect 8588 116890 8616 119200
rect 8576 116884 8628 116890
rect 8576 116826 8628 116832
rect 8576 116748 8628 116754
rect 8576 116690 8628 116696
rect 8392 115796 8444 115802
rect 8392 115738 8444 115744
rect 8392 114912 8444 114918
rect 8392 114854 8444 114860
rect 8208 114572 8260 114578
rect 8208 114514 8260 114520
rect 8300 114436 8352 114442
rect 8300 114378 8352 114384
rect 8312 113626 8340 114378
rect 8404 113898 8432 114854
rect 8588 114510 8616 116690
rect 8668 115728 8720 115734
rect 8668 115670 8720 115676
rect 8576 114504 8628 114510
rect 8576 114446 8628 114452
rect 8392 113892 8444 113898
rect 8392 113834 8444 113840
rect 8300 113620 8352 113626
rect 8300 113562 8352 113568
rect 8208 113552 8260 113558
rect 8260 113500 8432 113506
rect 8208 113494 8432 113500
rect 8220 113490 8432 113494
rect 8220 113484 8444 113490
rect 8220 113478 8392 113484
rect 8392 113426 8444 113432
rect 8116 113348 8168 113354
rect 8116 113290 8168 113296
rect 8680 109274 8708 115670
rect 8772 113966 8800 119200
rect 8956 117298 8984 119200
rect 9140 117586 9168 119200
rect 9140 117558 9352 117586
rect 8944 117292 8996 117298
rect 8944 117234 8996 117240
rect 9324 116890 9352 117558
rect 9312 116884 9364 116890
rect 9312 116826 9364 116832
rect 9416 114986 9444 119200
rect 9600 117230 9628 119200
rect 9784 117858 9812 119200
rect 9692 117830 9812 117858
rect 9588 117224 9640 117230
rect 9588 117166 9640 117172
rect 9496 117156 9548 117162
rect 9496 117098 9548 117104
rect 9508 116210 9536 117098
rect 9692 116822 9720 117830
rect 9772 117156 9824 117162
rect 9772 117098 9824 117104
rect 9680 116816 9732 116822
rect 9680 116758 9732 116764
rect 9496 116204 9548 116210
rect 9496 116146 9548 116152
rect 9784 115802 9812 117098
rect 9864 116748 9916 116754
rect 9864 116690 9916 116696
rect 9772 115796 9824 115802
rect 9772 115738 9824 115744
rect 9876 115258 9904 116690
rect 10060 115462 10088 119200
rect 10244 117298 10272 119200
rect 10232 117292 10284 117298
rect 10232 117234 10284 117240
rect 10428 116346 10456 119200
rect 10600 116748 10652 116754
rect 10600 116690 10652 116696
rect 10416 116340 10468 116346
rect 10416 116282 10468 116288
rect 10048 115456 10100 115462
rect 10048 115398 10100 115404
rect 10612 115258 10640 116690
rect 9864 115252 9916 115258
rect 9864 115194 9916 115200
rect 10600 115252 10652 115258
rect 10600 115194 10652 115200
rect 10704 115122 10732 119200
rect 10888 117230 10916 119200
rect 10876 117224 10928 117230
rect 10876 117166 10928 117172
rect 11072 116346 11100 119200
rect 11256 117314 11284 119200
rect 11256 117286 11468 117314
rect 11532 117298 11560 119200
rect 11152 117156 11204 117162
rect 11152 117098 11204 117104
rect 11336 117156 11388 117162
rect 11336 117098 11388 117104
rect 11060 116340 11112 116346
rect 11060 116282 11112 116288
rect 10968 116068 11020 116074
rect 10968 116010 11020 116016
rect 10876 115456 10928 115462
rect 10876 115398 10928 115404
rect 9864 115116 9916 115122
rect 9864 115058 9916 115064
rect 10692 115116 10744 115122
rect 10692 115058 10744 115064
rect 9404 114980 9456 114986
rect 9404 114922 9456 114928
rect 9876 114374 9904 115058
rect 10508 114980 10560 114986
rect 10508 114922 10560 114928
rect 10416 114708 10468 114714
rect 10416 114650 10468 114656
rect 9864 114368 9916 114374
rect 9864 114310 9916 114316
rect 10428 114034 10456 114650
rect 10520 114578 10548 114922
rect 10888 114578 10916 115398
rect 10980 115258 11008 116010
rect 11164 115802 11192 117098
rect 11244 116068 11296 116074
rect 11244 116010 11296 116016
rect 11152 115796 11204 115802
rect 11152 115738 11204 115744
rect 11256 115258 11284 116010
rect 11348 115734 11376 117098
rect 11336 115728 11388 115734
rect 11336 115670 11388 115676
rect 10968 115252 11020 115258
rect 10968 115194 11020 115200
rect 11244 115252 11296 115258
rect 11244 115194 11296 115200
rect 10968 115048 11020 115054
rect 10968 114990 11020 114996
rect 10508 114572 10560 114578
rect 10508 114514 10560 114520
rect 10876 114572 10928 114578
rect 10876 114514 10928 114520
rect 10980 114374 11008 114990
rect 11440 114578 11468 117286
rect 11520 117292 11572 117298
rect 11520 117234 11572 117240
rect 11716 116890 11744 119200
rect 11704 116884 11756 116890
rect 11704 116826 11756 116832
rect 11900 114986 11928 119200
rect 12176 117094 12204 119200
rect 12164 117088 12216 117094
rect 12164 117030 12216 117036
rect 12360 116872 12388 119200
rect 12440 116884 12492 116890
rect 12360 116844 12440 116872
rect 12440 116826 12492 116832
rect 12164 116748 12216 116754
rect 12164 116690 12216 116696
rect 12176 115666 12204 116690
rect 12164 115660 12216 115666
rect 12164 115602 12216 115608
rect 11888 114980 11940 114986
rect 11888 114922 11940 114928
rect 12544 114918 12572 119200
rect 12820 117366 12848 119200
rect 13004 117450 13032 119200
rect 13188 117586 13216 119200
rect 13188 117558 13308 117586
rect 13004 117422 13216 117450
rect 12808 117360 12860 117366
rect 12808 117302 12860 117308
rect 13084 117156 13136 117162
rect 13084 117098 13136 117104
rect 12900 116748 12952 116754
rect 12900 116690 12952 116696
rect 12992 116748 13044 116754
rect 12992 116690 13044 116696
rect 12912 115666 12940 116690
rect 12900 115660 12952 115666
rect 12900 115602 12952 115608
rect 13004 115258 13032 116690
rect 13096 116210 13124 117098
rect 13188 116822 13216 117422
rect 13176 116816 13228 116822
rect 13176 116758 13228 116764
rect 13084 116204 13136 116210
rect 13084 116146 13136 116152
rect 12992 115252 13044 115258
rect 12992 115194 13044 115200
rect 12900 114980 12952 114986
rect 12900 114922 12952 114928
rect 12532 114912 12584 114918
rect 12532 114854 12584 114860
rect 12912 114578 12940 114922
rect 13280 114578 13308 117558
rect 13464 117094 13492 119200
rect 13452 117088 13504 117094
rect 13452 117030 13504 117036
rect 13648 116890 13676 119200
rect 13832 117280 13860 119200
rect 14016 117366 14044 119200
rect 14004 117360 14056 117366
rect 14004 117302 14056 117308
rect 13832 117252 13952 117280
rect 13820 117156 13872 117162
rect 13820 117098 13872 117104
rect 13636 116884 13688 116890
rect 13636 116826 13688 116832
rect 13832 116142 13860 117098
rect 13820 116136 13872 116142
rect 13820 116078 13872 116084
rect 13544 114912 13596 114918
rect 13544 114854 13596 114860
rect 13556 114578 13584 114854
rect 13924 114578 13952 117252
rect 14096 117224 14148 117230
rect 14096 117166 14148 117172
rect 14108 115802 14136 117166
rect 14292 116822 14320 119200
rect 14280 116816 14332 116822
rect 14280 116758 14332 116764
rect 14372 116748 14424 116754
rect 14372 116690 14424 116696
rect 14096 115796 14148 115802
rect 14096 115738 14148 115744
rect 14384 115258 14412 116690
rect 14372 115252 14424 115258
rect 14372 115194 14424 115200
rect 14476 114714 14504 119200
rect 14660 116686 14688 119200
rect 14936 117586 14964 119200
rect 14752 117558 14964 117586
rect 14752 116890 14780 117558
rect 15120 117280 15148 119200
rect 15304 117450 15332 119200
rect 15304 117422 15424 117450
rect 15396 117366 15424 117422
rect 15384 117360 15436 117366
rect 15384 117302 15436 117308
rect 14936 117252 15148 117280
rect 14740 116884 14792 116890
rect 14740 116826 14792 116832
rect 14648 116680 14700 116686
rect 14648 116622 14700 116628
rect 14464 114708 14516 114714
rect 14464 114650 14516 114656
rect 14936 114578 14964 117252
rect 15016 117156 15068 117162
rect 15016 117098 15068 117104
rect 15028 116210 15056 117098
rect 15580 116872 15608 119200
rect 15580 116844 15700 116872
rect 15108 116748 15160 116754
rect 15108 116690 15160 116696
rect 15568 116748 15620 116754
rect 15568 116690 15620 116696
rect 15016 116204 15068 116210
rect 15016 116146 15068 116152
rect 15120 115258 15148 116690
rect 15580 115258 15608 116690
rect 15672 116346 15700 116844
rect 15660 116340 15712 116346
rect 15660 116282 15712 116288
rect 15660 116068 15712 116074
rect 15660 116010 15712 116016
rect 15672 115258 15700 116010
rect 15108 115252 15160 115258
rect 15108 115194 15160 115200
rect 15568 115252 15620 115258
rect 15568 115194 15620 115200
rect 15660 115252 15712 115258
rect 15660 115194 15712 115200
rect 15292 115048 15344 115054
rect 15292 114990 15344 114996
rect 11428 114572 11480 114578
rect 11428 114514 11480 114520
rect 12900 114572 12952 114578
rect 12900 114514 12952 114520
rect 13268 114572 13320 114578
rect 13268 114514 13320 114520
rect 13544 114572 13596 114578
rect 13544 114514 13596 114520
rect 13912 114572 13964 114578
rect 13912 114514 13964 114520
rect 14924 114572 14976 114578
rect 14924 114514 14976 114520
rect 15304 114442 15332 114990
rect 15292 114436 15344 114442
rect 15292 114378 15344 114384
rect 10968 114368 11020 114374
rect 10968 114310 11020 114316
rect 13360 114368 13412 114374
rect 13360 114310 13412 114316
rect 14648 114368 14700 114374
rect 14648 114310 14700 114316
rect 10416 114028 10468 114034
rect 10416 113970 10468 113976
rect 8760 113960 8812 113966
rect 8760 113902 8812 113908
rect 13372 113422 13400 114310
rect 14660 113558 14688 114310
rect 15764 113966 15792 119200
rect 15948 117314 15976 119200
rect 15948 117286 16068 117314
rect 15844 117224 15896 117230
rect 15844 117166 15896 117172
rect 15856 115802 15884 117166
rect 15936 117156 15988 117162
rect 15936 117098 15988 117104
rect 15948 116142 15976 117098
rect 16040 116822 16068 117286
rect 16028 116816 16080 116822
rect 16028 116758 16080 116764
rect 16132 116278 16160 119200
rect 16304 117088 16356 117094
rect 16304 117030 16356 117036
rect 16316 116686 16344 117030
rect 16304 116680 16356 116686
rect 16304 116622 16356 116628
rect 16120 116272 16172 116278
rect 16120 116214 16172 116220
rect 16408 116226 16436 119200
rect 16592 117434 16620 119200
rect 16580 117428 16632 117434
rect 16580 117370 16632 117376
rect 16580 117156 16632 117162
rect 16580 117098 16632 117104
rect 16408 116198 16528 116226
rect 15936 116136 15988 116142
rect 15936 116078 15988 116084
rect 16396 116068 16448 116074
rect 16396 116010 16448 116016
rect 15844 115796 15896 115802
rect 15844 115738 15896 115744
rect 16408 115258 16436 116010
rect 16396 115252 16448 115258
rect 16396 115194 16448 115200
rect 16500 113966 16528 116198
rect 16592 115734 16620 117098
rect 16776 116890 16804 119200
rect 16764 116884 16816 116890
rect 16764 116826 16816 116832
rect 16580 115728 16632 115734
rect 16580 115670 16632 115676
rect 17052 114578 17080 119200
rect 17236 116686 17264 119200
rect 17420 117586 17448 119200
rect 17420 117558 17632 117586
rect 17604 116890 17632 117558
rect 17592 116884 17644 116890
rect 17592 116826 17644 116832
rect 17408 116748 17460 116754
rect 17408 116690 17460 116696
rect 17224 116680 17276 116686
rect 17224 116622 17276 116628
rect 17420 115666 17448 116690
rect 17408 115660 17460 115666
rect 17408 115602 17460 115608
rect 17316 114980 17368 114986
rect 17316 114922 17368 114928
rect 17328 114714 17356 114922
rect 17316 114708 17368 114714
rect 17316 114650 17368 114656
rect 17040 114572 17092 114578
rect 17040 114514 17092 114520
rect 17696 113966 17724 119200
rect 17776 117224 17828 117230
rect 17776 117166 17828 117172
rect 17880 117178 17908 119200
rect 17788 115598 17816 117166
rect 17880 117150 18000 117178
rect 17868 117088 17920 117094
rect 17868 117030 17920 117036
rect 17880 116822 17908 117030
rect 17868 116816 17920 116822
rect 17868 116758 17920 116764
rect 17972 116618 18000 117150
rect 18064 116822 18092 119200
rect 18052 116816 18104 116822
rect 18052 116758 18104 116764
rect 18144 116748 18196 116754
rect 18144 116690 18196 116696
rect 17960 116612 18012 116618
rect 17960 116554 18012 116560
rect 17776 115592 17828 115598
rect 17776 115534 17828 115540
rect 18156 115258 18184 116690
rect 18144 115252 18196 115258
rect 18144 115194 18196 115200
rect 18052 114572 18104 114578
rect 18052 114514 18104 114520
rect 18064 114170 18092 114514
rect 18052 114164 18104 114170
rect 18052 114106 18104 114112
rect 18248 113966 18276 119200
rect 18524 117638 18552 119200
rect 18512 117632 18564 117638
rect 18512 117574 18564 117580
rect 18708 116890 18736 119200
rect 18696 116884 18748 116890
rect 18892 116872 18920 119200
rect 19064 117632 19116 117638
rect 19064 117574 19116 117580
rect 19076 117366 19104 117574
rect 19064 117360 19116 117366
rect 19064 117302 19116 117308
rect 19064 117156 19116 117162
rect 19064 117098 19116 117104
rect 18892 116844 19012 116872
rect 18696 116826 18748 116832
rect 18880 116748 18932 116754
rect 18880 116690 18932 116696
rect 18696 115184 18748 115190
rect 18696 115126 18748 115132
rect 18708 114578 18736 115126
rect 18892 115122 18920 116690
rect 18880 115116 18932 115122
rect 18880 115058 18932 115064
rect 18880 114912 18932 114918
rect 18880 114854 18932 114860
rect 18696 114572 18748 114578
rect 18696 114514 18748 114520
rect 18892 114442 18920 114854
rect 18984 114578 19012 116844
rect 19076 116686 19104 117098
rect 19168 116822 19196 119200
rect 19352 117230 19380 119200
rect 19340 117224 19392 117230
rect 19340 117166 19392 117172
rect 19536 117076 19564 119200
rect 19812 117434 19840 119200
rect 19800 117428 19852 117434
rect 19800 117370 19852 117376
rect 19892 117360 19944 117366
rect 19890 117328 19892 117337
rect 19944 117328 19946 117337
rect 19890 117263 19946 117272
rect 19892 117156 19944 117162
rect 19892 117098 19944 117104
rect 19444 117048 19564 117076
rect 19156 116816 19208 116822
rect 19156 116758 19208 116764
rect 19340 116748 19392 116754
rect 19340 116690 19392 116696
rect 19064 116680 19116 116686
rect 19064 116622 19116 116628
rect 19352 115258 19380 116690
rect 19340 115252 19392 115258
rect 19340 115194 19392 115200
rect 19340 115116 19392 115122
rect 19340 115058 19392 115064
rect 18972 114572 19024 114578
rect 18972 114514 19024 114520
rect 19352 114442 19380 115058
rect 19444 114646 19472 117048
rect 19580 116988 19876 117008
rect 19636 116986 19660 116988
rect 19716 116986 19740 116988
rect 19796 116986 19820 116988
rect 19658 116934 19660 116986
rect 19722 116934 19734 116986
rect 19796 116934 19798 116986
rect 19636 116932 19660 116934
rect 19716 116932 19740 116934
rect 19796 116932 19820 116934
rect 19580 116912 19876 116932
rect 19904 116210 19932 117098
rect 19996 116346 20024 119200
rect 20076 116680 20128 116686
rect 20076 116622 20128 116628
rect 19984 116340 20036 116346
rect 19984 116282 20036 116288
rect 19892 116204 19944 116210
rect 19892 116146 19944 116152
rect 19580 115900 19876 115920
rect 19636 115898 19660 115900
rect 19716 115898 19740 115900
rect 19796 115898 19820 115900
rect 19658 115846 19660 115898
rect 19722 115846 19734 115898
rect 19796 115846 19798 115898
rect 19636 115844 19660 115846
rect 19716 115844 19740 115846
rect 19796 115844 19820 115846
rect 19580 115824 19876 115844
rect 20088 115802 20116 116622
rect 20076 115796 20128 115802
rect 20076 115738 20128 115744
rect 19580 114812 19876 114832
rect 19636 114810 19660 114812
rect 19716 114810 19740 114812
rect 19796 114810 19820 114812
rect 19658 114758 19660 114810
rect 19722 114758 19734 114810
rect 19796 114758 19798 114810
rect 19636 114756 19660 114758
rect 19716 114756 19740 114758
rect 19796 114756 19820 114758
rect 19580 114736 19876 114756
rect 19432 114640 19484 114646
rect 19432 114582 19484 114588
rect 18880 114436 18932 114442
rect 18880 114378 18932 114384
rect 19340 114436 19392 114442
rect 19340 114378 19392 114384
rect 20180 113966 20208 119200
rect 20364 117706 20392 119200
rect 20352 117700 20404 117706
rect 20352 117642 20404 117648
rect 20260 117428 20312 117434
rect 20260 117370 20312 117376
rect 20272 115841 20300 117370
rect 20444 117224 20496 117230
rect 20444 117166 20496 117172
rect 20456 116890 20484 117166
rect 20536 117156 20588 117162
rect 20536 117098 20588 117104
rect 20444 116884 20496 116890
rect 20444 116826 20496 116832
rect 20352 116748 20404 116754
rect 20352 116690 20404 116696
rect 20258 115832 20314 115841
rect 20258 115767 20314 115776
rect 20364 115258 20392 116690
rect 20548 116074 20576 117098
rect 20640 116872 20668 119200
rect 20720 116884 20772 116890
rect 20640 116844 20720 116872
rect 20720 116826 20772 116832
rect 20536 116068 20588 116074
rect 20536 116010 20588 116016
rect 20720 116000 20772 116006
rect 20720 115942 20772 115948
rect 20732 115258 20760 115942
rect 20352 115252 20404 115258
rect 20352 115194 20404 115200
rect 20720 115252 20772 115258
rect 20720 115194 20772 115200
rect 20720 114708 20772 114714
rect 20720 114650 20772 114656
rect 20732 114617 20760 114650
rect 20718 114608 20774 114617
rect 20260 114572 20312 114578
rect 20718 114543 20774 114552
rect 20260 114514 20312 114520
rect 20272 114170 20300 114514
rect 20720 114504 20772 114510
rect 20720 114446 20772 114452
rect 20260 114164 20312 114170
rect 20260 114106 20312 114112
rect 20732 114034 20760 114446
rect 20720 114028 20772 114034
rect 20720 113970 20772 113976
rect 20824 113966 20852 119200
rect 21008 117434 21036 119200
rect 20996 117428 21048 117434
rect 20996 117370 21048 117376
rect 21088 116544 21140 116550
rect 21088 116486 21140 116492
rect 21100 115666 21128 116486
rect 21284 116346 21312 119200
rect 21364 117156 21416 117162
rect 21364 117098 21416 117104
rect 21272 116340 21324 116346
rect 21272 116282 21324 116288
rect 21376 116278 21404 117098
rect 21468 116906 21496 119200
rect 21652 117638 21680 119200
rect 21640 117632 21692 117638
rect 21640 117574 21692 117580
rect 21640 117224 21692 117230
rect 21640 117166 21692 117172
rect 21468 116878 21588 116906
rect 21454 116648 21510 116657
rect 21454 116583 21510 116592
rect 21364 116272 21416 116278
rect 21364 116214 21416 116220
rect 21088 115660 21140 115666
rect 21088 115602 21140 115608
rect 20902 115288 20958 115297
rect 20902 115223 20958 115232
rect 20916 114918 20944 115223
rect 20904 114912 20956 114918
rect 20904 114854 20956 114860
rect 20996 114912 21048 114918
rect 20996 114854 21048 114860
rect 20904 114572 20956 114578
rect 21008 114560 21036 114854
rect 21468 114730 21496 116583
rect 21376 114714 21496 114730
rect 21364 114708 21496 114714
rect 21416 114702 21496 114708
rect 21364 114650 21416 114656
rect 21560 114594 21588 116878
rect 21652 115666 21680 117166
rect 21732 117088 21784 117094
rect 21732 117030 21784 117036
rect 21744 116618 21772 117030
rect 21732 116612 21784 116618
rect 21732 116554 21784 116560
rect 21824 116612 21876 116618
rect 21824 116554 21876 116560
rect 21836 115934 21864 116554
rect 21928 116362 21956 119200
rect 22008 117224 22060 117230
rect 22008 117166 22060 117172
rect 22112 117178 22140 119200
rect 22020 116686 22048 117166
rect 22112 117150 22232 117178
rect 22204 116770 22232 117150
rect 22296 116890 22324 119200
rect 22376 117428 22428 117434
rect 22376 117370 22428 117376
rect 22284 116884 22336 116890
rect 22284 116826 22336 116832
rect 22388 116822 22416 117370
rect 22376 116816 22428 116822
rect 22204 116742 22324 116770
rect 22376 116758 22428 116764
rect 22008 116680 22060 116686
rect 22100 116680 22152 116686
rect 22008 116622 22060 116628
rect 22098 116648 22100 116657
rect 22152 116648 22154 116657
rect 22098 116583 22154 116592
rect 21928 116346 22140 116362
rect 21928 116340 22152 116346
rect 21928 116334 22100 116340
rect 22100 116282 22152 116288
rect 21914 116240 21970 116249
rect 21914 116175 21970 116184
rect 21744 115906 21864 115934
rect 21640 115660 21692 115666
rect 21640 115602 21692 115608
rect 21640 115524 21692 115530
rect 21640 115466 21692 115472
rect 21652 115258 21680 115466
rect 21640 115252 21692 115258
rect 21640 115194 21692 115200
rect 21744 114714 21772 115906
rect 21732 114708 21784 114714
rect 21732 114650 21784 114656
rect 21824 114640 21876 114646
rect 21560 114588 21824 114594
rect 21560 114582 21876 114588
rect 21560 114566 21864 114582
rect 20956 114532 21036 114560
rect 20904 114514 20956 114520
rect 15752 113960 15804 113966
rect 15752 113902 15804 113908
rect 16488 113960 16540 113966
rect 16488 113902 16540 113908
rect 17684 113960 17736 113966
rect 17684 113902 17736 113908
rect 18236 113960 18288 113966
rect 18236 113902 18288 113908
rect 20168 113960 20220 113966
rect 20168 113902 20220 113908
rect 20812 113960 20864 113966
rect 20812 113902 20864 113908
rect 19580 113724 19876 113744
rect 19636 113722 19660 113724
rect 19716 113722 19740 113724
rect 19796 113722 19820 113724
rect 19658 113670 19660 113722
rect 19722 113670 19734 113722
rect 19796 113670 19798 113722
rect 19636 113668 19660 113670
rect 19716 113668 19740 113670
rect 19796 113668 19820 113670
rect 19580 113648 19876 113668
rect 14648 113552 14700 113558
rect 14648 113494 14700 113500
rect 13360 113416 13412 113422
rect 13360 113358 13412 113364
rect 21640 113416 21692 113422
rect 21640 113358 21692 113364
rect 16028 112736 16080 112742
rect 16028 112678 16080 112684
rect 12716 112396 12768 112402
rect 12716 112338 12768 112344
rect 11060 109540 11112 109546
rect 11060 109482 11112 109488
rect 8668 109268 8720 109274
rect 8668 109210 8720 109216
rect 8944 105120 8996 105126
rect 8944 105062 8996 105068
rect 8956 85270 8984 105062
rect 10324 104576 10376 104582
rect 10324 104518 10376 104524
rect 9036 103556 9088 103562
rect 9036 103498 9088 103504
rect 9048 87446 9076 103498
rect 9128 98116 9180 98122
rect 9128 98058 9180 98064
rect 9140 88602 9168 98058
rect 9220 88868 9272 88874
rect 9220 88810 9272 88816
rect 9128 88596 9180 88602
rect 9128 88538 9180 88544
rect 9036 87440 9088 87446
rect 9036 87382 9088 87388
rect 8944 85264 8996 85270
rect 8944 85206 8996 85212
rect 9232 84182 9260 88810
rect 10336 85610 10364 104518
rect 11072 103834 11100 109482
rect 11060 103828 11112 103834
rect 11060 103770 11112 103776
rect 12532 103692 12584 103698
rect 12532 103634 12584 103640
rect 12624 103692 12676 103698
rect 12624 103634 12676 103640
rect 12440 102740 12492 102746
rect 12440 102682 12492 102688
rect 12072 102536 12124 102542
rect 12072 102478 12124 102484
rect 12084 101998 12112 102478
rect 12072 101992 12124 101998
rect 12072 101934 12124 101940
rect 12256 101924 12308 101930
rect 12256 101866 12308 101872
rect 12268 101538 12296 101866
rect 12452 101862 12480 102682
rect 12544 102542 12572 103634
rect 12636 102678 12664 103634
rect 12624 102672 12676 102678
rect 12624 102614 12676 102620
rect 12532 102536 12584 102542
rect 12532 102478 12584 102484
rect 12440 101856 12492 101862
rect 12440 101798 12492 101804
rect 12452 101658 12480 101798
rect 12440 101652 12492 101658
rect 12440 101594 12492 101600
rect 12544 101538 12572 102478
rect 12624 102060 12676 102066
rect 12624 102002 12676 102008
rect 12636 101862 12664 102002
rect 12624 101856 12676 101862
rect 12624 101798 12676 101804
rect 12636 101590 12664 101798
rect 12728 101658 12756 112338
rect 13084 109132 13136 109138
rect 13084 109074 13136 109080
rect 12716 101652 12768 101658
rect 12716 101594 12768 101600
rect 12268 101510 12572 101538
rect 12624 101584 12676 101590
rect 12624 101526 12676 101532
rect 12544 101454 12572 101510
rect 12900 101516 12952 101522
rect 12900 101458 12952 101464
rect 10876 101448 10928 101454
rect 10876 101390 10928 101396
rect 12532 101448 12584 101454
rect 12532 101390 12584 101396
rect 10888 91866 10916 101390
rect 12072 100020 12124 100026
rect 12072 99962 12124 99968
rect 11704 96960 11756 96966
rect 11704 96902 11756 96908
rect 10876 91860 10928 91866
rect 10876 91802 10928 91808
rect 10784 91724 10836 91730
rect 10784 91666 10836 91672
rect 10324 85604 10376 85610
rect 10324 85546 10376 85552
rect 9220 84176 9272 84182
rect 9220 84118 9272 84124
rect 8852 82952 8904 82958
rect 8852 82894 8904 82900
rect 8864 79898 8892 82894
rect 8852 79892 8904 79898
rect 8852 79834 8904 79840
rect 8300 76288 8352 76294
rect 8300 76230 8352 76236
rect 8312 73234 8340 76230
rect 9680 75744 9732 75750
rect 9680 75686 9732 75692
rect 9220 74724 9272 74730
rect 9220 74666 9272 74672
rect 8944 74180 8996 74186
rect 8944 74122 8996 74128
rect 8300 73228 8352 73234
rect 8300 73170 8352 73176
rect 8956 62898 8984 74122
rect 9036 68196 9088 68202
rect 9036 68138 9088 68144
rect 8944 62892 8996 62898
rect 8944 62834 8996 62840
rect 8024 62824 8076 62830
rect 8024 62766 8076 62772
rect 7840 62144 7892 62150
rect 7840 62086 7892 62092
rect 7852 52562 7880 62086
rect 8484 61600 8536 61606
rect 8484 61542 8536 61548
rect 8300 56976 8352 56982
rect 8300 56918 8352 56924
rect 7932 53440 7984 53446
rect 7932 53382 7984 53388
rect 7840 52556 7892 52562
rect 7840 52498 7892 52504
rect 7656 49700 7708 49706
rect 7656 49642 7708 49648
rect 7748 49700 7800 49706
rect 7748 49642 7800 49648
rect 7564 47116 7616 47122
rect 7564 47058 7616 47064
rect 7472 47048 7524 47054
rect 7472 46990 7524 46996
rect 7840 46980 7892 46986
rect 7840 46922 7892 46928
rect 7748 46504 7800 46510
rect 7748 46446 7800 46452
rect 7760 45966 7788 46446
rect 7748 45960 7800 45966
rect 7748 45902 7800 45908
rect 7760 45626 7788 45902
rect 7748 45620 7800 45626
rect 7748 45562 7800 45568
rect 7380 45484 7432 45490
rect 7380 45426 7432 45432
rect 7288 45416 7340 45422
rect 7288 45358 7340 45364
rect 7300 43790 7328 45358
rect 7392 44334 7420 45426
rect 7380 44328 7432 44334
rect 7380 44270 7432 44276
rect 7748 44192 7800 44198
rect 7748 44134 7800 44140
rect 7288 43784 7340 43790
rect 7288 43726 7340 43732
rect 7196 42152 7248 42158
rect 7196 42094 7248 42100
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 7116 16574 7144 36722
rect 7484 17882 7512 40870
rect 7564 22500 7616 22506
rect 7564 22442 7616 22448
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7116 16546 7236 16574
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 3670 6960 8910
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6196 800 6224 2450
rect 6472 800 6500 2926
rect 6840 800 6868 3334
rect 7116 800 7144 4014
rect 7208 2582 7236 16546
rect 7576 14618 7604 22442
rect 7760 20058 7788 44134
rect 7852 35766 7880 46922
rect 7944 45554 7972 53382
rect 8024 52964 8076 52970
rect 8024 52906 8076 52912
rect 8036 49366 8064 52906
rect 8312 52086 8340 56918
rect 8392 56160 8444 56166
rect 8392 56102 8444 56108
rect 8300 52080 8352 52086
rect 8300 52022 8352 52028
rect 8300 51060 8352 51066
rect 8300 51002 8352 51008
rect 8024 49360 8076 49366
rect 8024 49302 8076 49308
rect 8208 49156 8260 49162
rect 8208 49098 8260 49104
rect 8220 47530 8248 49098
rect 8208 47524 8260 47530
rect 8208 47466 8260 47472
rect 8312 47122 8340 51002
rect 8404 49910 8432 56102
rect 8392 49904 8444 49910
rect 8392 49846 8444 49852
rect 8392 49700 8444 49706
rect 8392 49642 8444 49648
rect 8404 47598 8432 49642
rect 8392 47592 8444 47598
rect 8392 47534 8444 47540
rect 8392 47252 8444 47258
rect 8392 47194 8444 47200
rect 8300 47116 8352 47122
rect 8300 47058 8352 47064
rect 8404 46510 8432 47194
rect 8392 46504 8444 46510
rect 8392 46446 8444 46452
rect 7944 45526 8064 45554
rect 7932 42152 7984 42158
rect 7932 42094 7984 42100
rect 7944 41614 7972 42094
rect 7932 41608 7984 41614
rect 7932 41550 7984 41556
rect 7944 41070 7972 41550
rect 7932 41064 7984 41070
rect 7932 41006 7984 41012
rect 7944 40526 7972 41006
rect 7932 40520 7984 40526
rect 7932 40462 7984 40468
rect 7932 40384 7984 40390
rect 7932 40326 7984 40332
rect 7944 39982 7972 40326
rect 8036 40050 8064 45526
rect 8116 44736 8168 44742
rect 8116 44678 8168 44684
rect 8128 40474 8156 44678
rect 8208 44328 8260 44334
rect 8208 44270 8260 44276
rect 8220 43858 8248 44270
rect 8496 43858 8524 61542
rect 8944 59968 8996 59974
rect 8944 59910 8996 59916
rect 8760 52556 8812 52562
rect 8760 52498 8812 52504
rect 8576 46368 8628 46374
rect 8576 46310 8628 46316
rect 8208 43852 8260 43858
rect 8208 43794 8260 43800
rect 8484 43852 8536 43858
rect 8484 43794 8536 43800
rect 8588 43738 8616 46310
rect 8668 45280 8720 45286
rect 8668 45222 8720 45228
rect 8208 43716 8260 43722
rect 8208 43658 8260 43664
rect 8496 43710 8616 43738
rect 8220 41138 8248 43658
rect 8496 42906 8524 43710
rect 8576 43648 8628 43654
rect 8576 43590 8628 43596
rect 8484 42900 8536 42906
rect 8484 42842 8536 42848
rect 8588 42090 8616 43590
rect 8576 42084 8628 42090
rect 8576 42026 8628 42032
rect 8300 41472 8352 41478
rect 8300 41414 8352 41420
rect 8208 41132 8260 41138
rect 8208 41074 8260 41080
rect 8220 40594 8248 41074
rect 8208 40588 8260 40594
rect 8208 40530 8260 40536
rect 8128 40446 8248 40474
rect 8116 40384 8168 40390
rect 8116 40326 8168 40332
rect 8024 40044 8076 40050
rect 8024 39986 8076 39992
rect 7932 39976 7984 39982
rect 7932 39918 7984 39924
rect 7840 35760 7892 35766
rect 7840 35702 7892 35708
rect 7840 33924 7892 33930
rect 7840 33866 7892 33872
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7392 800 7420 3538
rect 7852 3194 7880 33866
rect 8128 27538 8156 40326
rect 8220 39506 8248 40446
rect 8208 39500 8260 39506
rect 8208 39442 8260 39448
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 3040 7972 26386
rect 8312 17270 8340 41414
rect 8576 40452 8628 40458
rect 8576 40394 8628 40400
rect 8392 39840 8444 39846
rect 8392 39782 8444 39788
rect 8404 35562 8432 39782
rect 8392 35556 8444 35562
rect 8392 35498 8444 35504
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8220 11014 8248 15642
rect 8404 15026 8432 17818
rect 8588 16574 8616 40394
rect 8680 19174 8708 45222
rect 8772 44334 8800 52498
rect 8956 49706 8984 59910
rect 9048 57934 9076 68138
rect 9128 65136 9180 65142
rect 9128 65078 9180 65084
rect 9036 57928 9088 57934
rect 9036 57870 9088 57876
rect 9140 56506 9168 65078
rect 9128 56500 9180 56506
rect 9128 56442 9180 56448
rect 8944 49700 8996 49706
rect 8944 49642 8996 49648
rect 9232 47122 9260 74666
rect 9496 63232 9548 63238
rect 9496 63174 9548 63180
rect 9220 47116 9272 47122
rect 9220 47058 9272 47064
rect 9036 47048 9088 47054
rect 9036 46990 9088 46996
rect 9048 46442 9076 46990
rect 9220 46980 9272 46986
rect 9220 46922 9272 46928
rect 9036 46436 9088 46442
rect 9036 46378 9088 46384
rect 9036 44736 9088 44742
rect 9036 44678 9088 44684
rect 8760 44328 8812 44334
rect 8760 44270 8812 44276
rect 9048 42838 9076 44678
rect 9036 42832 9088 42838
rect 9036 42774 9088 42780
rect 9128 41472 9180 41478
rect 9128 41414 9180 41420
rect 8760 36576 8812 36582
rect 8760 36518 8812 36524
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8588 16546 8708 16574
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7852 3012 7972 3040
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7668 800 7696 2926
rect 7852 2378 7880 3012
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7932 2916 7984 2922
rect 7932 2858 7984 2864
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 7944 800 7972 2858
rect 8220 800 8248 2926
rect 8588 800 8616 3538
rect 8680 2650 8708 16546
rect 8772 3738 8800 36518
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 4486 8984 19178
rect 9140 17542 9168 41414
rect 9232 39370 9260 46922
rect 9404 46912 9456 46918
rect 9404 46854 9456 46860
rect 9416 46578 9444 46854
rect 9404 46572 9456 46578
rect 9404 46514 9456 46520
rect 9312 45824 9364 45830
rect 9312 45766 9364 45772
rect 9220 39364 9272 39370
rect 9220 39306 9272 39312
rect 9324 31142 9352 45766
rect 9508 45554 9536 63174
rect 9692 46510 9720 75686
rect 10048 62892 10100 62898
rect 10048 62834 10100 62840
rect 9772 56500 9824 56506
rect 9772 56442 9824 56448
rect 9784 47598 9812 56442
rect 9956 53100 10008 53106
rect 9956 53042 10008 53048
rect 9772 47592 9824 47598
rect 9772 47534 9824 47540
rect 9680 46504 9732 46510
rect 9680 46446 9732 46452
rect 9864 46368 9916 46374
rect 9864 46310 9916 46316
rect 9416 45526 9536 45554
rect 9416 45422 9444 45526
rect 9404 45416 9456 45422
rect 9404 45358 9456 45364
rect 9496 45416 9548 45422
rect 9496 45358 9548 45364
rect 9508 44878 9536 45358
rect 9496 44872 9548 44878
rect 9496 44814 9548 44820
rect 9508 43994 9536 44814
rect 9876 44402 9904 46310
rect 9968 45422 9996 53042
rect 10060 47122 10088 62834
rect 10508 57928 10560 57934
rect 10508 57870 10560 57876
rect 10140 49700 10192 49706
rect 10140 49642 10192 49648
rect 10048 47116 10100 47122
rect 10048 47058 10100 47064
rect 9956 45416 10008 45422
rect 9956 45358 10008 45364
rect 9864 44396 9916 44402
rect 9864 44338 9916 44344
rect 10152 44334 10180 49642
rect 10232 47456 10284 47462
rect 10232 47398 10284 47404
rect 10140 44328 10192 44334
rect 10140 44270 10192 44276
rect 9864 44192 9916 44198
rect 9864 44134 9916 44140
rect 9496 43988 9548 43994
rect 9496 43930 9548 43936
rect 9588 43920 9640 43926
rect 9588 43862 9640 43868
rect 9496 41744 9548 41750
rect 9496 41686 9548 41692
rect 9508 39438 9536 41686
rect 9600 41070 9628 43862
rect 9588 41064 9640 41070
rect 9588 41006 9640 41012
rect 9876 40050 9904 44134
rect 9956 40928 10008 40934
rect 9956 40870 10008 40876
rect 9864 40044 9916 40050
rect 9864 39986 9916 39992
rect 9496 39432 9548 39438
rect 9496 39374 9548 39380
rect 9312 31136 9364 31142
rect 9312 31078 9364 31084
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9416 16726 9444 25094
rect 9968 23118 9996 40870
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 9404 16720 9456 16726
rect 9404 16662 9456 16668
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8864 800 8892 3334
rect 8956 3194 8984 3946
rect 9416 3670 9444 10406
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 9140 800 9168 2450
rect 9416 800 9444 2926
rect 9600 2922 9628 4762
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 9692 800 9720 3334
rect 10152 2582 10180 33254
rect 10244 27606 10272 47398
rect 10520 44946 10548 57870
rect 10508 44940 10560 44946
rect 10508 44882 10560 44888
rect 10692 44736 10744 44742
rect 10692 44678 10744 44684
rect 10324 42084 10376 42090
rect 10324 42026 10376 42032
rect 10232 27600 10284 27606
rect 10232 27542 10284 27548
rect 10336 18873 10364 42026
rect 10704 34542 10732 44678
rect 10692 34536 10744 34542
rect 10692 34478 10744 34484
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10322 18864 10378 18873
rect 10322 18799 10378 18808
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 3670 10272 11834
rect 10428 3942 10456 13262
rect 10520 11762 10548 23802
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10612 11082 10640 21558
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10796 8430 10824 91666
rect 11716 87922 11744 96902
rect 11704 87916 11756 87922
rect 11704 87858 11756 87864
rect 11980 59016 12032 59022
rect 11980 58958 12032 58964
rect 11992 58410 12020 58958
rect 11980 58404 12032 58410
rect 11980 58346 12032 58352
rect 11992 58002 12020 58346
rect 11980 57996 12032 58002
rect 11980 57938 12032 57944
rect 11060 51332 11112 51338
rect 11060 51274 11112 51280
rect 10968 40996 11020 41002
rect 10968 40938 11020 40944
rect 10980 39574 11008 40938
rect 10968 39568 11020 39574
rect 10968 39510 11020 39516
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 4078 11008 7754
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10140 2576 10192 2582
rect 10140 2518 10192 2524
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 9968 800 9996 2450
rect 10336 800 10364 2450
rect 10612 800 10640 3878
rect 11072 3738 11100 51274
rect 11152 44940 11204 44946
rect 11152 44882 11204 44888
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10888 800 10916 2926
rect 11072 1850 11100 3538
rect 11164 3194 11192 44882
rect 11888 44804 11940 44810
rect 11888 44746 11940 44752
rect 11704 40044 11756 40050
rect 11704 39986 11756 39992
rect 11716 17746 11744 39986
rect 11900 34542 11928 44746
rect 11796 34536 11848 34542
rect 11796 34478 11848 34484
rect 11888 34536 11940 34542
rect 11888 34478 11940 34484
rect 11808 24750 11836 34478
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 12084 6914 12112 99962
rect 12544 97510 12572 101390
rect 12912 99278 12940 101458
rect 12900 99272 12952 99278
rect 12900 99214 12952 99220
rect 12532 97504 12584 97510
rect 12532 97446 12584 97452
rect 12256 77376 12308 77382
rect 12256 77318 12308 77324
rect 12164 73228 12216 73234
rect 12164 73170 12216 73176
rect 12176 58002 12204 73170
rect 12268 59090 12296 77318
rect 12992 65544 13044 65550
rect 12992 65486 13044 65492
rect 12256 59084 12308 59090
rect 12256 59026 12308 59032
rect 13004 58478 13032 65486
rect 12992 58472 13044 58478
rect 12992 58414 13044 58420
rect 12348 58336 12400 58342
rect 12348 58278 12400 58284
rect 12164 57996 12216 58002
rect 12164 57938 12216 57944
rect 12256 50380 12308 50386
rect 12256 50322 12308 50328
rect 11992 6886 12112 6914
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4078 11744 4966
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11072 1822 11192 1850
rect 11164 800 11192 1822
rect 11440 800 11468 3878
rect 11992 3058 12020 6886
rect 12268 3738 12296 50322
rect 12360 39370 12388 58278
rect 12440 57996 12492 58002
rect 12440 57938 12492 57944
rect 12452 45558 12480 57938
rect 12440 45552 12492 45558
rect 12440 45494 12492 45500
rect 12348 39364 12400 39370
rect 12348 39306 12400 39312
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12360 7886 12388 15574
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11808 800 11836 2926
rect 12084 800 12112 3538
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12360 800 12388 3334
rect 12452 2582 12480 5034
rect 12912 3670 12940 11018
rect 13096 6866 13124 109074
rect 13452 108044 13504 108050
rect 13452 107986 13504 107992
rect 13176 102604 13228 102610
rect 13176 102546 13228 102552
rect 13188 99278 13216 102546
rect 13360 102400 13412 102406
rect 13360 102342 13412 102348
rect 13176 99272 13228 99278
rect 13176 99214 13228 99220
rect 13188 90778 13216 99214
rect 13176 90772 13228 90778
rect 13176 90714 13228 90720
rect 13268 47524 13320 47530
rect 13268 47466 13320 47472
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 19922 13216 23054
rect 13280 22574 13308 47466
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13280 9382 13308 18362
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13372 5574 13400 102342
rect 13464 102134 13492 107986
rect 14464 103692 14516 103698
rect 14464 103634 14516 103640
rect 13544 103488 13596 103494
rect 13544 103430 13596 103436
rect 13556 102746 13584 103430
rect 13544 102740 13596 102746
rect 13544 102682 13596 102688
rect 13452 102128 13504 102134
rect 13452 102070 13504 102076
rect 13556 102066 13584 102682
rect 13544 102060 13596 102066
rect 13544 102002 13596 102008
rect 13728 99408 13780 99414
rect 13728 99350 13780 99356
rect 13452 44260 13504 44266
rect 13452 44202 13504 44208
rect 13464 20466 13492 44202
rect 13544 40384 13596 40390
rect 13544 40326 13596 40332
rect 13556 23322 13584 40326
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13452 19168 13504 19174
rect 13450 19136 13452 19145
rect 13504 19136 13506 19145
rect 13450 19071 13506 19080
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13464 8362 13492 16730
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13740 3058 13768 99350
rect 13820 98728 13872 98734
rect 13820 98670 13872 98676
rect 13832 7562 13860 98670
rect 14004 97300 14056 97306
rect 14004 97242 14056 97248
rect 13832 7534 13952 7562
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12636 800 12664 2450
rect 12912 800 12940 2926
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13188 800 13216 2790
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13556 800 13584 2450
rect 13832 800 13860 3538
rect 13924 2582 13952 7534
rect 14016 3670 14044 97242
rect 14476 33318 14504 103634
rect 15200 103012 15252 103018
rect 15200 102954 15252 102960
rect 15212 99414 15240 102954
rect 15936 100428 15988 100434
rect 15936 100370 15988 100376
rect 15200 99408 15252 99414
rect 15200 99350 15252 99356
rect 15200 99272 15252 99278
rect 15200 99214 15252 99220
rect 15212 97578 15240 99214
rect 15200 97572 15252 97578
rect 15200 97514 15252 97520
rect 15844 97572 15896 97578
rect 15844 97514 15896 97520
rect 15108 97504 15160 97510
rect 15108 97446 15160 97452
rect 15120 95470 15148 97446
rect 15108 95464 15160 95470
rect 15108 95406 15160 95412
rect 15856 91866 15884 97514
rect 15844 91860 15896 91866
rect 15844 91802 15896 91808
rect 15292 71052 15344 71058
rect 15292 70994 15344 71000
rect 15304 64122 15332 70994
rect 15292 64116 15344 64122
rect 15292 64058 15344 64064
rect 15200 63844 15252 63850
rect 15200 63786 15252 63792
rect 14648 48000 14700 48006
rect 14648 47942 14700 47948
rect 14556 42016 14608 42022
rect 14556 41958 14608 41964
rect 14464 33312 14516 33318
rect 14464 33254 14516 33260
rect 14462 28792 14518 28801
rect 14462 28727 14518 28736
rect 14476 21418 14504 28727
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14464 18896 14516 18902
rect 14464 18838 14516 18844
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14384 13190 14412 17274
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14476 6322 14504 18838
rect 14568 14958 14596 41958
rect 14660 22234 14688 47942
rect 15108 47048 15160 47054
rect 15108 46990 15160 46996
rect 15120 46646 15148 46990
rect 15108 46640 15160 46646
rect 15108 46582 15160 46588
rect 15108 44532 15160 44538
rect 15108 44474 15160 44480
rect 14740 42832 14792 42838
rect 14740 42774 14792 42780
rect 14752 25838 14780 42774
rect 15120 41614 15148 44474
rect 15108 41608 15160 41614
rect 15108 41550 15160 41556
rect 14832 35760 14884 35766
rect 14832 35702 14884 35708
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14844 21486 14872 35702
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14936 15570 14964 27474
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 14108 800 14136 3334
rect 14568 2922 14596 3606
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14384 800 14412 2450
rect 14660 800 14688 4626
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14752 2990 14780 4082
rect 14844 3602 14872 10542
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14832 2916 14884 2922
rect 14936 2904 14964 6258
rect 15028 4078 15056 7822
rect 15212 6798 15240 63786
rect 15844 45280 15896 45286
rect 15844 45222 15896 45228
rect 15752 35556 15804 35562
rect 15752 35498 15804 35504
rect 15292 31952 15344 31958
rect 15292 31894 15344 31900
rect 15304 29646 15332 31894
rect 15292 29640 15344 29646
rect 15292 29582 15344 29588
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15304 21010 15332 27542
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15764 18834 15792 35498
rect 15856 24818 15884 45222
rect 15948 36786 15976 100370
rect 16040 91866 16068 112678
rect 19580 112636 19876 112656
rect 19636 112634 19660 112636
rect 19716 112634 19740 112636
rect 19796 112634 19820 112636
rect 19658 112582 19660 112634
rect 19722 112582 19734 112634
rect 19796 112582 19798 112634
rect 19636 112580 19660 112582
rect 19716 112580 19740 112582
rect 19796 112580 19820 112582
rect 19580 112560 19876 112580
rect 20720 112464 20772 112470
rect 20720 112406 20772 112412
rect 19580 111548 19876 111568
rect 19636 111546 19660 111548
rect 19716 111546 19740 111548
rect 19796 111546 19820 111548
rect 19658 111494 19660 111546
rect 19722 111494 19734 111546
rect 19796 111494 19798 111546
rect 19636 111492 19660 111494
rect 19716 111492 19740 111494
rect 19796 111492 19820 111494
rect 19580 111472 19876 111492
rect 19580 110460 19876 110480
rect 19636 110458 19660 110460
rect 19716 110458 19740 110460
rect 19796 110458 19820 110460
rect 19658 110406 19660 110458
rect 19722 110406 19734 110458
rect 19796 110406 19798 110458
rect 19636 110404 19660 110406
rect 19716 110404 19740 110406
rect 19796 110404 19820 110406
rect 19580 110384 19876 110404
rect 19580 109372 19876 109392
rect 19636 109370 19660 109372
rect 19716 109370 19740 109372
rect 19796 109370 19820 109372
rect 19658 109318 19660 109370
rect 19722 109318 19734 109370
rect 19796 109318 19798 109370
rect 19636 109316 19660 109318
rect 19716 109316 19740 109318
rect 19796 109316 19820 109318
rect 19580 109296 19876 109316
rect 19580 108284 19876 108304
rect 19636 108282 19660 108284
rect 19716 108282 19740 108284
rect 19796 108282 19820 108284
rect 19658 108230 19660 108282
rect 19722 108230 19734 108282
rect 19796 108230 19798 108282
rect 19636 108228 19660 108230
rect 19716 108228 19740 108230
rect 19796 108228 19820 108230
rect 19580 108208 19876 108228
rect 19580 107196 19876 107216
rect 19636 107194 19660 107196
rect 19716 107194 19740 107196
rect 19796 107194 19820 107196
rect 19658 107142 19660 107194
rect 19722 107142 19734 107194
rect 19796 107142 19798 107194
rect 19636 107140 19660 107142
rect 19716 107140 19740 107142
rect 19796 107140 19820 107142
rect 19580 107120 19876 107140
rect 19580 106108 19876 106128
rect 19636 106106 19660 106108
rect 19716 106106 19740 106108
rect 19796 106106 19820 106108
rect 19658 106054 19660 106106
rect 19722 106054 19734 106106
rect 19796 106054 19798 106106
rect 19636 106052 19660 106054
rect 19716 106052 19740 106054
rect 19796 106052 19820 106054
rect 19580 106032 19876 106052
rect 20628 105188 20680 105194
rect 20628 105130 20680 105136
rect 19580 105020 19876 105040
rect 19636 105018 19660 105020
rect 19716 105018 19740 105020
rect 19796 105018 19820 105020
rect 19658 104966 19660 105018
rect 19722 104966 19734 105018
rect 19796 104966 19798 105018
rect 19636 104964 19660 104966
rect 19716 104964 19740 104966
rect 19796 104964 19820 104966
rect 19580 104944 19876 104964
rect 20444 104848 20496 104854
rect 20444 104790 20496 104796
rect 19580 103932 19876 103952
rect 19636 103930 19660 103932
rect 19716 103930 19740 103932
rect 19796 103930 19820 103932
rect 19658 103878 19660 103930
rect 19722 103878 19734 103930
rect 19796 103878 19798 103930
rect 19636 103876 19660 103878
rect 19716 103876 19740 103878
rect 19796 103876 19820 103878
rect 19580 103856 19876 103876
rect 20456 103766 20484 104790
rect 18328 103760 18380 103766
rect 18328 103702 18380 103708
rect 20444 103760 20496 103766
rect 20444 103702 20496 103708
rect 20536 103760 20588 103766
rect 20536 103702 20588 103708
rect 18052 103624 18104 103630
rect 18052 103566 18104 103572
rect 16580 103488 16632 103494
rect 16580 103430 16632 103436
rect 16396 99340 16448 99346
rect 16396 99282 16448 99288
rect 16408 97646 16436 99282
rect 16592 97782 16620 103430
rect 18064 101998 18092 103566
rect 18340 103494 18368 103702
rect 18328 103488 18380 103494
rect 18328 103430 18380 103436
rect 19340 103488 19392 103494
rect 19340 103430 19392 103436
rect 18052 101992 18104 101998
rect 18052 101934 18104 101940
rect 17224 101516 17276 101522
rect 17224 101458 17276 101464
rect 16580 97776 16632 97782
rect 16580 97718 16632 97724
rect 16396 97640 16448 97646
rect 16396 97582 16448 97588
rect 16580 96416 16632 96422
rect 16580 96358 16632 96364
rect 16028 91860 16080 91866
rect 16028 91802 16080 91808
rect 16488 91724 16540 91730
rect 16488 91666 16540 91672
rect 16500 90030 16528 91666
rect 16488 90024 16540 90030
rect 16488 89966 16540 89972
rect 16304 46028 16356 46034
rect 16304 45970 16356 45976
rect 16028 42900 16080 42906
rect 16028 42842 16080 42848
rect 15936 36780 15988 36786
rect 15936 36722 15988 36728
rect 16040 28014 16068 42842
rect 16028 28008 16080 28014
rect 16028 27950 16080 27956
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14884 2876 14964 2904
rect 14832 2858 14884 2864
rect 15120 2774 15148 3878
rect 15028 2746 15148 2774
rect 15028 1986 15056 2746
rect 15304 2582 15332 13738
rect 15856 9178 15884 15506
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15396 3534 15424 3946
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15764 3058 15792 5510
rect 15948 4078 15976 23190
rect 16132 19334 16160 23258
rect 16040 19306 16160 19334
rect 16040 19174 16068 19306
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16028 19168 16080 19174
rect 16224 19122 16252 19246
rect 16028 19110 16080 19116
rect 16132 19094 16252 19122
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16040 14550 16068 18770
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 16132 11762 16160 19094
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16224 9926 16252 18906
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 14936 1958 15056 1986
rect 14936 800 14964 1958
rect 15304 800 15332 2382
rect 15580 800 15608 2926
rect 15856 800 15884 3878
rect 16316 3738 16344 45970
rect 16500 22094 16528 89966
rect 16592 88534 16620 96358
rect 16580 88528 16632 88534
rect 16580 88470 16632 88476
rect 17236 60734 17264 101458
rect 17316 100224 17368 100230
rect 17316 100166 17368 100172
rect 17328 90098 17356 100166
rect 18064 96490 18092 101934
rect 18604 99748 18656 99754
rect 18604 99690 18656 99696
rect 18236 97640 18288 97646
rect 18236 97582 18288 97588
rect 18248 96558 18276 97582
rect 18236 96552 18288 96558
rect 18236 96494 18288 96500
rect 18052 96484 18104 96490
rect 18052 96426 18104 96432
rect 17316 90092 17368 90098
rect 17316 90034 17368 90040
rect 18064 84194 18092 96426
rect 18248 86630 18276 96494
rect 18236 86624 18288 86630
rect 18236 86566 18288 86572
rect 17972 84166 18092 84194
rect 17868 73296 17920 73302
rect 17868 73238 17920 73244
rect 17776 69216 17828 69222
rect 17776 69158 17828 69164
rect 17144 60706 17264 60734
rect 17144 55894 17172 60706
rect 17316 58880 17368 58886
rect 17316 58822 17368 58828
rect 17224 57316 17276 57322
rect 17224 57258 17276 57264
rect 17236 56982 17264 57258
rect 17224 56976 17276 56982
rect 17224 56918 17276 56924
rect 17132 55888 17184 55894
rect 17132 55830 17184 55836
rect 17224 46980 17276 46986
rect 17224 46922 17276 46928
rect 16856 39432 16908 39438
rect 16856 39374 16908 39380
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16592 23254 16620 24890
rect 16672 24336 16724 24342
rect 16672 24278 16724 24284
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16408 22066 16528 22094
rect 16408 13802 16436 22066
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 19446 16528 19722
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 16500 18834 16528 19382
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16592 18222 16620 19994
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16592 16046 16620 17206
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 14482 16620 14894
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 12714 16436 13738
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16684 11014 16712 24278
rect 16868 21690 16896 39374
rect 17236 28626 17264 46922
rect 17328 40050 17356 58822
rect 17500 58336 17552 58342
rect 17500 58278 17552 58284
rect 17408 46572 17460 46578
rect 17408 46514 17460 46520
rect 17316 40044 17368 40050
rect 17316 39986 17368 39992
rect 17420 29102 17448 46514
rect 17512 45354 17540 58278
rect 17684 45552 17736 45558
rect 17684 45494 17736 45500
rect 17500 45348 17552 45354
rect 17500 45290 17552 45296
rect 17592 44396 17644 44402
rect 17592 44338 17644 44344
rect 17500 39500 17552 39506
rect 17500 39442 17552 39448
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17224 28620 17276 28626
rect 17224 28562 17276 28568
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17144 24138 17172 24618
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 17132 22024 17184 22030
rect 17130 21992 17132 22001
rect 17184 21992 17186 22001
rect 17130 21927 17186 21936
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16948 21480 17000 21486
rect 17132 21480 17184 21486
rect 16948 21422 17000 21428
rect 17130 21448 17132 21457
rect 17184 21448 17186 21457
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 19990 16804 20198
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16776 19514 16804 19654
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16776 18766 16804 19450
rect 16868 18834 16896 20402
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17270 16804 18158
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16868 15502 16896 15914
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16868 15366 16896 15438
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 14952 16816 14958
rect 16868 14940 16896 15302
rect 16816 14912 16896 14940
rect 16764 14894 16816 14900
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16960 9586 16988 21422
rect 17040 21412 17092 21418
rect 17130 21383 17186 21392
rect 17040 21354 17092 21360
rect 17052 21078 17080 21354
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17144 15978 17172 20742
rect 17236 19315 17264 24754
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 24614 17356 24686
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 17314 23760 17370 23769
rect 17314 23695 17370 23704
rect 17328 19446 17356 23695
rect 17420 23594 17448 24550
rect 17512 24274 17540 39442
rect 17604 29714 17632 44338
rect 17696 38894 17724 45494
rect 17684 38888 17736 38894
rect 17684 38830 17736 38836
rect 17788 38486 17816 69158
rect 17776 38480 17828 38486
rect 17776 38422 17828 38428
rect 17880 37330 17908 73238
rect 17868 37324 17920 37330
rect 17868 37266 17920 37272
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17788 25362 17816 34478
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17696 24274 17724 24618
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17696 24138 17724 24210
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17408 23588 17460 23594
rect 17408 23530 17460 23536
rect 17696 23322 17724 24074
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21690 17448 21966
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17420 21146 17448 21286
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17512 19990 17540 23122
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17682 21584 17738 21593
rect 17682 21519 17738 21528
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 17512 19718 17540 19926
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17222 19306 17278 19315
rect 17222 19241 17278 19250
rect 17224 19168 17276 19174
rect 17222 19136 17224 19145
rect 17500 19168 17552 19174
rect 17276 19136 17278 19145
rect 17500 19110 17552 19116
rect 17222 19071 17278 19080
rect 17314 19000 17370 19009
rect 17314 18935 17370 18944
rect 17328 18884 17356 18935
rect 17328 18856 17448 18884
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17132 15972 17184 15978
rect 17132 15914 17184 15920
rect 17144 15638 17172 15914
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 14822 17080 14894
rect 17144 14890 17172 15574
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16040 1850 16068 3538
rect 16040 1822 16160 1850
rect 16132 800 16160 1822
rect 16408 800 16436 3538
rect 16868 3466 16896 7278
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 800 16712 3334
rect 16960 3126 16988 3402
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17052 800 17080 2926
rect 17144 2582 17172 11086
rect 17236 10538 17264 18702
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17328 15570 17356 17478
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 17420 7750 17448 18856
rect 17512 17202 17540 19110
rect 17604 18834 17632 19382
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17604 18358 17632 18770
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17604 17814 17632 18294
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 17338 17632 17614
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17592 15564 17644 15570
rect 17696 15552 17724 21519
rect 17788 18222 17816 22034
rect 17972 22030 18000 84166
rect 18328 60308 18380 60314
rect 18328 60250 18380 60256
rect 18052 58336 18104 58342
rect 18052 58278 18104 58284
rect 18064 52494 18092 58278
rect 18236 56772 18288 56778
rect 18236 56714 18288 56720
rect 18052 52488 18104 52494
rect 18052 52430 18104 52436
rect 18052 37868 18104 37874
rect 18052 37810 18104 37816
rect 18064 33862 18092 37810
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 18248 28257 18276 56714
rect 18340 34134 18368 60250
rect 18512 60240 18564 60246
rect 18512 60182 18564 60188
rect 18420 50720 18472 50726
rect 18420 50662 18472 50668
rect 18328 34128 18380 34134
rect 18328 34070 18380 34076
rect 18432 33930 18460 50662
rect 18524 34950 18552 60182
rect 18616 35154 18644 99690
rect 19352 96762 19380 103430
rect 19580 102844 19876 102864
rect 19636 102842 19660 102844
rect 19716 102842 19740 102844
rect 19796 102842 19820 102844
rect 19658 102790 19660 102842
rect 19722 102790 19734 102842
rect 19796 102790 19798 102842
rect 19636 102788 19660 102790
rect 19716 102788 19740 102790
rect 19796 102788 19820 102790
rect 19580 102768 19876 102788
rect 19432 101924 19484 101930
rect 19432 101866 19484 101872
rect 19444 100910 19472 101866
rect 19580 101756 19876 101776
rect 19636 101754 19660 101756
rect 19716 101754 19740 101756
rect 19796 101754 19820 101756
rect 19658 101702 19660 101754
rect 19722 101702 19734 101754
rect 19796 101702 19798 101754
rect 19636 101700 19660 101702
rect 19716 101700 19740 101702
rect 19796 101700 19820 101702
rect 19580 101680 19876 101700
rect 20548 100910 20576 103702
rect 20640 101862 20668 105130
rect 20628 101856 20680 101862
rect 20628 101798 20680 101804
rect 19432 100904 19484 100910
rect 19432 100846 19484 100852
rect 20536 100904 20588 100910
rect 20536 100846 20588 100852
rect 19340 96756 19392 96762
rect 19340 96698 19392 96704
rect 19352 95538 19380 96698
rect 19340 95532 19392 95538
rect 19340 95474 19392 95480
rect 19444 93854 19472 100846
rect 19580 100668 19876 100688
rect 19636 100666 19660 100668
rect 19716 100666 19740 100668
rect 19796 100666 19820 100668
rect 19658 100614 19660 100666
rect 19722 100614 19734 100666
rect 19796 100614 19798 100666
rect 19636 100612 19660 100614
rect 19716 100612 19740 100614
rect 19796 100612 19820 100614
rect 19580 100592 19876 100612
rect 19580 99580 19876 99600
rect 19636 99578 19660 99580
rect 19716 99578 19740 99580
rect 19796 99578 19820 99580
rect 19658 99526 19660 99578
rect 19722 99526 19734 99578
rect 19796 99526 19798 99578
rect 19636 99524 19660 99526
rect 19716 99524 19740 99526
rect 19796 99524 19820 99526
rect 19580 99504 19876 99524
rect 20076 99204 20128 99210
rect 20076 99146 20128 99152
rect 19580 98492 19876 98512
rect 19636 98490 19660 98492
rect 19716 98490 19740 98492
rect 19796 98490 19820 98492
rect 19658 98438 19660 98490
rect 19722 98438 19734 98490
rect 19796 98438 19798 98490
rect 19636 98436 19660 98438
rect 19716 98436 19740 98438
rect 19796 98436 19820 98438
rect 19580 98416 19876 98436
rect 19580 97404 19876 97424
rect 19636 97402 19660 97404
rect 19716 97402 19740 97404
rect 19796 97402 19820 97404
rect 19658 97350 19660 97402
rect 19722 97350 19734 97402
rect 19796 97350 19798 97402
rect 19636 97348 19660 97350
rect 19716 97348 19740 97350
rect 19796 97348 19820 97350
rect 19580 97328 19876 97348
rect 19580 96316 19876 96336
rect 19636 96314 19660 96316
rect 19716 96314 19740 96316
rect 19796 96314 19820 96316
rect 19658 96262 19660 96314
rect 19722 96262 19734 96314
rect 19796 96262 19798 96314
rect 19636 96260 19660 96262
rect 19716 96260 19740 96262
rect 19796 96260 19820 96262
rect 19580 96240 19876 96260
rect 19984 95396 20036 95402
rect 19984 95338 20036 95344
rect 19580 95228 19876 95248
rect 19636 95226 19660 95228
rect 19716 95226 19740 95228
rect 19796 95226 19820 95228
rect 19658 95174 19660 95226
rect 19722 95174 19734 95226
rect 19796 95174 19798 95226
rect 19636 95172 19660 95174
rect 19716 95172 19740 95174
rect 19796 95172 19820 95174
rect 19580 95152 19876 95172
rect 19580 94140 19876 94160
rect 19636 94138 19660 94140
rect 19716 94138 19740 94140
rect 19796 94138 19820 94140
rect 19658 94086 19660 94138
rect 19722 94086 19734 94138
rect 19796 94086 19798 94138
rect 19636 94084 19660 94086
rect 19716 94084 19740 94086
rect 19796 94084 19820 94086
rect 19580 94064 19876 94084
rect 19352 93826 19472 93854
rect 19064 91792 19116 91798
rect 19064 91734 19116 91740
rect 18972 69352 19024 69358
rect 18972 69294 19024 69300
rect 18788 59628 18840 59634
rect 18788 59570 18840 59576
rect 18696 45484 18748 45490
rect 18696 45426 18748 45432
rect 18604 35148 18656 35154
rect 18604 35090 18656 35096
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18420 33924 18472 33930
rect 18420 33866 18472 33872
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18340 29034 18368 29582
rect 18328 29028 18380 29034
rect 18328 28970 18380 28976
rect 18340 28694 18368 28970
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18234 28248 18290 28257
rect 18234 28183 18290 28192
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 18064 24154 18092 28086
rect 18340 27946 18368 28630
rect 18604 28484 18656 28490
rect 18604 28426 18656 28432
rect 18328 27940 18380 27946
rect 18328 27882 18380 27888
rect 18340 27674 18368 27882
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 18616 26518 18644 28426
rect 18604 26512 18656 26518
rect 18604 26454 18656 26460
rect 18236 25764 18288 25770
rect 18156 25724 18236 25752
rect 18156 25362 18184 25724
rect 18420 25764 18472 25770
rect 18236 25706 18288 25712
rect 18340 25724 18420 25752
rect 18236 25424 18288 25430
rect 18340 25412 18368 25724
rect 18420 25706 18472 25712
rect 18288 25384 18368 25412
rect 18236 25366 18288 25372
rect 18144 25356 18196 25362
rect 18144 25298 18196 25304
rect 18156 24682 18184 25298
rect 18340 24682 18368 25384
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18328 24676 18380 24682
rect 18328 24618 18380 24624
rect 18340 24342 18368 24618
rect 18432 24410 18460 24686
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18064 24126 18276 24154
rect 18144 24064 18196 24070
rect 18050 24032 18106 24041
rect 18144 24006 18196 24012
rect 18050 23967 18106 23976
rect 18064 23866 18092 23967
rect 18156 23866 18184 24006
rect 18052 23860 18104 23866
rect 18052 23802 18104 23808
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18248 23338 18276 24126
rect 18156 23310 18276 23338
rect 18340 23322 18368 24278
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18328 23316 18380 23322
rect 18156 23050 18184 23310
rect 18328 23258 18380 23264
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17880 19394 17908 20946
rect 17972 19990 18000 21830
rect 18064 21622 18092 22646
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18064 21078 18092 21558
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 18052 20528 18104 20534
rect 18052 20470 18104 20476
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17880 19366 18000 19394
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17880 18970 17908 19246
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17972 18850 18000 19366
rect 17880 18822 18000 18850
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17644 15524 17724 15552
rect 17592 15506 17644 15512
rect 17512 11830 17540 15506
rect 17696 15094 17724 15524
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17696 9382 17724 14894
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17328 2774 17356 6802
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17420 3670 17448 5510
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17604 3194 17632 3878
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17328 2746 17448 2774
rect 17420 2582 17448 2746
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17328 800 17356 2450
rect 17696 1714 17724 3334
rect 17788 2854 17816 18158
rect 17880 13258 17908 18822
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17972 18426 18000 18702
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18064 16538 18092 20470
rect 18156 17218 18184 22510
rect 18248 21894 18276 23122
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18248 20262 18276 20946
rect 18340 20942 18368 21422
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18248 18902 18276 19178
rect 18432 18970 18460 24006
rect 18524 23662 18552 24618
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18616 23730 18644 24550
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18524 23186 18552 23598
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18512 23044 18564 23050
rect 18512 22986 18564 22992
rect 18524 21690 18552 22986
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18616 22234 18644 22646
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18616 21593 18644 21626
rect 18602 21584 18658 21593
rect 18602 21519 18658 21528
rect 18510 21448 18566 21457
rect 18510 21383 18512 21392
rect 18564 21383 18566 21392
rect 18512 21354 18564 21360
rect 18524 21078 18552 21354
rect 18512 21072 18564 21078
rect 18512 21014 18564 21020
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18616 18902 18644 19450
rect 18236 18896 18288 18902
rect 18604 18896 18656 18902
rect 18236 18838 18288 18844
rect 18418 18864 18474 18873
rect 18248 18290 18276 18838
rect 18604 18838 18656 18844
rect 18418 18799 18420 18808
rect 18472 18799 18474 18808
rect 18420 18770 18472 18776
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 17746 18276 18226
rect 18340 17882 18368 18702
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18156 17190 18276 17218
rect 18064 16510 18184 16538
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14414 18092 14894
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17604 1686 17724 1714
rect 17604 800 17632 1686
rect 17880 800 17908 4014
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 2990 18000 3878
rect 18156 3670 18184 16510
rect 18248 9654 18276 17190
rect 18432 15978 18460 17546
rect 18616 16794 18644 18702
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18156 800 18184 2926
rect 18524 800 18552 3334
rect 18708 3194 18736 45426
rect 18800 33590 18828 59570
rect 18880 57792 18932 57798
rect 18880 57734 18932 57740
rect 18788 33584 18840 33590
rect 18788 33526 18840 33532
rect 18892 29510 18920 57734
rect 18984 39642 19012 69294
rect 18972 39636 19024 39642
rect 18972 39578 19024 39584
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 18892 29102 18920 29242
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 18800 21593 18828 28018
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 18892 25362 18920 26182
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18878 23896 18934 23905
rect 18878 23831 18934 23840
rect 18892 22778 18920 23831
rect 18880 22772 18932 22778
rect 18880 22714 18932 22720
rect 18892 22166 18920 22714
rect 18880 22160 18932 22166
rect 18880 22102 18932 22108
rect 18880 22024 18932 22030
rect 18878 21992 18880 22001
rect 18932 21992 18934 22001
rect 18878 21927 18934 21936
rect 18880 21616 18932 21622
rect 18786 21584 18842 21593
rect 18880 21558 18932 21564
rect 18786 21519 18842 21528
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18800 11082 18828 21422
rect 18892 18222 18920 21558
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18892 17542 18920 18158
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18984 11558 19012 29650
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18892 3602 18920 6326
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18800 800 18828 3470
rect 19076 2582 19104 91734
rect 19352 89962 19380 93826
rect 19580 93052 19876 93072
rect 19636 93050 19660 93052
rect 19716 93050 19740 93052
rect 19796 93050 19820 93052
rect 19658 92998 19660 93050
rect 19722 92998 19734 93050
rect 19796 92998 19798 93050
rect 19636 92996 19660 92998
rect 19716 92996 19740 92998
rect 19796 92996 19820 92998
rect 19580 92976 19876 92996
rect 19996 92410 20024 95338
rect 20088 93854 20116 99146
rect 20640 95402 20668 101798
rect 20628 95396 20680 95402
rect 20628 95338 20680 95344
rect 20088 93826 20208 93854
rect 19984 92404 20036 92410
rect 19984 92346 20036 92352
rect 20076 92132 20128 92138
rect 20076 92074 20128 92080
rect 19580 91964 19876 91984
rect 19636 91962 19660 91964
rect 19716 91962 19740 91964
rect 19796 91962 19820 91964
rect 19658 91910 19660 91962
rect 19722 91910 19734 91962
rect 19796 91910 19798 91962
rect 19636 91908 19660 91910
rect 19716 91908 19740 91910
rect 19796 91908 19820 91910
rect 19580 91888 19876 91908
rect 19580 90876 19876 90896
rect 19636 90874 19660 90876
rect 19716 90874 19740 90876
rect 19796 90874 19820 90876
rect 19658 90822 19660 90874
rect 19722 90822 19734 90874
rect 19796 90822 19798 90874
rect 19636 90820 19660 90822
rect 19716 90820 19740 90822
rect 19796 90820 19820 90822
rect 19580 90800 19876 90820
rect 19892 90636 19944 90642
rect 19892 90578 19944 90584
rect 19340 89956 19392 89962
rect 19340 89898 19392 89904
rect 19352 86766 19380 89898
rect 19580 89788 19876 89808
rect 19636 89786 19660 89788
rect 19716 89786 19740 89788
rect 19796 89786 19820 89788
rect 19658 89734 19660 89786
rect 19722 89734 19734 89786
rect 19796 89734 19798 89786
rect 19636 89732 19660 89734
rect 19716 89732 19740 89734
rect 19796 89732 19820 89734
rect 19580 89712 19876 89732
rect 19580 88700 19876 88720
rect 19636 88698 19660 88700
rect 19716 88698 19740 88700
rect 19796 88698 19820 88700
rect 19658 88646 19660 88698
rect 19722 88646 19734 88698
rect 19796 88646 19798 88698
rect 19636 88644 19660 88646
rect 19716 88644 19740 88646
rect 19796 88644 19820 88646
rect 19580 88624 19876 88644
rect 19580 87612 19876 87632
rect 19636 87610 19660 87612
rect 19716 87610 19740 87612
rect 19796 87610 19820 87612
rect 19658 87558 19660 87610
rect 19722 87558 19734 87610
rect 19796 87558 19798 87610
rect 19636 87556 19660 87558
rect 19716 87556 19740 87558
rect 19796 87556 19820 87558
rect 19580 87536 19876 87556
rect 19340 86760 19392 86766
rect 19340 86702 19392 86708
rect 19432 86692 19484 86698
rect 19432 86634 19484 86640
rect 19340 86624 19392 86630
rect 19340 86566 19392 86572
rect 19248 76288 19300 76294
rect 19248 76230 19300 76236
rect 19156 75540 19208 75546
rect 19156 75482 19208 75488
rect 19168 43314 19196 75482
rect 19260 44402 19288 76230
rect 19248 44396 19300 44402
rect 19248 44338 19300 44344
rect 19156 43308 19208 43314
rect 19156 43250 19208 43256
rect 19248 29844 19300 29850
rect 19168 29804 19248 29832
rect 19168 29034 19196 29804
rect 19248 29786 19300 29792
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28422 19196 28970
rect 19248 28688 19300 28694
rect 19248 28630 19300 28636
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19168 27946 19196 28358
rect 19156 27940 19208 27946
rect 19156 27882 19208 27888
rect 19168 23798 19196 27882
rect 19260 27674 19288 28630
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19260 24750 19288 27610
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19260 23905 19288 24346
rect 19246 23896 19302 23905
rect 19246 23831 19302 23840
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 22642 19196 23598
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19168 22166 19196 22578
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19168 21418 19196 22102
rect 19246 21584 19302 21593
rect 19246 21519 19302 21528
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19260 21298 19288 21519
rect 19168 21270 19288 21298
rect 19168 15026 19196 21270
rect 19352 19786 19380 86566
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19444 19394 19472 86634
rect 19580 86524 19876 86544
rect 19636 86522 19660 86524
rect 19716 86522 19740 86524
rect 19796 86522 19820 86524
rect 19658 86470 19660 86522
rect 19722 86470 19734 86522
rect 19796 86470 19798 86522
rect 19636 86468 19660 86470
rect 19716 86468 19740 86470
rect 19796 86468 19820 86470
rect 19580 86448 19876 86468
rect 19904 86290 19932 90578
rect 20088 86834 20116 92074
rect 20076 86828 20128 86834
rect 20076 86770 20128 86776
rect 20088 86426 20116 86770
rect 20180 86698 20208 93826
rect 20168 86692 20220 86698
rect 20168 86634 20220 86640
rect 20076 86420 20128 86426
rect 20076 86362 20128 86368
rect 19892 86284 19944 86290
rect 19892 86226 19944 86232
rect 19580 85436 19876 85456
rect 19636 85434 19660 85436
rect 19716 85434 19740 85436
rect 19796 85434 19820 85436
rect 19658 85382 19660 85434
rect 19722 85382 19734 85434
rect 19796 85382 19798 85434
rect 19636 85380 19660 85382
rect 19716 85380 19740 85382
rect 19796 85380 19820 85382
rect 19580 85360 19876 85380
rect 19580 84348 19876 84368
rect 19636 84346 19660 84348
rect 19716 84346 19740 84348
rect 19796 84346 19820 84348
rect 19658 84294 19660 84346
rect 19722 84294 19734 84346
rect 19796 84294 19798 84346
rect 19636 84292 19660 84294
rect 19716 84292 19740 84294
rect 19796 84292 19820 84294
rect 19580 84272 19876 84292
rect 19580 83260 19876 83280
rect 19636 83258 19660 83260
rect 19716 83258 19740 83260
rect 19796 83258 19820 83260
rect 19658 83206 19660 83258
rect 19722 83206 19734 83258
rect 19796 83206 19798 83258
rect 19636 83204 19660 83206
rect 19716 83204 19740 83206
rect 19796 83204 19820 83206
rect 19580 83184 19876 83204
rect 19580 82172 19876 82192
rect 19636 82170 19660 82172
rect 19716 82170 19740 82172
rect 19796 82170 19820 82172
rect 19658 82118 19660 82170
rect 19722 82118 19734 82170
rect 19796 82118 19798 82170
rect 19636 82116 19660 82118
rect 19716 82116 19740 82118
rect 19796 82116 19820 82118
rect 19580 82096 19876 82116
rect 19580 81084 19876 81104
rect 19636 81082 19660 81084
rect 19716 81082 19740 81084
rect 19796 81082 19820 81084
rect 19658 81030 19660 81082
rect 19722 81030 19734 81082
rect 19796 81030 19798 81082
rect 19636 81028 19660 81030
rect 19716 81028 19740 81030
rect 19796 81028 19820 81030
rect 19580 81008 19876 81028
rect 19580 79996 19876 80016
rect 19636 79994 19660 79996
rect 19716 79994 19740 79996
rect 19796 79994 19820 79996
rect 19658 79942 19660 79994
rect 19722 79942 19734 79994
rect 19796 79942 19798 79994
rect 19636 79940 19660 79942
rect 19716 79940 19740 79942
rect 19796 79940 19820 79942
rect 19580 79920 19876 79940
rect 19580 78908 19876 78928
rect 19636 78906 19660 78908
rect 19716 78906 19740 78908
rect 19796 78906 19820 78908
rect 19658 78854 19660 78906
rect 19722 78854 19734 78906
rect 19796 78854 19798 78906
rect 19636 78852 19660 78854
rect 19716 78852 19740 78854
rect 19796 78852 19820 78854
rect 19580 78832 19876 78852
rect 19580 77820 19876 77840
rect 19636 77818 19660 77820
rect 19716 77818 19740 77820
rect 19796 77818 19820 77820
rect 19658 77766 19660 77818
rect 19722 77766 19734 77818
rect 19796 77766 19798 77818
rect 19636 77764 19660 77766
rect 19716 77764 19740 77766
rect 19796 77764 19820 77766
rect 19580 77744 19876 77764
rect 19580 76732 19876 76752
rect 19636 76730 19660 76732
rect 19716 76730 19740 76732
rect 19796 76730 19820 76732
rect 19658 76678 19660 76730
rect 19722 76678 19734 76730
rect 19796 76678 19798 76730
rect 19636 76676 19660 76678
rect 19716 76676 19740 76678
rect 19796 76676 19820 76678
rect 19580 76656 19876 76676
rect 19580 75644 19876 75664
rect 19636 75642 19660 75644
rect 19716 75642 19740 75644
rect 19796 75642 19820 75644
rect 19658 75590 19660 75642
rect 19722 75590 19734 75642
rect 19796 75590 19798 75642
rect 19636 75588 19660 75590
rect 19716 75588 19740 75590
rect 19796 75588 19820 75590
rect 19580 75568 19876 75588
rect 19580 74556 19876 74576
rect 19636 74554 19660 74556
rect 19716 74554 19740 74556
rect 19796 74554 19820 74556
rect 19658 74502 19660 74554
rect 19722 74502 19734 74554
rect 19796 74502 19798 74554
rect 19636 74500 19660 74502
rect 19716 74500 19740 74502
rect 19796 74500 19820 74502
rect 19580 74480 19876 74500
rect 19580 73468 19876 73488
rect 19636 73466 19660 73468
rect 19716 73466 19740 73468
rect 19796 73466 19820 73468
rect 19658 73414 19660 73466
rect 19722 73414 19734 73466
rect 19796 73414 19798 73466
rect 19636 73412 19660 73414
rect 19716 73412 19740 73414
rect 19796 73412 19820 73414
rect 19580 73392 19876 73412
rect 19580 72380 19876 72400
rect 19636 72378 19660 72380
rect 19716 72378 19740 72380
rect 19796 72378 19820 72380
rect 19658 72326 19660 72378
rect 19722 72326 19734 72378
rect 19796 72326 19798 72378
rect 19636 72324 19660 72326
rect 19716 72324 19740 72326
rect 19796 72324 19820 72326
rect 19580 72304 19876 72324
rect 19580 71292 19876 71312
rect 19636 71290 19660 71292
rect 19716 71290 19740 71292
rect 19796 71290 19820 71292
rect 19658 71238 19660 71290
rect 19722 71238 19734 71290
rect 19796 71238 19798 71290
rect 19636 71236 19660 71238
rect 19716 71236 19740 71238
rect 19796 71236 19820 71238
rect 19580 71216 19876 71236
rect 19580 70204 19876 70224
rect 19636 70202 19660 70204
rect 19716 70202 19740 70204
rect 19796 70202 19820 70204
rect 19658 70150 19660 70202
rect 19722 70150 19734 70202
rect 19796 70150 19798 70202
rect 19636 70148 19660 70150
rect 19716 70148 19740 70150
rect 19796 70148 19820 70150
rect 19580 70128 19876 70148
rect 19580 69116 19876 69136
rect 19636 69114 19660 69116
rect 19716 69114 19740 69116
rect 19796 69114 19820 69116
rect 19658 69062 19660 69114
rect 19722 69062 19734 69114
rect 19796 69062 19798 69114
rect 19636 69060 19660 69062
rect 19716 69060 19740 69062
rect 19796 69060 19820 69062
rect 19580 69040 19876 69060
rect 19580 68028 19876 68048
rect 19636 68026 19660 68028
rect 19716 68026 19740 68028
rect 19796 68026 19820 68028
rect 19658 67974 19660 68026
rect 19722 67974 19734 68026
rect 19796 67974 19798 68026
rect 19636 67972 19660 67974
rect 19716 67972 19740 67974
rect 19796 67972 19820 67974
rect 19580 67952 19876 67972
rect 19580 66940 19876 66960
rect 19636 66938 19660 66940
rect 19716 66938 19740 66940
rect 19796 66938 19820 66940
rect 19658 66886 19660 66938
rect 19722 66886 19734 66938
rect 19796 66886 19798 66938
rect 19636 66884 19660 66886
rect 19716 66884 19740 66886
rect 19796 66884 19820 66886
rect 19580 66864 19876 66884
rect 19580 65852 19876 65872
rect 19636 65850 19660 65852
rect 19716 65850 19740 65852
rect 19796 65850 19820 65852
rect 19658 65798 19660 65850
rect 19722 65798 19734 65850
rect 19796 65798 19798 65850
rect 19636 65796 19660 65798
rect 19716 65796 19740 65798
rect 19796 65796 19820 65798
rect 19580 65776 19876 65796
rect 19580 64764 19876 64784
rect 19636 64762 19660 64764
rect 19716 64762 19740 64764
rect 19796 64762 19820 64764
rect 19658 64710 19660 64762
rect 19722 64710 19734 64762
rect 19796 64710 19798 64762
rect 19636 64708 19660 64710
rect 19716 64708 19740 64710
rect 19796 64708 19820 64710
rect 19580 64688 19876 64708
rect 19580 63676 19876 63696
rect 19636 63674 19660 63676
rect 19716 63674 19740 63676
rect 19796 63674 19820 63676
rect 19658 63622 19660 63674
rect 19722 63622 19734 63674
rect 19796 63622 19798 63674
rect 19636 63620 19660 63622
rect 19716 63620 19740 63622
rect 19796 63620 19820 63622
rect 19580 63600 19876 63620
rect 19580 62588 19876 62608
rect 19636 62586 19660 62588
rect 19716 62586 19740 62588
rect 19796 62586 19820 62588
rect 19658 62534 19660 62586
rect 19722 62534 19734 62586
rect 19796 62534 19798 62586
rect 19636 62532 19660 62534
rect 19716 62532 19740 62534
rect 19796 62532 19820 62534
rect 19580 62512 19876 62532
rect 19580 61500 19876 61520
rect 19636 61498 19660 61500
rect 19716 61498 19740 61500
rect 19796 61498 19820 61500
rect 19658 61446 19660 61498
rect 19722 61446 19734 61498
rect 19796 61446 19798 61498
rect 19636 61444 19660 61446
rect 19716 61444 19740 61446
rect 19796 61444 19820 61446
rect 19580 61424 19876 61444
rect 19580 60412 19876 60432
rect 19636 60410 19660 60412
rect 19716 60410 19740 60412
rect 19796 60410 19820 60412
rect 19658 60358 19660 60410
rect 19722 60358 19734 60410
rect 19796 60358 19798 60410
rect 19636 60356 19660 60358
rect 19716 60356 19740 60358
rect 19796 60356 19820 60358
rect 19580 60336 19876 60356
rect 19580 59324 19876 59344
rect 19636 59322 19660 59324
rect 19716 59322 19740 59324
rect 19796 59322 19820 59324
rect 19658 59270 19660 59322
rect 19722 59270 19734 59322
rect 19796 59270 19798 59322
rect 19636 59268 19660 59270
rect 19716 59268 19740 59270
rect 19796 59268 19820 59270
rect 19580 59248 19876 59268
rect 19580 58236 19876 58256
rect 19636 58234 19660 58236
rect 19716 58234 19740 58236
rect 19796 58234 19820 58236
rect 19658 58182 19660 58234
rect 19722 58182 19734 58234
rect 19796 58182 19798 58234
rect 19636 58180 19660 58182
rect 19716 58180 19740 58182
rect 19796 58180 19820 58182
rect 19580 58160 19876 58180
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 19904 48498 19932 86226
rect 20168 77716 20220 77722
rect 20168 77658 20220 77664
rect 19984 64932 20036 64938
rect 19984 64874 20036 64880
rect 19996 60734 20024 64874
rect 19996 60706 20116 60734
rect 19984 59968 20036 59974
rect 19984 59910 20036 59916
rect 19996 54874 20024 59910
rect 20088 55350 20116 60706
rect 20180 57934 20208 77658
rect 20260 74656 20312 74662
rect 20260 74598 20312 74604
rect 20168 57928 20220 57934
rect 20168 57870 20220 57876
rect 20076 55344 20128 55350
rect 20076 55286 20128 55292
rect 19984 54868 20036 54874
rect 19984 54810 20036 54816
rect 20168 52556 20220 52562
rect 20168 52498 20220 52504
rect 20076 48748 20128 48754
rect 20076 48690 20128 48696
rect 19982 48512 20038 48521
rect 19904 48470 19982 48498
rect 19580 48444 19876 48464
rect 19982 48447 20038 48456
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 19984 48272 20036 48278
rect 19890 48240 19946 48249
rect 19984 48214 20036 48220
rect 19890 48175 19946 48184
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19614 28656 19670 28665
rect 19614 28591 19670 28600
rect 19798 28656 19854 28665
rect 19798 28591 19800 28600
rect 19628 28490 19656 28591
rect 19852 28591 19854 28600
rect 19800 28562 19852 28568
rect 19616 28484 19668 28490
rect 19616 28426 19668 28432
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19614 27568 19670 27577
rect 19614 27503 19670 27512
rect 19628 27334 19656 27503
rect 19616 27328 19668 27334
rect 19616 27270 19668 27276
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19798 24168 19854 24177
rect 19798 24103 19854 24112
rect 19616 24064 19668 24070
rect 19614 24032 19616 24041
rect 19668 24032 19670 24041
rect 19614 23967 19670 23976
rect 19812 23662 19840 24103
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19352 19366 19472 19394
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19260 18970 19288 19178
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19352 18426 19380 19366
rect 19432 19304 19484 19310
rect 19536 19281 19564 19926
rect 19432 19246 19484 19252
rect 19522 19272 19578 19281
rect 19444 18834 19472 19246
rect 19522 19207 19578 19216
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19522 18864 19578 18873
rect 19432 18828 19484 18834
rect 19522 18799 19578 18808
rect 19432 18770 19484 18776
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19444 18290 19472 18770
rect 19536 18698 19564 18799
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19444 17746 19472 18226
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19352 13326 19380 17002
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19904 12374 19932 48175
rect 19996 30054 20024 48214
rect 20088 41682 20116 48690
rect 20076 41676 20128 41682
rect 20076 41618 20128 41624
rect 20180 41562 20208 52498
rect 20088 41534 20208 41562
rect 20088 36530 20116 41534
rect 20168 41472 20220 41478
rect 20168 41414 20220 41420
rect 20180 36650 20208 41414
rect 20272 40186 20300 74598
rect 20352 73364 20404 73370
rect 20352 73306 20404 73312
rect 20260 40180 20312 40186
rect 20260 40122 20312 40128
rect 20364 37194 20392 73306
rect 20536 63300 20588 63306
rect 20536 63242 20588 63248
rect 20548 60734 20576 63242
rect 20456 60706 20576 60734
rect 20352 37188 20404 37194
rect 20352 37130 20404 37136
rect 20168 36644 20220 36650
rect 20168 36586 20220 36592
rect 20088 36502 20208 36530
rect 20076 31136 20128 31142
rect 20076 31078 20128 31084
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19982 28792 20038 28801
rect 19982 28727 19984 28736
rect 20036 28727 20038 28736
rect 19984 28698 20036 28704
rect 20088 28665 20116 31078
rect 20180 28762 20208 36502
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20168 28756 20220 28762
rect 20168 28698 20220 28704
rect 20074 28656 20130 28665
rect 19984 28620 20036 28626
rect 20074 28591 20130 28600
rect 19984 28562 20036 28568
rect 19996 27946 20024 28562
rect 20272 28370 20300 29242
rect 20180 28342 20300 28370
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 20074 27704 20130 27713
rect 20074 27639 20076 27648
rect 20128 27639 20130 27648
rect 20076 27610 20128 27616
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19996 26994 20024 27406
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19996 26246 20024 26930
rect 20076 26852 20128 26858
rect 20076 26794 20128 26800
rect 20088 26586 20116 26794
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19984 26240 20036 26246
rect 19984 26182 20036 26188
rect 19996 24274 20024 26182
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 20088 24682 20116 25162
rect 20180 25158 20208 28342
rect 20260 27872 20312 27878
rect 20260 27814 20312 27820
rect 20272 27470 20300 27814
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20260 26512 20312 26518
rect 20260 26454 20312 26460
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19982 23896 20038 23905
rect 19982 23831 20038 23840
rect 19996 23662 20024 23831
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19996 21434 20024 23258
rect 20088 23186 20116 24618
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20180 23118 20208 24210
rect 20168 23112 20220 23118
rect 20168 23054 20220 23060
rect 20180 22098 20208 23054
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 20180 21554 20208 22034
rect 20168 21548 20220 21554
rect 20168 21490 20220 21496
rect 19996 21406 20208 21434
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19996 21026 20024 21286
rect 19996 20998 20116 21026
rect 19984 20868 20036 20874
rect 19984 20810 20036 20816
rect 19996 19310 20024 20810
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19996 18902 20024 19110
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 20088 16946 20116 20998
rect 19996 16918 20116 16946
rect 19996 14618 20024 16918
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19892 12368 19944 12374
rect 19892 12310 19944 12316
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19904 11150 19932 12310
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 20088 10470 20116 16730
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 19168 2446 19196 8366
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19076 800 19104 2382
rect 19352 800 19380 2790
rect 19444 2122 19472 4014
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19996 3398 20024 3674
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19536 3058 19564 3334
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 20088 2990 20116 6938
rect 20180 6186 20208 21406
rect 20272 11150 20300 26454
rect 20364 19990 20392 29650
rect 20352 19984 20404 19990
rect 20352 19926 20404 19932
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20364 6254 20392 19790
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20456 3738 20484 60706
rect 20628 57928 20680 57934
rect 20628 57870 20680 57876
rect 20536 57520 20588 57526
rect 20536 57462 20588 57468
rect 20548 35766 20576 57462
rect 20640 55146 20668 57870
rect 20628 55140 20680 55146
rect 20628 55082 20680 55088
rect 20628 54868 20680 54874
rect 20628 54810 20680 54816
rect 20536 35760 20588 35766
rect 20536 35702 20588 35708
rect 20640 34610 20668 54810
rect 20732 51066 20760 112406
rect 21548 108452 21600 108458
rect 21548 108394 21600 108400
rect 21272 104712 21324 104718
rect 21272 104654 21324 104660
rect 21284 103834 21312 104654
rect 21272 103828 21324 103834
rect 21272 103770 21324 103776
rect 21456 101448 21508 101454
rect 21456 101390 21508 101396
rect 21468 98870 21496 101390
rect 21456 98864 21508 98870
rect 21456 98806 21508 98812
rect 21272 98660 21324 98666
rect 21272 98602 21324 98608
rect 20904 63368 20956 63374
rect 20904 63310 20956 63316
rect 20812 58880 20864 58886
rect 20812 58822 20864 58828
rect 20720 51060 20772 51066
rect 20720 51002 20772 51008
rect 20720 45824 20772 45830
rect 20720 45766 20772 45772
rect 20732 43450 20760 45766
rect 20720 43444 20772 43450
rect 20720 43386 20772 43392
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20824 33153 20852 58822
rect 20916 35086 20944 63310
rect 21180 62280 21232 62286
rect 21180 62222 21232 62228
rect 20996 50312 21048 50318
rect 20996 50254 21048 50260
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20810 33144 20866 33153
rect 20810 33079 20866 33088
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20536 27940 20588 27946
rect 20536 27882 20588 27888
rect 20548 20602 20576 27882
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20640 23322 20668 27542
rect 20732 23769 20760 28970
rect 20812 28416 20864 28422
rect 20812 28358 20864 28364
rect 20824 27538 20852 28358
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 20812 27532 20864 27538
rect 20812 27474 20864 27480
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20824 25906 20852 26862
rect 20916 26382 20944 27610
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20812 25356 20864 25362
rect 20812 25298 20864 25304
rect 20718 23760 20774 23769
rect 20718 23695 20774 23704
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20640 21672 20668 22918
rect 20732 22166 20760 23598
rect 20824 23322 20852 25298
rect 20904 25152 20956 25158
rect 20904 25094 20956 25100
rect 20916 24954 20944 25094
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20902 24848 20958 24857
rect 20902 24783 20958 24792
rect 20916 23662 20944 24783
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20904 23520 20956 23526
rect 20904 23462 20956 23468
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20640 21644 20760 21672
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20640 20874 20668 21490
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20732 20346 20760 21644
rect 20824 21078 20852 23122
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20640 20318 20760 20346
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20548 15722 20576 19722
rect 20640 18970 20668 20318
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20732 18834 20760 20198
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20824 18970 20852 19110
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20548 15694 20668 15722
rect 20640 12782 20668 15694
rect 20732 12850 20760 18362
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 12374 20576 12582
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20640 7546 20668 12718
rect 20824 11898 20852 18906
rect 20916 17134 20944 23462
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20916 4826 20944 16934
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 4214 20760 4422
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19444 2094 19656 2122
rect 19628 800 19656 2094
rect 19904 800 19932 2450
rect 20272 800 20300 2858
rect 20548 800 20576 4014
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20640 3126 20668 3878
rect 21008 3194 21036 50254
rect 21088 50244 21140 50250
rect 21088 50186 21140 50192
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20628 3120 20680 3126
rect 21100 3074 21128 50186
rect 21192 4282 21220 62222
rect 21284 54602 21312 98602
rect 21456 62824 21508 62830
rect 21456 62766 21508 62772
rect 21272 54596 21324 54602
rect 21272 54538 21324 54544
rect 21272 51468 21324 51474
rect 21272 51410 21324 51416
rect 21284 48754 21312 51410
rect 21364 49904 21416 49910
rect 21364 49846 21416 49852
rect 21272 48748 21324 48754
rect 21272 48690 21324 48696
rect 21376 46034 21404 49846
rect 21364 46028 21416 46034
rect 21364 45970 21416 45976
rect 21364 40384 21416 40390
rect 21364 40326 21416 40332
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21284 26790 21312 27882
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 21284 26246 21312 26726
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21270 25936 21326 25945
rect 21270 25871 21326 25880
rect 21284 24886 21312 25871
rect 21376 25362 21404 40326
rect 21468 36242 21496 62766
rect 21560 51610 21588 108394
rect 21652 103834 21680 113358
rect 21928 109034 21956 116175
rect 22008 115592 22060 115598
rect 22008 115534 22060 115540
rect 22098 115560 22154 115569
rect 22020 115433 22048 115534
rect 22098 115495 22154 115504
rect 22006 115424 22062 115433
rect 22006 115359 22062 115368
rect 22112 115258 22140 115495
rect 22100 115252 22152 115258
rect 22100 115194 22152 115200
rect 22296 114646 22324 116742
rect 22480 116550 22508 119200
rect 22558 117192 22614 117201
rect 22558 117127 22614 117136
rect 22376 116544 22428 116550
rect 22376 116486 22428 116492
rect 22468 116544 22520 116550
rect 22468 116486 22520 116492
rect 22388 116278 22416 116486
rect 22376 116272 22428 116278
rect 22376 116214 22428 116220
rect 22572 115682 22600 117127
rect 22652 116816 22704 116822
rect 22652 116758 22704 116764
rect 22664 116346 22692 116758
rect 22652 116340 22704 116346
rect 22652 116282 22704 116288
rect 22480 115654 22600 115682
rect 22192 114640 22244 114646
rect 22192 114582 22244 114588
rect 22284 114640 22336 114646
rect 22284 114582 22336 114588
rect 22204 113966 22232 114582
rect 22192 113960 22244 113966
rect 22192 113902 22244 113908
rect 22480 109034 22508 115654
rect 22560 115592 22612 115598
rect 22756 115580 22784 119200
rect 22940 117366 22968 119200
rect 22928 117360 22980 117366
rect 22928 117302 22980 117308
rect 23124 116346 23152 119200
rect 23202 117328 23258 117337
rect 23202 117263 23258 117272
rect 23216 117162 23244 117263
rect 23204 117156 23256 117162
rect 23204 117098 23256 117104
rect 23296 117156 23348 117162
rect 23296 117098 23348 117104
rect 23202 117056 23258 117065
rect 23202 116991 23258 117000
rect 22928 116340 22980 116346
rect 22928 116282 22980 116288
rect 23112 116340 23164 116346
rect 23112 116282 23164 116288
rect 22940 115666 22968 116282
rect 23112 116204 23164 116210
rect 23112 116146 23164 116152
rect 23020 116068 23072 116074
rect 23020 116010 23072 116016
rect 23032 115666 23060 116010
rect 22928 115660 22980 115666
rect 22928 115602 22980 115608
rect 23020 115660 23072 115666
rect 23020 115602 23072 115608
rect 22756 115552 22876 115580
rect 22560 115534 22612 115540
rect 22572 114714 22600 115534
rect 22560 114708 22612 114714
rect 22560 114650 22612 114656
rect 22744 114572 22796 114578
rect 22744 114514 22796 114520
rect 22756 114102 22784 114514
rect 22744 114096 22796 114102
rect 22744 114038 22796 114044
rect 22848 113966 22876 115552
rect 23124 114986 23152 116146
rect 23216 115530 23244 116991
rect 23308 115802 23336 117098
rect 23296 115796 23348 115802
rect 23296 115738 23348 115744
rect 23204 115524 23256 115530
rect 23204 115466 23256 115472
rect 23294 115152 23350 115161
rect 23294 115087 23350 115096
rect 23112 114980 23164 114986
rect 23112 114922 23164 114928
rect 23308 114918 23336 115087
rect 23296 114912 23348 114918
rect 23296 114854 23348 114860
rect 23400 113966 23428 119200
rect 23584 115802 23612 119200
rect 23664 116884 23716 116890
rect 23664 116826 23716 116832
rect 23572 115796 23624 115802
rect 23572 115738 23624 115744
rect 23676 114714 23704 116826
rect 23768 116346 23796 119200
rect 23940 117088 23992 117094
rect 23940 117030 23992 117036
rect 23756 116340 23808 116346
rect 23756 116282 23808 116288
rect 23952 115841 23980 117030
rect 23938 115832 23994 115841
rect 23938 115767 23994 115776
rect 23848 115660 23900 115666
rect 23848 115602 23900 115608
rect 23664 114708 23716 114714
rect 23664 114650 23716 114656
rect 23860 114578 23888 115602
rect 23848 114572 23900 114578
rect 23848 114514 23900 114520
rect 24044 113966 24072 119200
rect 24124 117156 24176 117162
rect 24124 117098 24176 117104
rect 24136 115530 24164 117098
rect 24228 116890 24256 119200
rect 24412 116906 24440 119200
rect 24412 116890 24532 116906
rect 24216 116884 24268 116890
rect 24412 116884 24544 116890
rect 24412 116878 24492 116884
rect 24216 116826 24268 116832
rect 24492 116826 24544 116832
rect 24308 116748 24360 116754
rect 24308 116690 24360 116696
rect 24320 115666 24348 116690
rect 24490 115968 24546 115977
rect 24490 115903 24546 115912
rect 24308 115660 24360 115666
rect 24308 115602 24360 115608
rect 24124 115524 24176 115530
rect 24124 115466 24176 115472
rect 24504 114170 24532 115903
rect 24492 114164 24544 114170
rect 24492 114106 24544 114112
rect 22836 113960 22888 113966
rect 22836 113902 22888 113908
rect 23388 113960 23440 113966
rect 23388 113902 23440 113908
rect 24032 113960 24084 113966
rect 24032 113902 24084 113908
rect 24596 113490 24624 119200
rect 24872 117774 24900 119200
rect 24860 117768 24912 117774
rect 24860 117710 24912 117716
rect 24676 117700 24728 117706
rect 24676 117642 24728 117648
rect 24688 117094 24716 117642
rect 24768 117156 24820 117162
rect 24768 117098 24820 117104
rect 24676 117088 24728 117094
rect 24676 117030 24728 117036
rect 24780 116278 24808 117098
rect 25056 116550 25084 119200
rect 25134 116920 25190 116929
rect 25134 116855 25190 116864
rect 25044 116544 25096 116550
rect 25044 116486 25096 116492
rect 24768 116272 24820 116278
rect 24768 116214 24820 116220
rect 24676 115796 24728 115802
rect 24676 115738 24728 115744
rect 24688 115530 24716 115738
rect 24676 115524 24728 115530
rect 24676 115466 24728 115472
rect 25148 115462 25176 116855
rect 25136 115456 25188 115462
rect 25136 115398 25188 115404
rect 25240 113490 25268 119200
rect 25516 117978 25544 119200
rect 25504 117972 25556 117978
rect 25504 117914 25556 117920
rect 25700 116890 25728 119200
rect 25688 116884 25740 116890
rect 25688 116826 25740 116832
rect 25596 116748 25648 116754
rect 25596 116690 25648 116696
rect 25780 116748 25832 116754
rect 25780 116690 25832 116696
rect 25502 116240 25558 116249
rect 25502 116175 25558 116184
rect 25320 116136 25372 116142
rect 25320 116078 25372 116084
rect 25332 114442 25360 116078
rect 25412 115728 25464 115734
rect 25412 115670 25464 115676
rect 25320 114436 25372 114442
rect 25320 114378 25372 114384
rect 25424 114170 25452 115670
rect 25516 115666 25544 116175
rect 25504 115660 25556 115666
rect 25504 115602 25556 115608
rect 25608 114170 25636 116690
rect 25792 115258 25820 116690
rect 25884 116346 25912 119200
rect 25964 117088 26016 117094
rect 25964 117030 26016 117036
rect 25872 116340 25924 116346
rect 25872 116282 25924 116288
rect 25872 116068 25924 116074
rect 25872 116010 25924 116016
rect 25884 115530 25912 116010
rect 25976 115802 26004 117030
rect 26160 116822 26188 119200
rect 26056 116816 26108 116822
rect 26056 116758 26108 116764
rect 26148 116816 26200 116822
rect 26148 116758 26200 116764
rect 25964 115796 26016 115802
rect 25964 115738 26016 115744
rect 25872 115524 25924 115530
rect 25872 115466 25924 115472
rect 25780 115252 25832 115258
rect 25780 115194 25832 115200
rect 26068 114918 26096 116758
rect 26240 116204 26292 116210
rect 26240 116146 26292 116152
rect 26148 116068 26200 116074
rect 26148 116010 26200 116016
rect 26160 115433 26188 116010
rect 26146 115424 26202 115433
rect 26146 115359 26202 115368
rect 26056 114912 26108 114918
rect 26056 114854 26108 114860
rect 25412 114164 25464 114170
rect 25412 114106 25464 114112
rect 25596 114164 25648 114170
rect 25596 114106 25648 114112
rect 26160 113966 26188 115359
rect 26252 114442 26280 116146
rect 26344 115802 26372 119200
rect 26528 116872 26556 119200
rect 26700 117224 26752 117230
rect 26700 117166 26752 117172
rect 26528 116844 26648 116872
rect 26516 116748 26568 116754
rect 26516 116690 26568 116696
rect 26332 115796 26384 115802
rect 26332 115738 26384 115744
rect 26424 115660 26476 115666
rect 26424 115602 26476 115608
rect 26436 115569 26464 115602
rect 26422 115560 26478 115569
rect 26422 115495 26478 115504
rect 26528 115258 26556 116690
rect 26620 116346 26648 116844
rect 26608 116340 26660 116346
rect 26608 116282 26660 116288
rect 26712 116278 26740 117166
rect 26804 116890 26832 119200
rect 26792 116884 26844 116890
rect 26792 116826 26844 116832
rect 26988 116278 27016 119200
rect 27172 117314 27200 119200
rect 27252 117632 27304 117638
rect 27252 117574 27304 117580
rect 27264 117434 27292 117574
rect 27252 117428 27304 117434
rect 27252 117370 27304 117376
rect 27172 117286 27292 117314
rect 27160 117156 27212 117162
rect 27160 117098 27212 117104
rect 27172 117065 27200 117098
rect 27158 117056 27214 117065
rect 27158 116991 27214 117000
rect 26700 116272 26752 116278
rect 26700 116214 26752 116220
rect 26976 116272 27028 116278
rect 26976 116214 27028 116220
rect 27264 115802 27292 117286
rect 27356 116006 27384 119200
rect 27528 116068 27580 116074
rect 27528 116010 27580 116016
rect 27344 116000 27396 116006
rect 27344 115942 27396 115948
rect 27252 115796 27304 115802
rect 27252 115738 27304 115744
rect 26516 115252 26568 115258
rect 26516 115194 26568 115200
rect 26424 115184 26476 115190
rect 26424 115126 26476 115132
rect 26436 114578 26464 115126
rect 27540 115122 27568 116010
rect 27632 115258 27660 119200
rect 27620 115252 27672 115258
rect 27620 115194 27672 115200
rect 27528 115116 27580 115122
rect 27528 115058 27580 115064
rect 27816 115054 27844 119200
rect 26700 115048 26752 115054
rect 26700 114990 26752 114996
rect 27804 115048 27856 115054
rect 27804 114990 27856 114996
rect 26424 114572 26476 114578
rect 26424 114514 26476 114520
rect 26712 114442 26740 114990
rect 27712 114980 27764 114986
rect 27712 114922 27764 114928
rect 27724 114617 27752 114922
rect 27896 114912 27948 114918
rect 27896 114854 27948 114860
rect 27908 114714 27936 114854
rect 27896 114708 27948 114714
rect 27896 114650 27948 114656
rect 27710 114608 27766 114617
rect 28000 114578 28028 119200
rect 28276 116770 28304 119200
rect 28356 117156 28408 117162
rect 28356 117098 28408 117104
rect 28368 116929 28396 117098
rect 28354 116920 28410 116929
rect 28354 116855 28410 116864
rect 28276 116742 28396 116770
rect 28172 116340 28224 116346
rect 28172 116282 28224 116288
rect 27710 114543 27766 114552
rect 27988 114572 28040 114578
rect 27988 114514 28040 114520
rect 26240 114436 26292 114442
rect 26240 114378 26292 114384
rect 26700 114436 26752 114442
rect 26700 114378 26752 114384
rect 26148 113960 26200 113966
rect 26148 113902 26200 113908
rect 25412 113824 25464 113830
rect 25412 113766 25464 113772
rect 24584 113484 24636 113490
rect 24584 113426 24636 113432
rect 25228 113484 25280 113490
rect 25228 113426 25280 113432
rect 23572 112464 23624 112470
rect 23572 112406 23624 112412
rect 23296 112192 23348 112198
rect 23296 112134 23348 112140
rect 22560 110084 22612 110090
rect 22560 110026 22612 110032
rect 21928 109006 22048 109034
rect 21640 103828 21692 103834
rect 21640 103770 21692 103776
rect 22020 103514 22048 109006
rect 21928 103486 22048 103514
rect 22296 109006 22508 109034
rect 21824 85672 21876 85678
rect 21824 85614 21876 85620
rect 21732 79280 21784 79286
rect 21732 79222 21784 79228
rect 21640 70440 21692 70446
rect 21640 70382 21692 70388
rect 21548 51604 21600 51610
rect 21548 51546 21600 51552
rect 21548 50856 21600 50862
rect 21548 50798 21600 50804
rect 21560 40458 21588 50798
rect 21548 40452 21600 40458
rect 21548 40394 21600 40400
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21456 36236 21508 36242
rect 21456 36178 21508 36184
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 28121 21496 29582
rect 21560 28200 21588 37334
rect 21652 31929 21680 70382
rect 21744 52358 21772 79222
rect 21836 57594 21864 85614
rect 21824 57588 21876 57594
rect 21824 57530 21876 57536
rect 21928 55758 21956 103486
rect 22008 98660 22060 98666
rect 22008 98602 22060 98608
rect 22020 68338 22048 98602
rect 22100 82272 22152 82278
rect 22100 82214 22152 82220
rect 22112 79218 22140 82214
rect 22100 79212 22152 79218
rect 22100 79154 22152 79160
rect 22192 74112 22244 74118
rect 22192 74054 22244 74060
rect 22008 68332 22060 68338
rect 22008 68274 22060 68280
rect 22008 63572 22060 63578
rect 22008 63514 22060 63520
rect 21916 55752 21968 55758
rect 21916 55694 21968 55700
rect 21732 52352 21784 52358
rect 21732 52294 21784 52300
rect 21732 52148 21784 52154
rect 21732 52090 21784 52096
rect 21744 45490 21772 52090
rect 21732 45484 21784 45490
rect 21732 45426 21784 45432
rect 21732 45348 21784 45354
rect 21732 45290 21784 45296
rect 21744 37806 21772 45290
rect 21928 42566 21956 55694
rect 22020 43926 22048 63514
rect 22204 55842 22232 74054
rect 22296 57934 22324 109006
rect 22468 106956 22520 106962
rect 22468 106898 22520 106904
rect 22284 57928 22336 57934
rect 22284 57870 22336 57876
rect 22204 55814 22416 55842
rect 22100 55344 22152 55350
rect 22100 55286 22152 55292
rect 22112 48074 22140 55286
rect 22284 55140 22336 55146
rect 22284 55082 22336 55088
rect 22192 51808 22244 51814
rect 22192 51750 22244 51756
rect 22204 49230 22232 51750
rect 22192 49224 22244 49230
rect 22192 49166 22244 49172
rect 22100 48068 22152 48074
rect 22100 48010 22152 48016
rect 22296 48006 22324 55082
rect 22284 48000 22336 48006
rect 22284 47942 22336 47948
rect 22192 44872 22244 44878
rect 22192 44814 22244 44820
rect 22008 43920 22060 43926
rect 22008 43862 22060 43868
rect 21916 42560 21968 42566
rect 21916 42502 21968 42508
rect 22100 41744 22152 41750
rect 22098 41712 22100 41721
rect 22152 41712 22154 41721
rect 22098 41647 22154 41656
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 21732 37800 21784 37806
rect 21732 37742 21784 37748
rect 21732 37256 21784 37262
rect 21732 37198 21784 37204
rect 21744 36786 21772 37198
rect 21732 36780 21784 36786
rect 21732 36722 21784 36728
rect 21638 31920 21694 31929
rect 21638 31855 21694 31864
rect 21732 31204 21784 31210
rect 21732 31146 21784 31152
rect 21640 28212 21692 28218
rect 21560 28172 21640 28200
rect 21640 28154 21692 28160
rect 21454 28112 21510 28121
rect 21454 28047 21510 28056
rect 21456 27940 21508 27946
rect 21456 27882 21508 27888
rect 21468 27334 21496 27882
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21652 27470 21680 27814
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21456 27056 21508 27062
rect 21456 26998 21508 27004
rect 21364 25356 21416 25362
rect 21364 25298 21416 25304
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21272 24744 21324 24750
rect 21376 24732 21404 25298
rect 21468 24857 21496 26998
rect 21454 24848 21510 24857
rect 21560 24834 21588 27066
rect 21652 26518 21680 27270
rect 21744 27062 21772 31146
rect 21732 27056 21784 27062
rect 21836 27033 21864 38830
rect 21916 38820 21968 38826
rect 21968 38780 22048 38808
rect 21916 38762 21968 38768
rect 22020 38418 22048 38780
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 22008 38412 22060 38418
rect 22008 38354 22060 38360
rect 21916 37936 21968 37942
rect 21914 37904 21916 37913
rect 21968 37904 21970 37913
rect 21914 37839 21970 37848
rect 21916 37800 21968 37806
rect 21916 37742 21968 37748
rect 21732 26998 21784 27004
rect 21822 27024 21878 27033
rect 21822 26959 21878 26968
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 21640 26512 21692 26518
rect 21640 26454 21692 26460
rect 21730 26480 21786 26489
rect 21652 25838 21680 26454
rect 21836 26450 21864 26862
rect 21730 26415 21786 26424
rect 21824 26444 21876 26450
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21560 24806 21680 24834
rect 21454 24783 21510 24792
rect 21548 24744 21600 24750
rect 21376 24704 21496 24732
rect 21272 24686 21324 24692
rect 21284 17338 21312 24686
rect 21468 24274 21496 24704
rect 21548 24686 21600 24692
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21376 22098 21404 24142
rect 21468 23662 21496 24210
rect 21560 24206 21588 24686
rect 21652 24342 21680 24806
rect 21640 24336 21692 24342
rect 21640 24278 21692 24284
rect 21548 24200 21600 24206
rect 21744 24154 21772 26415
rect 21824 26386 21876 26392
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21548 24142 21600 24148
rect 21652 24126 21772 24154
rect 21456 23656 21508 23662
rect 21508 23604 21588 23610
rect 21456 23598 21588 23604
rect 21468 23582 21588 23598
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21468 23118 21496 23462
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21468 22574 21496 23054
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21364 22092 21416 22098
rect 21364 22034 21416 22040
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21376 17746 21404 20742
rect 21468 18698 21496 21830
rect 21560 21418 21588 23582
rect 21548 21412 21600 21418
rect 21548 21354 21600 21360
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 21560 18630 21588 20266
rect 21652 18766 21680 24126
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21744 21978 21772 23598
rect 21836 23186 21864 24618
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21744 21950 21864 21978
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21744 21690 21772 21830
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21836 21026 21864 21950
rect 21744 20998 21864 21026
rect 21744 19514 21772 20998
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21548 18624 21600 18630
rect 21468 18572 21548 18578
rect 21468 18566 21600 18572
rect 21468 18550 21588 18566
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21376 16794 21404 17478
rect 21468 16998 21496 18550
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21560 18086 21588 18362
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21560 8974 21588 18022
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21744 17134 21772 17546
rect 21836 17542 21864 20878
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21744 11082 21772 12650
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 20628 3062 20680 3068
rect 21008 3046 21128 3074
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20824 800 20852 2926
rect 21008 2650 21036 3046
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21100 800 21128 2790
rect 21284 2378 21312 6734
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 21376 800 21404 4014
rect 21836 2990 21864 13466
rect 21928 13190 21956 37742
rect 22020 37738 22048 38354
rect 22008 37732 22060 37738
rect 22008 37674 22060 37680
rect 22112 31890 22140 38490
rect 22100 31884 22152 31890
rect 22100 31826 22152 31832
rect 22112 28370 22140 31826
rect 22204 28506 22232 44814
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22296 39522 22324 44270
rect 22388 41070 22416 55814
rect 22480 51610 22508 106898
rect 22468 51604 22520 51610
rect 22468 51546 22520 51552
rect 22572 51066 22600 110026
rect 23112 108384 23164 108390
rect 23112 108326 23164 108332
rect 23124 100570 23152 108326
rect 23308 101658 23336 112134
rect 23296 101652 23348 101658
rect 23296 101594 23348 101600
rect 23112 100564 23164 100570
rect 23112 100506 23164 100512
rect 23388 91860 23440 91866
rect 23388 91802 23440 91808
rect 23400 88942 23428 91802
rect 23388 88936 23440 88942
rect 23388 88878 23440 88884
rect 23400 87378 23428 88878
rect 23388 87372 23440 87378
rect 23388 87314 23440 87320
rect 23400 86766 23428 87314
rect 23388 86760 23440 86766
rect 23388 86702 23440 86708
rect 22744 86692 22796 86698
rect 22744 86634 22796 86640
rect 22756 80054 22784 86634
rect 23400 86290 23428 86702
rect 23388 86284 23440 86290
rect 23388 86226 23440 86232
rect 23296 86080 23348 86086
rect 23296 86022 23348 86028
rect 23308 85134 23336 86022
rect 23400 85202 23428 86226
rect 23388 85196 23440 85202
rect 23388 85138 23440 85144
rect 23296 85128 23348 85134
rect 23296 85070 23348 85076
rect 22664 80026 22784 80054
rect 22560 51060 22612 51066
rect 22560 51002 22612 51008
rect 22468 50992 22520 50998
rect 22468 50934 22520 50940
rect 22480 46918 22508 50934
rect 22468 46912 22520 46918
rect 22468 46854 22520 46860
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22468 40044 22520 40050
rect 22468 39986 22520 39992
rect 22296 39494 22416 39522
rect 22282 38584 22338 38593
rect 22282 38519 22338 38528
rect 22296 38486 22324 38519
rect 22284 38480 22336 38486
rect 22284 38422 22336 38428
rect 22284 38344 22336 38350
rect 22282 38312 22284 38321
rect 22336 38312 22338 38321
rect 22282 38247 22338 38256
rect 22388 37992 22416 39494
rect 22296 37964 22416 37992
rect 22296 37874 22324 37964
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 22480 37806 22508 39986
rect 22560 39364 22612 39370
rect 22560 39306 22612 39312
rect 22572 38418 22600 39306
rect 22560 38412 22612 38418
rect 22560 38354 22612 38360
rect 22376 37800 22428 37806
rect 22282 37768 22338 37777
rect 22376 37742 22428 37748
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22282 37703 22284 37712
rect 22336 37703 22338 37712
rect 22284 37674 22336 37680
rect 22284 36576 22336 36582
rect 22284 36518 22336 36524
rect 22296 36174 22324 36518
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22296 34542 22324 36110
rect 22284 34536 22336 34542
rect 22284 34478 22336 34484
rect 22282 34368 22338 34377
rect 22282 34303 22338 34312
rect 22296 28801 22324 34303
rect 22388 31113 22416 37742
rect 22560 37664 22612 37670
rect 22480 37624 22560 37652
rect 22480 36718 22508 37624
rect 22560 37606 22612 37612
rect 22560 37188 22612 37194
rect 22560 37130 22612 37136
rect 22572 36854 22600 37130
rect 22560 36848 22612 36854
rect 22560 36790 22612 36796
rect 22468 36712 22520 36718
rect 22468 36654 22520 36660
rect 22480 36174 22508 36654
rect 22468 36168 22520 36174
rect 22520 36128 22600 36156
rect 22468 36110 22520 36116
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22374 31104 22430 31113
rect 22374 31039 22430 31048
rect 22376 30116 22428 30122
rect 22376 30058 22428 30064
rect 22282 28792 22338 28801
rect 22388 28762 22416 30058
rect 22480 29102 22508 35090
rect 22572 34678 22600 36128
rect 22560 34672 22612 34678
rect 22560 34614 22612 34620
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 22572 29170 22600 34478
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22468 29096 22520 29102
rect 22572 29073 22600 29106
rect 22468 29038 22520 29044
rect 22558 29064 22614 29073
rect 22558 28999 22614 29008
rect 22468 28960 22520 28966
rect 22466 28928 22468 28937
rect 22520 28928 22522 28937
rect 22466 28863 22522 28872
rect 22664 28762 22692 80026
rect 22928 77444 22980 77450
rect 22928 77386 22980 77392
rect 22744 75880 22796 75886
rect 22744 75822 22796 75828
rect 22756 38554 22784 75822
rect 22836 62416 22888 62422
rect 22836 62358 22888 62364
rect 22848 41274 22876 62358
rect 22836 41268 22888 41274
rect 22836 41210 22888 41216
rect 22836 40520 22888 40526
rect 22836 40462 22888 40468
rect 22848 39098 22876 40462
rect 22836 39092 22888 39098
rect 22836 39034 22888 39040
rect 22834 38992 22890 39001
rect 22834 38927 22890 38936
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22744 38276 22796 38282
rect 22744 38218 22796 38224
rect 22282 28727 22338 28736
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 22558 28656 22614 28665
rect 22558 28591 22560 28600
rect 22612 28591 22614 28600
rect 22560 28562 22612 28568
rect 22468 28552 22520 28558
rect 22204 28478 22324 28506
rect 22468 28494 22520 28500
rect 22112 28342 22232 28370
rect 22098 28248 22154 28257
rect 22098 28183 22100 28192
rect 22152 28183 22154 28192
rect 22100 28154 22152 28160
rect 22006 27840 22062 27849
rect 22006 27775 22062 27784
rect 22020 25129 22048 27775
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22112 26926 22140 27474
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22204 26382 22232 28342
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22192 25764 22244 25770
rect 22192 25706 22244 25712
rect 22204 25498 22232 25706
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22006 25120 22062 25129
rect 22006 25055 22062 25064
rect 22296 24970 22324 28478
rect 22480 27946 22508 28494
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22468 27940 22520 27946
rect 22468 27882 22520 27888
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22388 27674 22416 27814
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22376 26920 22428 26926
rect 22376 26862 22428 26868
rect 22388 26489 22416 26862
rect 22374 26480 22430 26489
rect 22374 26415 22430 26424
rect 22020 24942 22324 24970
rect 22020 24750 22048 24942
rect 22192 24812 22244 24818
rect 22192 24754 22244 24760
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 22008 24200 22060 24206
rect 22006 24168 22008 24177
rect 22060 24168 22062 24177
rect 22006 24103 22062 24112
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 22020 23610 22048 24006
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22112 23610 22140 23734
rect 22020 23582 22140 23610
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22020 16250 22048 23258
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 21146 22140 22918
rect 22204 21486 22232 24754
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 21690 22324 24686
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22296 19334 22324 21626
rect 22204 19306 22324 19334
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 22204 5030 22232 19306
rect 22388 16574 22416 22714
rect 22480 17066 22508 27270
rect 22572 26382 22600 27950
rect 22652 27600 22704 27606
rect 22652 27542 22704 27548
rect 22560 26376 22612 26382
rect 22560 26318 22612 26324
rect 22572 25838 22600 26318
rect 22664 26314 22692 27542
rect 22756 26568 22784 38218
rect 22848 37670 22876 38927
rect 22836 37664 22888 37670
rect 22836 37606 22888 37612
rect 22836 37324 22888 37330
rect 22836 37266 22888 37272
rect 22848 36242 22876 37266
rect 22836 36236 22888 36242
rect 22836 36178 22888 36184
rect 22848 35698 22876 36178
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22836 33040 22888 33046
rect 22834 33008 22836 33017
rect 22888 33008 22890 33017
rect 22834 32943 22890 32952
rect 22836 32292 22888 32298
rect 22836 32234 22888 32240
rect 22848 31890 22876 32234
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22940 29714 22968 77386
rect 23020 76628 23072 76634
rect 23020 76570 23072 76576
rect 23032 50998 23060 76570
rect 23204 69760 23256 69766
rect 23204 69702 23256 69708
rect 23112 62212 23164 62218
rect 23112 62154 23164 62160
rect 23020 50992 23072 50998
rect 23020 50934 23072 50940
rect 23020 50788 23072 50794
rect 23020 50730 23072 50736
rect 23032 44946 23060 50730
rect 23020 44940 23072 44946
rect 23020 44882 23072 44888
rect 23124 41206 23152 62154
rect 23216 51074 23244 69702
rect 23308 59634 23336 85070
rect 23388 61328 23440 61334
rect 23388 61270 23440 61276
rect 23296 59628 23348 59634
rect 23296 59570 23348 59576
rect 23216 51046 23336 51074
rect 23204 49768 23256 49774
rect 23204 49710 23256 49716
rect 23216 47734 23244 49710
rect 23204 47728 23256 47734
rect 23204 47670 23256 47676
rect 23112 41200 23164 41206
rect 23112 41142 23164 41148
rect 23112 41064 23164 41070
rect 23112 41006 23164 41012
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 23032 39001 23060 40462
rect 23018 38992 23074 39001
rect 23018 38927 23074 38936
rect 23020 38888 23072 38894
rect 23020 38830 23072 38836
rect 22928 29708 22980 29714
rect 22928 29650 22980 29656
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22848 27334 22876 28902
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22940 27130 22968 29446
rect 23032 28994 23060 38830
rect 23124 38457 23152 41006
rect 23308 39302 23336 51046
rect 23400 39370 23428 61270
rect 23584 51066 23612 112406
rect 25320 111376 25372 111382
rect 25320 111318 25372 111324
rect 24676 109812 24728 109818
rect 24676 109754 24728 109760
rect 24032 107024 24084 107030
rect 24032 106966 24084 106972
rect 23664 98660 23716 98666
rect 23664 98602 23716 98608
rect 23572 51060 23624 51066
rect 23572 51002 23624 51008
rect 23480 49224 23532 49230
rect 23480 49166 23532 49172
rect 23492 45336 23520 49166
rect 23492 45308 23612 45336
rect 23480 45076 23532 45082
rect 23480 45018 23532 45024
rect 23388 39364 23440 39370
rect 23388 39306 23440 39312
rect 23296 39296 23348 39302
rect 23296 39238 23348 39244
rect 23294 38992 23350 39001
rect 23492 38962 23520 45018
rect 23294 38927 23350 38936
rect 23480 38956 23532 38962
rect 23110 38448 23166 38457
rect 23110 38383 23166 38392
rect 23204 38412 23256 38418
rect 23204 38354 23256 38360
rect 23216 38321 23244 38354
rect 23308 38350 23336 38927
rect 23480 38898 23532 38904
rect 23386 38584 23442 38593
rect 23386 38519 23388 38528
rect 23440 38519 23442 38528
rect 23388 38490 23440 38496
rect 23492 38486 23520 38898
rect 23480 38480 23532 38486
rect 23480 38422 23532 38428
rect 23388 38412 23440 38418
rect 23388 38354 23440 38360
rect 23296 38344 23348 38350
rect 23202 38312 23258 38321
rect 23296 38286 23348 38292
rect 23400 38282 23428 38354
rect 23202 38247 23258 38256
rect 23388 38276 23440 38282
rect 23388 38218 23440 38224
rect 23492 37924 23520 38422
rect 23400 37896 23520 37924
rect 23296 37800 23348 37806
rect 23124 37760 23296 37788
rect 23124 35222 23152 37760
rect 23400 37777 23428 37896
rect 23480 37800 23532 37806
rect 23296 37742 23348 37748
rect 23386 37768 23442 37777
rect 23480 37742 23532 37748
rect 23386 37703 23388 37712
rect 23440 37703 23442 37712
rect 23388 37674 23440 37680
rect 23400 37643 23428 37674
rect 23388 37324 23440 37330
rect 23388 37266 23440 37272
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23216 36650 23244 37130
rect 23400 36802 23428 37266
rect 23492 36922 23520 37742
rect 23584 37262 23612 45308
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23584 37126 23612 37198
rect 23572 37120 23624 37126
rect 23572 37062 23624 37068
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23400 36786 23520 36802
rect 23400 36780 23532 36786
rect 23400 36774 23480 36780
rect 23480 36722 23532 36728
rect 23204 36644 23256 36650
rect 23204 36586 23256 36592
rect 23216 35834 23244 36586
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23216 35290 23244 35770
rect 23204 35284 23256 35290
rect 23204 35226 23256 35232
rect 23112 35216 23164 35222
rect 23112 35158 23164 35164
rect 23112 33992 23164 33998
rect 23112 33934 23164 33940
rect 23124 29578 23152 33934
rect 23308 30122 23336 36518
rect 23388 36032 23440 36038
rect 23388 35974 23440 35980
rect 23400 35154 23428 35974
rect 23492 35494 23520 36722
rect 23584 36718 23612 36858
rect 23572 36712 23624 36718
rect 23572 36654 23624 36660
rect 23584 35630 23612 36654
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23386 32056 23442 32065
rect 23386 31991 23442 32000
rect 23400 31958 23428 31991
rect 23388 31952 23440 31958
rect 23388 31894 23440 31900
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23400 30122 23428 30194
rect 23296 30116 23348 30122
rect 23296 30058 23348 30064
rect 23388 30116 23440 30122
rect 23388 30058 23440 30064
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23296 29164 23348 29170
rect 23296 29106 23348 29112
rect 23032 28966 23152 28994
rect 23020 28756 23072 28762
rect 23020 28698 23072 28704
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22756 26540 22968 26568
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22652 26308 22704 26314
rect 22652 26250 22704 26256
rect 22664 26042 22692 26250
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 22756 25922 22784 26386
rect 22664 25894 22784 25922
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22572 25294 22600 25774
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22572 24138 22600 25230
rect 22560 24132 22612 24138
rect 22560 24074 22612 24080
rect 22572 23118 22600 24074
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22572 22098 22600 23054
rect 22560 22092 22612 22098
rect 22664 22094 22692 25894
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22756 24206 22784 24550
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22664 22066 22876 22094
rect 22560 22034 22612 22040
rect 22572 21554 22600 22034
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22572 21010 22600 21082
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22848 20534 22876 22066
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22296 16546 22416 16574
rect 22296 6322 22324 16546
rect 22572 15162 22600 20334
rect 22940 17814 22968 26540
rect 22928 17808 22980 17814
rect 22928 17750 22980 17756
rect 23032 17660 23060 28698
rect 23124 28626 23152 28966
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23112 27940 23164 27946
rect 23112 27882 23164 27888
rect 23124 27577 23152 27882
rect 23110 27568 23166 27577
rect 23110 27503 23166 27512
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23124 22778 23152 24346
rect 23216 24342 23244 25638
rect 23308 25498 23336 29106
rect 23492 29102 23520 35430
rect 23570 31648 23626 31657
rect 23570 31583 23626 31592
rect 23584 31346 23612 31583
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 23400 24970 23428 28698
rect 23584 28665 23612 29582
rect 23570 28656 23626 28665
rect 23570 28591 23626 28600
rect 23572 27396 23624 27402
rect 23572 27338 23624 27344
rect 23480 27056 23532 27062
rect 23480 26998 23532 27004
rect 23308 24942 23428 24970
rect 23204 24336 23256 24342
rect 23204 24278 23256 24284
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23308 22386 23336 24942
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23400 22574 23428 24550
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23216 22358 23336 22386
rect 23216 22234 23244 22358
rect 23294 22264 23350 22273
rect 23204 22228 23256 22234
rect 23294 22199 23350 22208
rect 23204 22170 23256 22176
rect 23204 21888 23256 21894
rect 22940 17632 23060 17660
rect 23124 21836 23204 21842
rect 23124 21830 23256 21836
rect 23124 21814 23244 21830
rect 22940 16794 22968 17632
rect 23020 17060 23072 17066
rect 23020 17002 23072 17008
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 22112 3126 22140 3878
rect 22204 3670 22232 3878
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22192 3528 22244 3534
rect 22190 3496 22192 3505
rect 22244 3496 22246 3505
rect 22190 3431 22246 3440
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 21652 800 21680 2450
rect 22020 800 22048 2790
rect 22112 2650 22140 2858
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22296 800 22324 4626
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22388 3058 22416 4218
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22480 2938 22508 7482
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22560 4480 22612 4486
rect 22560 4422 22612 4428
rect 22572 3058 22600 4422
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22388 2922 22508 2938
rect 22376 2916 22508 2922
rect 22428 2910 22508 2916
rect 22376 2858 22428 2864
rect 22664 2774 22692 4558
rect 22848 3482 22876 8978
rect 22940 3602 22968 9658
rect 23032 9042 23060 17002
rect 23124 10606 23152 21814
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23216 10470 23244 20538
rect 23308 19174 23336 22199
rect 23492 21894 23520 26998
rect 23584 25430 23612 27338
rect 23572 25424 23624 25430
rect 23572 25366 23624 25372
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23584 24070 23612 24890
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 23308 9738 23336 19110
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23216 9710 23336 9738
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 23124 5642 23152 9522
rect 23216 7818 23244 9710
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23204 7812 23256 7818
rect 23204 7754 23256 7760
rect 23308 7206 23336 9590
rect 23400 9110 23428 17138
rect 23492 15094 23520 20946
rect 23584 19310 23612 22374
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23480 15088 23532 15094
rect 23480 15030 23532 15036
rect 23388 9104 23440 9110
rect 23388 9046 23440 9052
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23112 5636 23164 5642
rect 23112 5578 23164 5584
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22848 3454 22968 3482
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22572 2746 22692 2774
rect 22572 800 22600 2746
rect 22848 800 22876 3334
rect 22940 2854 22968 3454
rect 22928 2848 22980 2854
rect 22928 2790 22980 2796
rect 23124 800 23152 3946
rect 23308 3738 23336 4014
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23400 3534 23428 3878
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23676 2582 23704 98602
rect 23940 95328 23992 95334
rect 23940 95270 23992 95276
rect 23848 81796 23900 81802
rect 23848 81738 23900 81744
rect 23756 77512 23808 77518
rect 23756 77454 23808 77460
rect 23768 21078 23796 77454
rect 23860 25786 23888 81738
rect 23952 30666 23980 95270
rect 24044 44946 24072 106966
rect 24124 90228 24176 90234
rect 24124 90170 24176 90176
rect 24136 88058 24164 90170
rect 24124 88052 24176 88058
rect 24124 87994 24176 88000
rect 24584 81252 24636 81258
rect 24584 81194 24636 81200
rect 24124 80368 24176 80374
rect 24124 80310 24176 80316
rect 24032 44940 24084 44946
rect 24032 44882 24084 44888
rect 24032 39364 24084 39370
rect 24032 39306 24084 39312
rect 24044 38962 24072 39306
rect 24032 38956 24084 38962
rect 24032 38898 24084 38904
rect 24032 38752 24084 38758
rect 24032 38694 24084 38700
rect 24044 37398 24072 38694
rect 24032 37392 24084 37398
rect 24032 37334 24084 37340
rect 24044 32502 24072 37334
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 23940 30660 23992 30666
rect 23940 30602 23992 30608
rect 23940 30252 23992 30258
rect 23940 30194 23992 30200
rect 23952 29850 23980 30194
rect 23940 29844 23992 29850
rect 23940 29786 23992 29792
rect 24044 29714 24072 32438
rect 24032 29708 24084 29714
rect 24032 29650 24084 29656
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23952 29238 23980 29446
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 24044 28966 24072 29650
rect 24032 28960 24084 28966
rect 24032 28902 24084 28908
rect 24136 28234 24164 80310
rect 24216 78192 24268 78198
rect 24216 78134 24268 78140
rect 24228 53174 24256 78134
rect 24596 62830 24624 81194
rect 24688 67634 24716 109754
rect 24860 105256 24912 105262
rect 24860 105198 24912 105204
rect 24872 104786 24900 105198
rect 24860 104780 24912 104786
rect 24860 104722 24912 104728
rect 24872 103766 24900 104722
rect 24952 104236 25004 104242
rect 24952 104178 25004 104184
rect 24860 103760 24912 103766
rect 24860 103702 24912 103708
rect 24860 93152 24912 93158
rect 24860 93094 24912 93100
rect 24872 86834 24900 93094
rect 24860 86828 24912 86834
rect 24860 86770 24912 86776
rect 24860 76900 24912 76906
rect 24860 76842 24912 76848
rect 24872 76498 24900 76842
rect 24860 76492 24912 76498
rect 24860 76434 24912 76440
rect 24872 75886 24900 76434
rect 24860 75880 24912 75886
rect 24860 75822 24912 75828
rect 24688 67606 24808 67634
rect 24780 62914 24808 67606
rect 24688 62886 24808 62914
rect 24584 62824 24636 62830
rect 24584 62766 24636 62772
rect 24308 62348 24360 62354
rect 24308 62290 24360 62296
rect 24216 53168 24268 53174
rect 24216 53110 24268 53116
rect 24320 40662 24348 62290
rect 24400 60580 24452 60586
rect 24400 60522 24452 60528
rect 24412 45082 24440 60522
rect 24492 59424 24544 59430
rect 24492 59366 24544 59372
rect 24504 49434 24532 59366
rect 24584 54528 24636 54534
rect 24584 54470 24636 54476
rect 24492 49428 24544 49434
rect 24492 49370 24544 49376
rect 24400 45076 24452 45082
rect 24400 45018 24452 45024
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 24308 40656 24360 40662
rect 24308 40598 24360 40604
rect 24320 38894 24348 40598
rect 24308 38888 24360 38894
rect 24308 38830 24360 38836
rect 24400 38820 24452 38826
rect 24400 38762 24452 38768
rect 24216 37936 24268 37942
rect 24214 37904 24216 37913
rect 24268 37904 24270 37913
rect 24214 37839 24270 37848
rect 24412 37806 24440 38762
rect 24504 38418 24532 44814
rect 24492 38412 24544 38418
rect 24492 38354 24544 38360
rect 24400 37800 24452 37806
rect 24400 37742 24452 37748
rect 24490 37768 24546 37777
rect 24490 37703 24546 37712
rect 24216 37664 24268 37670
rect 24216 37606 24268 37612
rect 24228 36242 24256 37606
rect 24308 37392 24360 37398
rect 24308 37334 24360 37340
rect 24216 36236 24268 36242
rect 24216 36178 24268 36184
rect 24320 35562 24348 37334
rect 24400 36780 24452 36786
rect 24400 36722 24452 36728
rect 24412 36038 24440 36722
rect 24400 36032 24452 36038
rect 24400 35974 24452 35980
rect 24308 35556 24360 35562
rect 24308 35498 24360 35504
rect 24216 34672 24268 34678
rect 24216 34614 24268 34620
rect 24228 29714 24256 34614
rect 24398 34504 24454 34513
rect 24398 34439 24454 34448
rect 24306 32328 24362 32337
rect 24306 32263 24308 32272
rect 24360 32263 24362 32272
rect 24308 32234 24360 32240
rect 24412 30258 24440 34439
rect 24400 30252 24452 30258
rect 24400 30194 24452 30200
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 24216 29096 24268 29102
rect 24216 29038 24268 29044
rect 24228 28966 24256 29038
rect 24216 28960 24268 28966
rect 24216 28902 24268 28908
rect 24228 28422 24256 28902
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24044 28206 24164 28234
rect 23938 27568 23994 27577
rect 23938 27503 23994 27512
rect 23952 27334 23980 27503
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23860 25758 23980 25786
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23860 23526 23888 24686
rect 23848 23520 23900 23526
rect 23848 23462 23900 23468
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 23860 22386 23888 23258
rect 23952 22778 23980 25758
rect 24044 24818 24072 28206
rect 24214 27704 24270 27713
rect 24214 27639 24270 27648
rect 24228 27606 24256 27639
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 26586 24164 27270
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24124 26580 24176 26586
rect 24124 26522 24176 26528
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 24136 25702 24164 25978
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 23940 22772 23992 22778
rect 23940 22714 23992 22720
rect 24044 22522 24072 24142
rect 24136 23254 24164 25094
rect 24124 23248 24176 23254
rect 24124 23190 24176 23196
rect 24228 22574 24256 26726
rect 24320 26042 24348 29174
rect 24504 28937 24532 37703
rect 24596 29170 24624 54470
rect 24688 40594 24716 62886
rect 24768 62824 24820 62830
rect 24768 62766 24820 62772
rect 24676 40588 24728 40594
rect 24676 40530 24728 40536
rect 24676 37664 24728 37670
rect 24676 37606 24728 37612
rect 24688 37466 24716 37606
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24676 36100 24728 36106
rect 24676 36042 24728 36048
rect 24688 33998 24716 36042
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24676 33108 24728 33114
rect 24676 33050 24728 33056
rect 24688 31890 24716 33050
rect 24676 31884 24728 31890
rect 24676 31826 24728 31832
rect 24676 30660 24728 30666
rect 24676 30602 24728 30608
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24490 28928 24546 28937
rect 24490 28863 24546 28872
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24412 26450 24440 28086
rect 24688 27946 24716 30602
rect 24676 27940 24728 27946
rect 24676 27882 24728 27888
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24400 26444 24452 26450
rect 24400 26386 24452 26392
rect 24308 26036 24360 26042
rect 24308 25978 24360 25984
rect 24320 24206 24348 25978
rect 24504 25498 24532 27542
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24400 25424 24452 25430
rect 24400 25366 24452 25372
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24216 22568 24268 22574
rect 24044 22494 24164 22522
rect 24216 22510 24268 22516
rect 24032 22432 24084 22438
rect 23860 22358 23980 22386
rect 24032 22374 24084 22380
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23860 21486 23888 22170
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 18426 23888 20878
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 23952 7886 23980 22358
rect 24044 16182 24072 22374
rect 24136 22094 24164 22494
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 24228 22273 24256 22374
rect 24214 22264 24270 22273
rect 24214 22199 24270 22208
rect 24136 22066 24256 22094
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24136 20398 24164 21014
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 24228 5574 24256 22066
rect 24320 17746 24348 23462
rect 24412 23322 24440 25366
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24412 22166 24440 22510
rect 24504 22234 24532 25162
rect 24596 22982 24624 27406
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24688 26926 24716 27270
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24688 23662 24716 24210
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 24412 21078 24440 22102
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24400 21072 24452 21078
rect 24400 21014 24452 21020
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24412 18222 24440 20742
rect 24504 19242 24532 21830
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 24492 19236 24544 19242
rect 24492 19178 24544 19184
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23768 3482 23796 3538
rect 23768 3454 23888 3482
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 23492 800 23520 2450
rect 23768 800 23796 3334
rect 23860 3126 23888 3454
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23952 2990 23980 4150
rect 24320 3670 24348 16594
rect 24596 15434 24624 20946
rect 24688 15706 24716 22034
rect 24780 21010 24808 62766
rect 24964 51610 24992 104178
rect 25044 91316 25096 91322
rect 25044 91258 25096 91264
rect 25056 84658 25084 91258
rect 25044 84652 25096 84658
rect 25044 84594 25096 84600
rect 25136 83700 25188 83706
rect 25136 83642 25188 83648
rect 25044 79144 25096 79150
rect 25044 79086 25096 79092
rect 24952 51604 25004 51610
rect 24952 51546 25004 51552
rect 24860 50992 24912 50998
rect 24860 50934 24912 50940
rect 24872 40730 24900 50934
rect 24860 40724 24912 40730
rect 24860 40666 24912 40672
rect 24872 37738 24900 40666
rect 24860 37732 24912 37738
rect 24860 37674 24912 37680
rect 24952 33856 25004 33862
rect 24952 33798 25004 33804
rect 24860 32972 24912 32978
rect 24860 32914 24912 32920
rect 24872 31770 24900 32914
rect 24964 31958 24992 33798
rect 24952 31952 25004 31958
rect 24952 31894 25004 31900
rect 24872 31742 24992 31770
rect 25056 31754 25084 79086
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24964 31634 24992 31742
rect 25044 31748 25096 31754
rect 25044 31690 25096 31696
rect 24872 25945 24900 31622
rect 24964 31606 25084 31634
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24964 30938 24992 31078
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24964 26858 24992 30874
rect 25056 30870 25084 31606
rect 25044 30864 25096 30870
rect 25044 30806 25096 30812
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25056 30190 25084 30670
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 25056 28626 25084 30126
rect 25044 28620 25096 28626
rect 25044 28562 25096 28568
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 25056 27334 25084 28426
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 24952 26852 25004 26858
rect 24952 26794 25004 26800
rect 25056 26602 25084 27270
rect 24964 26574 25084 26602
rect 24858 25936 24914 25945
rect 24858 25871 24914 25880
rect 24964 23905 24992 26574
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 25056 25906 25084 26318
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 25044 25492 25096 25498
rect 25044 25434 25096 25440
rect 25056 25226 25084 25434
rect 25148 25362 25176 83642
rect 25228 57860 25280 57866
rect 25228 57802 25280 57808
rect 25240 48278 25268 57802
rect 25332 50522 25360 111318
rect 25424 51066 25452 113766
rect 28184 112878 28212 116282
rect 28264 116068 28316 116074
rect 28264 116010 28316 116016
rect 28276 115977 28304 116010
rect 28262 115968 28318 115977
rect 28262 115903 28318 115912
rect 28368 115122 28396 116742
rect 28356 115116 28408 115122
rect 28356 115058 28408 115064
rect 28460 114578 28488 119200
rect 28540 116816 28592 116822
rect 28540 116758 28592 116764
rect 28448 114572 28500 114578
rect 28448 114514 28500 114520
rect 28552 113014 28580 116758
rect 28644 114646 28672 119200
rect 28816 116612 28868 116618
rect 28816 116554 28868 116560
rect 28828 116210 28856 116554
rect 28816 116204 28868 116210
rect 28816 116146 28868 116152
rect 28724 115660 28776 115666
rect 28724 115602 28776 115608
rect 28816 115660 28868 115666
rect 28816 115602 28868 115608
rect 28632 114640 28684 114646
rect 28632 114582 28684 114588
rect 28632 114368 28684 114374
rect 28632 114310 28684 114316
rect 28644 113966 28672 114310
rect 28736 114170 28764 115602
rect 28828 115297 28856 115602
rect 28814 115288 28870 115297
rect 28920 115258 28948 119200
rect 29104 116890 29132 119200
rect 29184 117088 29236 117094
rect 29184 117030 29236 117036
rect 29092 116884 29144 116890
rect 29092 116826 29144 116832
rect 29000 116068 29052 116074
rect 29000 116010 29052 116016
rect 28814 115223 28870 115232
rect 28908 115252 28960 115258
rect 28908 115194 28960 115200
rect 29012 115161 29040 116010
rect 29196 115462 29224 117030
rect 29184 115456 29236 115462
rect 29184 115398 29236 115404
rect 28998 115152 29054 115161
rect 28998 115087 29054 115096
rect 29092 114980 29144 114986
rect 29092 114922 29144 114928
rect 29104 114714 29132 114922
rect 29092 114708 29144 114714
rect 29092 114650 29144 114656
rect 28724 114164 28776 114170
rect 28724 114106 28776 114112
rect 29288 113966 29316 119200
rect 29368 116544 29420 116550
rect 29368 116486 29420 116492
rect 29380 114102 29408 116486
rect 29472 115802 29500 119200
rect 29644 116680 29696 116686
rect 29644 116622 29696 116628
rect 29552 116544 29604 116550
rect 29552 116486 29604 116492
rect 29460 115796 29512 115802
rect 29460 115738 29512 115744
rect 29564 114714 29592 116486
rect 29552 114708 29604 114714
rect 29552 114650 29604 114656
rect 29656 114170 29684 116622
rect 29748 115802 29776 119200
rect 29828 117768 29880 117774
rect 29828 117710 29880 117716
rect 29840 117434 29868 117710
rect 29828 117428 29880 117434
rect 29828 117370 29880 117376
rect 29828 116000 29880 116006
rect 29828 115942 29880 115948
rect 29736 115796 29788 115802
rect 29736 115738 29788 115744
rect 29736 115456 29788 115462
rect 29736 115398 29788 115404
rect 29644 114164 29696 114170
rect 29644 114106 29696 114112
rect 29368 114096 29420 114102
rect 29368 114038 29420 114044
rect 28632 113960 28684 113966
rect 28632 113902 28684 113908
rect 29276 113960 29328 113966
rect 29276 113902 29328 113908
rect 28540 113008 28592 113014
rect 28540 112950 28592 112956
rect 28172 112872 28224 112878
rect 28172 112814 28224 112820
rect 26240 112736 26292 112742
rect 26240 112678 26292 112684
rect 26252 109750 26280 112678
rect 26792 111172 26844 111178
rect 26792 111114 26844 111120
rect 26700 110016 26752 110022
rect 26700 109958 26752 109964
rect 26240 109744 26292 109750
rect 26240 109686 26292 109692
rect 25964 105732 26016 105738
rect 25964 105674 26016 105680
rect 25976 104922 26004 105674
rect 26056 105256 26108 105262
rect 26056 105198 26108 105204
rect 25964 104916 26016 104922
rect 25964 104858 26016 104864
rect 26068 104854 26096 105198
rect 26056 104848 26108 104854
rect 26056 104790 26108 104796
rect 26712 103514 26740 109958
rect 26804 103766 26832 111114
rect 28264 110900 28316 110906
rect 28264 110842 28316 110848
rect 27620 109744 27672 109750
rect 27620 109686 27672 109692
rect 27632 105466 27660 109686
rect 27620 105460 27672 105466
rect 27620 105402 27672 105408
rect 26884 104168 26936 104174
rect 26884 104110 26936 104116
rect 26792 103760 26844 103766
rect 26792 103702 26844 103708
rect 26712 103486 26832 103514
rect 26804 102746 26832 103486
rect 26792 102740 26844 102746
rect 26792 102682 26844 102688
rect 26700 102604 26752 102610
rect 26700 102546 26752 102552
rect 26712 98734 26740 102546
rect 26700 98728 26752 98734
rect 26700 98670 26752 98676
rect 25504 94784 25556 94790
rect 25504 94726 25556 94732
rect 25516 86358 25544 94726
rect 26896 91798 26924 104110
rect 28276 98870 28304 110842
rect 29644 106412 29696 106418
rect 29644 106354 29696 106360
rect 29656 99822 29684 106354
rect 29644 99816 29696 99822
rect 29644 99758 29696 99764
rect 29656 99414 29684 99758
rect 29644 99408 29696 99414
rect 29644 99350 29696 99356
rect 28264 98864 28316 98870
rect 28264 98806 28316 98812
rect 29460 98048 29512 98054
rect 29460 97990 29512 97996
rect 28908 96416 28960 96422
rect 28908 96358 28960 96364
rect 28448 95940 28500 95946
rect 28448 95882 28500 95888
rect 27068 95872 27120 95878
rect 27068 95814 27120 95820
rect 26976 93900 27028 93906
rect 26976 93842 27028 93848
rect 26884 91792 26936 91798
rect 26884 91734 26936 91740
rect 26792 90636 26844 90642
rect 26792 90578 26844 90584
rect 26240 87848 26292 87854
rect 26240 87790 26292 87796
rect 26148 87508 26200 87514
rect 26148 87450 26200 87456
rect 25504 86352 25556 86358
rect 25504 86294 25556 86300
rect 25872 85060 25924 85066
rect 25872 85002 25924 85008
rect 25502 81696 25558 81705
rect 25502 81631 25558 81640
rect 25516 79626 25544 81631
rect 25780 80844 25832 80850
rect 25780 80786 25832 80792
rect 25688 80232 25740 80238
rect 25688 80174 25740 80180
rect 25596 79756 25648 79762
rect 25596 79698 25648 79704
rect 25504 79620 25556 79626
rect 25504 79562 25556 79568
rect 25502 79520 25558 79529
rect 25502 79455 25558 79464
rect 25516 79354 25544 79455
rect 25504 79348 25556 79354
rect 25504 79290 25556 79296
rect 25608 78470 25636 79698
rect 25596 78464 25648 78470
rect 25596 78406 25648 78412
rect 25504 77920 25556 77926
rect 25504 77862 25556 77868
rect 25412 51060 25464 51066
rect 25412 51002 25464 51008
rect 25320 50516 25372 50522
rect 25320 50458 25372 50464
rect 25228 48272 25280 48278
rect 25228 48214 25280 48220
rect 25412 39092 25464 39098
rect 25412 39034 25464 39040
rect 25228 38888 25280 38894
rect 25228 38830 25280 38836
rect 25240 38214 25268 38830
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38486 25360 38694
rect 25320 38480 25372 38486
rect 25320 38422 25372 38428
rect 25228 38208 25280 38214
rect 25228 38150 25280 38156
rect 25320 38208 25372 38214
rect 25320 38150 25372 38156
rect 25240 36922 25268 38150
rect 25332 37874 25360 38150
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 25424 34184 25452 39034
rect 25516 38894 25544 77862
rect 25596 57384 25648 57390
rect 25596 57326 25648 57332
rect 25608 57089 25636 57326
rect 25594 57080 25650 57089
rect 25594 57015 25650 57024
rect 25596 54120 25648 54126
rect 25596 54062 25648 54068
rect 25504 38888 25556 38894
rect 25504 38830 25556 38836
rect 25504 38752 25556 38758
rect 25504 38694 25556 38700
rect 25332 34156 25452 34184
rect 25332 33318 25360 34156
rect 25412 34060 25464 34066
rect 25412 34002 25464 34008
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25332 32978 25360 33254
rect 25320 32972 25372 32978
rect 25320 32914 25372 32920
rect 25228 32496 25280 32502
rect 25226 32464 25228 32473
rect 25280 32464 25282 32473
rect 25226 32399 25282 32408
rect 25332 32366 25360 32914
rect 25320 32360 25372 32366
rect 25240 32320 25320 32348
rect 25240 31686 25268 32320
rect 25424 32337 25452 34002
rect 25516 33386 25544 38694
rect 25504 33380 25556 33386
rect 25504 33322 25556 33328
rect 25516 32842 25544 33322
rect 25504 32836 25556 32842
rect 25504 32778 25556 32784
rect 25516 32502 25544 32778
rect 25504 32496 25556 32502
rect 25504 32438 25556 32444
rect 25320 32302 25372 32308
rect 25410 32328 25466 32337
rect 25410 32263 25466 32272
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25228 31680 25280 31686
rect 25228 31622 25280 31628
rect 25332 31328 25360 32166
rect 25240 31300 25360 31328
rect 25240 29782 25268 31300
rect 25320 31204 25372 31210
rect 25424 31192 25452 32263
rect 25516 31958 25544 32438
rect 25504 31952 25556 31958
rect 25504 31894 25556 31900
rect 25516 31822 25544 31894
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25372 31164 25452 31192
rect 25320 31146 25372 31152
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25412 30864 25464 30870
rect 25412 30806 25464 30812
rect 25320 30116 25372 30122
rect 25320 30058 25372 30064
rect 25228 29776 25280 29782
rect 25228 29718 25280 29724
rect 25226 29064 25282 29073
rect 25332 29034 25360 30058
rect 25226 28999 25282 29008
rect 25320 29028 25372 29034
rect 25240 27130 25268 28999
rect 25320 28970 25372 28976
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25228 27124 25280 27130
rect 25228 27066 25280 27072
rect 25332 26858 25360 27270
rect 25320 26852 25372 26858
rect 25320 26794 25372 26800
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 24950 23896 25006 23905
rect 24950 23831 25006 23840
rect 25056 23526 25084 24754
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24964 18970 24992 21966
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 25148 18902 25176 25162
rect 25240 21894 25268 26726
rect 25424 25650 25452 30806
rect 25516 25838 25544 31078
rect 25608 26994 25636 54062
rect 25700 32842 25728 80174
rect 25792 33658 25820 80786
rect 25884 80782 25912 85002
rect 25962 84280 26018 84289
rect 25962 84215 26018 84224
rect 25872 80776 25924 80782
rect 25872 80718 25924 80724
rect 25884 80102 25912 80718
rect 25872 80096 25924 80102
rect 25872 80038 25924 80044
rect 25884 79082 25912 80038
rect 25872 79076 25924 79082
rect 25872 79018 25924 79024
rect 25872 60512 25924 60518
rect 25872 60454 25924 60460
rect 25884 49298 25912 60454
rect 25872 49292 25924 49298
rect 25872 49234 25924 49240
rect 25872 43104 25924 43110
rect 25872 43046 25924 43052
rect 25884 42838 25912 43046
rect 25872 42832 25924 42838
rect 25872 42774 25924 42780
rect 25884 41750 25912 42774
rect 25872 41744 25924 41750
rect 25872 41686 25924 41692
rect 25872 38412 25924 38418
rect 25872 38354 25924 38360
rect 25884 38321 25912 38354
rect 25870 38312 25926 38321
rect 25870 38247 25926 38256
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25884 34406 25912 34954
rect 25872 34400 25924 34406
rect 25872 34342 25924 34348
rect 25780 33652 25832 33658
rect 25780 33594 25832 33600
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25688 32836 25740 32842
rect 25688 32778 25740 32784
rect 25688 32496 25740 32502
rect 25688 32438 25740 32444
rect 25700 32298 25728 32438
rect 25688 32292 25740 32298
rect 25688 32234 25740 32240
rect 25688 32020 25740 32026
rect 25688 31962 25740 31968
rect 25700 29578 25728 31962
rect 25688 29572 25740 29578
rect 25688 29514 25740 29520
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25424 25622 25544 25650
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 25424 23798 25452 24686
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 25516 23254 25544 25622
rect 25504 23248 25556 23254
rect 25504 23190 25556 23196
rect 25228 21888 25280 21894
rect 25228 21830 25280 21836
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25412 18148 25464 18154
rect 25412 18090 25464 18096
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24952 15020 25004 15026
rect 24952 14962 25004 14968
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24768 11008 24820 11014
rect 24768 10950 24820 10956
rect 24780 8430 24808 10950
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24872 7818 24900 14418
rect 24964 9926 24992 14962
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 24400 3664 24452 3670
rect 24400 3606 24452 3612
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24044 800 24072 3538
rect 24412 3505 24440 3606
rect 24398 3496 24454 3505
rect 24398 3431 24454 3440
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24504 3194 24532 3334
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 24308 2508 24360 2514
rect 24308 2450 24360 2456
rect 24320 800 24348 2450
rect 24596 800 24624 2790
rect 24872 800 24900 4014
rect 25148 2774 25176 4626
rect 25228 4480 25280 4486
rect 25228 4422 25280 4428
rect 25240 4282 25268 4422
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 25240 3126 25268 3878
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 25332 2990 25360 18022
rect 25424 3670 25452 18090
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25412 3664 25464 3670
rect 25412 3606 25464 3612
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 25320 2984 25372 2990
rect 25320 2926 25372 2932
rect 25148 2746 25268 2774
rect 25240 800 25268 2746
rect 25516 800 25544 3334
rect 25608 2854 25636 8978
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 25700 2582 25728 29514
rect 25792 29322 25820 33458
rect 25884 33454 25912 34342
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25884 30802 25912 33390
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 25792 29294 25912 29322
rect 25780 27872 25832 27878
rect 25780 27814 25832 27820
rect 25792 26518 25820 27814
rect 25884 27418 25912 29294
rect 25976 27538 26004 84215
rect 26054 79928 26110 79937
rect 26054 79863 26110 79872
rect 26068 79694 26096 79863
rect 26056 79688 26108 79694
rect 26056 79630 26108 79636
rect 26056 79552 26108 79558
rect 26056 79494 26108 79500
rect 26068 32570 26096 79494
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26054 32464 26110 32473
rect 26054 32399 26110 32408
rect 26068 32026 26096 32399
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 26056 31884 26108 31890
rect 26056 31826 26108 31832
rect 25964 27532 26016 27538
rect 25964 27474 26016 27480
rect 25884 27390 26004 27418
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25780 26512 25832 26518
rect 25780 26454 25832 26460
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25792 24410 25820 24686
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25884 14482 25912 27066
rect 25976 26858 26004 27390
rect 26068 26908 26096 31826
rect 26160 28082 26188 87450
rect 26252 59650 26280 87790
rect 26608 86760 26660 86766
rect 26608 86702 26660 86708
rect 26332 86216 26384 86222
rect 26332 86158 26384 86164
rect 26344 60042 26372 86158
rect 26424 85196 26476 85202
rect 26424 85138 26476 85144
rect 26436 79830 26464 85138
rect 26424 79824 26476 79830
rect 26424 79766 26476 79772
rect 26436 78742 26464 79766
rect 26514 79656 26570 79665
rect 26514 79591 26570 79600
rect 26424 78736 26476 78742
rect 26424 78678 26476 78684
rect 26422 78568 26478 78577
rect 26422 78503 26478 78512
rect 26436 75750 26464 78503
rect 26424 75744 26476 75750
rect 26424 75686 26476 75692
rect 26424 75404 26476 75410
rect 26424 75346 26476 75352
rect 26332 60036 26384 60042
rect 26332 59978 26384 59984
rect 26252 59622 26372 59650
rect 26240 59560 26292 59566
rect 26240 59502 26292 59508
rect 26252 58546 26280 59502
rect 26240 58540 26292 58546
rect 26240 58482 26292 58488
rect 26240 58404 26292 58410
rect 26240 58346 26292 58352
rect 26252 57322 26280 58346
rect 26240 57316 26292 57322
rect 26240 57258 26292 57264
rect 26252 56953 26280 57258
rect 26238 56944 26294 56953
rect 26238 56879 26294 56888
rect 26252 56234 26280 56879
rect 26240 56228 26292 56234
rect 26240 56170 26292 56176
rect 26344 54890 26372 59622
rect 26252 54862 26372 54890
rect 26252 47734 26280 54862
rect 26332 52896 26384 52902
rect 26332 52838 26384 52844
rect 26344 51882 26372 52838
rect 26332 51876 26384 51882
rect 26332 51818 26384 51824
rect 26344 50794 26372 51818
rect 26332 50788 26384 50794
rect 26332 50730 26384 50736
rect 26240 47728 26292 47734
rect 26436 47682 26464 75346
rect 26528 75206 26556 79591
rect 26516 75200 26568 75206
rect 26516 75142 26568 75148
rect 26516 60648 26568 60654
rect 26516 60590 26568 60596
rect 26528 58546 26556 60590
rect 26516 58540 26568 58546
rect 26516 58482 26568 58488
rect 26528 57458 26556 58482
rect 26516 57452 26568 57458
rect 26516 57394 26568 57400
rect 26528 57050 26556 57394
rect 26516 57044 26568 57050
rect 26620 57032 26648 86702
rect 26700 86692 26752 86698
rect 26700 86634 26752 86640
rect 26712 86290 26740 86634
rect 26700 86284 26752 86290
rect 26700 86226 26752 86232
rect 26712 85202 26740 86226
rect 26700 85196 26752 85202
rect 26700 85138 26752 85144
rect 26700 82408 26752 82414
rect 26700 82350 26752 82356
rect 26620 57004 26653 57032
rect 26516 56986 26568 56992
rect 26514 56944 26570 56953
rect 26625 56896 26653 57004
rect 26514 56879 26516 56888
rect 26568 56879 26570 56888
rect 26516 56850 26568 56856
rect 26620 56868 26653 56896
rect 26514 56808 26570 56817
rect 26514 56743 26570 56752
rect 26528 56710 26556 56743
rect 26516 56704 26568 56710
rect 26516 56646 26568 56652
rect 26516 50856 26568 50862
rect 26516 50798 26568 50804
rect 26528 50250 26556 50798
rect 26516 50244 26568 50250
rect 26516 50186 26568 50192
rect 26240 47670 26292 47676
rect 26344 47654 26464 47682
rect 26620 47666 26648 56868
rect 26608 47660 26660 47666
rect 26240 47116 26292 47122
rect 26240 47058 26292 47064
rect 26252 46986 26280 47058
rect 26240 46980 26292 46986
rect 26240 46922 26292 46928
rect 26240 46368 26292 46374
rect 26240 46310 26292 46316
rect 26252 45898 26280 46310
rect 26240 45892 26292 45898
rect 26240 45834 26292 45840
rect 26252 45286 26280 45834
rect 26240 45280 26292 45286
rect 26240 45222 26292 45228
rect 26252 42362 26280 45222
rect 26240 42356 26292 42362
rect 26240 42298 26292 42304
rect 26240 42220 26292 42226
rect 26240 42162 26292 42168
rect 26252 41313 26280 42162
rect 26238 41304 26294 41313
rect 26238 41239 26294 41248
rect 26252 36802 26280 41239
rect 26344 38282 26372 47654
rect 26608 47602 26660 47608
rect 26424 47592 26476 47598
rect 26424 47534 26476 47540
rect 26436 47258 26464 47534
rect 26516 47524 26568 47530
rect 26516 47466 26568 47472
rect 26608 47524 26660 47530
rect 26608 47466 26660 47472
rect 26424 47252 26476 47258
rect 26424 47194 26476 47200
rect 26528 47138 26556 47466
rect 26620 47258 26648 47466
rect 26608 47252 26660 47258
rect 26608 47194 26660 47200
rect 26436 47122 26556 47138
rect 26424 47116 26556 47122
rect 26476 47110 26556 47116
rect 26424 47058 26476 47064
rect 26436 46594 26464 47058
rect 26436 46566 26556 46594
rect 26424 46504 26476 46510
rect 26424 46446 26476 46452
rect 26436 46170 26464 46446
rect 26528 46442 26556 46566
rect 26620 46442 26648 47194
rect 26516 46436 26568 46442
rect 26516 46378 26568 46384
rect 26608 46436 26660 46442
rect 26608 46378 26660 46384
rect 26424 46164 26476 46170
rect 26424 46106 26476 46112
rect 26424 46028 26476 46034
rect 26424 45970 26476 45976
rect 26436 45778 26464 45970
rect 26528 45778 26556 46378
rect 26436 45750 26556 45778
rect 26424 45416 26476 45422
rect 26424 45358 26476 45364
rect 26436 44538 26464 45358
rect 26528 45354 26556 45750
rect 26516 45348 26568 45354
rect 26516 45290 26568 45296
rect 26424 44532 26476 44538
rect 26424 44474 26476 44480
rect 26528 44418 26556 45290
rect 26608 44940 26660 44946
rect 26608 44882 26660 44888
rect 26436 44390 26556 44418
rect 26436 42158 26464 44390
rect 26516 43376 26568 43382
rect 26516 43318 26568 43324
rect 26528 43246 26556 43318
rect 26516 43240 26568 43246
rect 26516 43182 26568 43188
rect 26516 42696 26568 42702
rect 26514 42664 26516 42673
rect 26568 42664 26570 42673
rect 26514 42599 26570 42608
rect 26620 42226 26648 44882
rect 26608 42220 26660 42226
rect 26608 42162 26660 42168
rect 26424 42152 26476 42158
rect 26424 42094 26476 42100
rect 26516 42016 26568 42022
rect 26516 41958 26568 41964
rect 26424 41744 26476 41750
rect 26424 41686 26476 41692
rect 26436 41002 26464 41686
rect 26528 41682 26556 41958
rect 26606 41712 26662 41721
rect 26516 41676 26568 41682
rect 26606 41647 26608 41656
rect 26516 41618 26568 41624
rect 26660 41647 26662 41656
rect 26608 41618 26660 41624
rect 26516 41064 26568 41070
rect 26516 41006 26568 41012
rect 26424 40996 26476 41002
rect 26424 40938 26476 40944
rect 26528 40730 26556 41006
rect 26516 40724 26568 40730
rect 26516 40666 26568 40672
rect 26516 40588 26568 40594
rect 26516 40530 26568 40536
rect 26424 38480 26476 38486
rect 26424 38422 26476 38428
rect 26332 38276 26384 38282
rect 26332 38218 26384 38224
rect 26332 37868 26384 37874
rect 26332 37810 26384 37816
rect 26344 36922 26372 37810
rect 26436 37738 26464 38422
rect 26528 38418 26556 40530
rect 26516 38412 26568 38418
rect 26516 38354 26568 38360
rect 26528 37806 26556 38354
rect 26608 38004 26660 38010
rect 26608 37946 26660 37952
rect 26516 37800 26568 37806
rect 26516 37742 26568 37748
rect 26424 37732 26476 37738
rect 26424 37674 26476 37680
rect 26436 37398 26464 37674
rect 26424 37392 26476 37398
rect 26424 37334 26476 37340
rect 26332 36916 26384 36922
rect 26332 36858 26384 36864
rect 26252 36774 26372 36802
rect 26240 36712 26292 36718
rect 26240 36654 26292 36660
rect 26252 35630 26280 36654
rect 26344 36582 26372 36774
rect 26436 36650 26464 37334
rect 26528 37262 26556 37742
rect 26620 37330 26648 37946
rect 26608 37324 26660 37330
rect 26608 37266 26660 37272
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26528 36718 26556 37198
rect 26712 36922 26740 82350
rect 26804 58138 26832 90578
rect 26988 86086 27016 93842
rect 27080 87854 27108 95814
rect 28264 94784 28316 94790
rect 28264 94726 28316 94732
rect 27344 93288 27396 93294
rect 27344 93230 27396 93236
rect 27356 90710 27384 93230
rect 27344 90704 27396 90710
rect 27344 90646 27396 90652
rect 27804 90024 27856 90030
rect 27804 89966 27856 89972
rect 27816 89714 27844 89966
rect 27816 89686 28028 89714
rect 27712 89548 27764 89554
rect 27712 89490 27764 89496
rect 27160 88868 27212 88874
rect 27160 88810 27212 88816
rect 27068 87848 27120 87854
rect 27068 87790 27120 87796
rect 27172 86766 27200 88810
rect 27436 88460 27488 88466
rect 27436 88402 27488 88408
rect 27252 88324 27304 88330
rect 27252 88266 27304 88272
rect 27264 87786 27292 88266
rect 27252 87780 27304 87786
rect 27252 87722 27304 87728
rect 27160 86760 27212 86766
rect 27160 86702 27212 86708
rect 27172 86193 27200 86702
rect 27264 86222 27292 87722
rect 27344 87372 27396 87378
rect 27344 87314 27396 87320
rect 27252 86216 27304 86222
rect 27158 86184 27214 86193
rect 27252 86158 27304 86164
rect 27158 86119 27214 86128
rect 26976 86080 27028 86086
rect 26976 86022 27028 86028
rect 27264 85338 27292 86158
rect 27252 85332 27304 85338
rect 27252 85274 27304 85280
rect 27160 85196 27212 85202
rect 27160 85138 27212 85144
rect 27068 84584 27120 84590
rect 27068 84526 27120 84532
rect 26884 83496 26936 83502
rect 26884 83438 26936 83444
rect 26896 75410 26924 83438
rect 26976 83020 27028 83026
rect 26976 82962 27028 82968
rect 26884 75404 26936 75410
rect 26884 75346 26936 75352
rect 26988 75290 27016 82962
rect 26896 75262 27016 75290
rect 26792 58132 26844 58138
rect 26792 58074 26844 58080
rect 26896 58018 26924 75262
rect 26976 75200 27028 75206
rect 26976 75142 27028 75148
rect 26804 57990 26924 58018
rect 26804 55842 26832 57990
rect 26884 56976 26936 56982
rect 26884 56918 26936 56924
rect 26896 56370 26924 56918
rect 26884 56364 26936 56370
rect 26884 56306 26936 56312
rect 26884 56228 26936 56234
rect 26884 56170 26936 56176
rect 26896 55962 26924 56170
rect 26884 55956 26936 55962
rect 26884 55898 26936 55904
rect 26804 55814 26924 55842
rect 26792 52964 26844 52970
rect 26792 52906 26844 52912
rect 26804 51950 26832 52906
rect 26792 51944 26844 51950
rect 26792 51886 26844 51892
rect 26804 51542 26832 51886
rect 26792 51536 26844 51542
rect 26792 51478 26844 51484
rect 26804 50794 26832 51478
rect 26792 50788 26844 50794
rect 26792 50730 26844 50736
rect 26804 49706 26832 50730
rect 26792 49700 26844 49706
rect 26792 49642 26844 49648
rect 26804 44538 26832 49642
rect 26792 44532 26844 44538
rect 26792 44474 26844 44480
rect 26792 44260 26844 44266
rect 26792 44202 26844 44208
rect 26804 42294 26832 44202
rect 26792 42288 26844 42294
rect 26792 42230 26844 42236
rect 26792 42016 26844 42022
rect 26792 41958 26844 41964
rect 26804 41002 26832 41958
rect 26792 40996 26844 41002
rect 26792 40938 26844 40944
rect 26792 40112 26844 40118
rect 26792 40054 26844 40060
rect 26804 38010 26832 40054
rect 26792 38004 26844 38010
rect 26792 37946 26844 37952
rect 26896 37330 26924 55814
rect 26884 37324 26936 37330
rect 26884 37266 26936 37272
rect 26884 37188 26936 37194
rect 26884 37130 26936 37136
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 26700 36916 26752 36922
rect 26700 36858 26752 36864
rect 26620 36802 26648 36858
rect 26620 36774 26832 36802
rect 26516 36712 26568 36718
rect 26516 36654 26568 36660
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26424 36644 26476 36650
rect 26424 36586 26476 36592
rect 26332 36576 26384 36582
rect 26332 36518 26384 36524
rect 26332 36236 26384 36242
rect 26436 36224 26464 36586
rect 26528 36242 26556 36654
rect 26620 36378 26648 36654
rect 26700 36576 26752 36582
rect 26700 36518 26752 36524
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26384 36196 26464 36224
rect 26516 36236 26568 36242
rect 26332 36178 26384 36184
rect 26516 36178 26568 36184
rect 26332 35828 26384 35834
rect 26332 35770 26384 35776
rect 26240 35624 26292 35630
rect 26240 35566 26292 35572
rect 26240 35284 26292 35290
rect 26240 35226 26292 35232
rect 26252 31754 26280 35226
rect 26344 32910 26372 35770
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26516 34536 26568 34542
rect 26516 34478 26568 34484
rect 26528 33386 26556 34478
rect 26620 33998 26648 35430
rect 26712 34105 26740 36518
rect 26804 35698 26832 36774
rect 26792 35692 26844 35698
rect 26792 35634 26844 35640
rect 26896 34377 26924 37130
rect 26988 36242 27016 75142
rect 27080 50810 27108 84526
rect 27172 58682 27200 85138
rect 27252 83156 27304 83162
rect 27252 83098 27304 83104
rect 27264 82346 27292 83098
rect 27252 82340 27304 82346
rect 27252 82282 27304 82288
rect 27252 81728 27304 81734
rect 27252 81670 27304 81676
rect 27160 58676 27212 58682
rect 27160 58618 27212 58624
rect 27160 58132 27212 58138
rect 27160 58074 27212 58080
rect 27172 53242 27200 58074
rect 27160 53236 27212 53242
rect 27160 53178 27212 53184
rect 27160 52352 27212 52358
rect 27160 52294 27212 52300
rect 27172 51950 27200 52294
rect 27160 51944 27212 51950
rect 27160 51886 27212 51892
rect 27080 50782 27200 50810
rect 27068 47660 27120 47666
rect 27068 47602 27120 47608
rect 27080 42770 27108 47602
rect 27068 42764 27120 42770
rect 27068 42706 27120 42712
rect 27068 42356 27120 42362
rect 27068 42298 27120 42304
rect 26976 36236 27028 36242
rect 26976 36178 27028 36184
rect 26976 35556 27028 35562
rect 26976 35498 27028 35504
rect 26882 34368 26938 34377
rect 26882 34303 26938 34312
rect 26882 34232 26938 34241
rect 26882 34167 26938 34176
rect 26698 34096 26754 34105
rect 26698 34031 26754 34040
rect 26792 34060 26844 34066
rect 26792 34002 26844 34008
rect 26608 33992 26660 33998
rect 26608 33934 26660 33940
rect 26700 33992 26752 33998
rect 26700 33934 26752 33940
rect 26608 33856 26660 33862
rect 26608 33798 26660 33804
rect 26516 33380 26568 33386
rect 26516 33322 26568 33328
rect 26424 32972 26476 32978
rect 26424 32914 26476 32920
rect 26516 32972 26568 32978
rect 26516 32914 26568 32920
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26240 31748 26292 31754
rect 26240 31690 26292 31696
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26252 30258 26280 30534
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 26344 30190 26372 32710
rect 26436 30666 26464 32914
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26424 30320 26476 30326
rect 26528 30308 26556 32914
rect 26620 30870 26648 33798
rect 26608 30864 26660 30870
rect 26608 30806 26660 30812
rect 26608 30660 26660 30666
rect 26608 30602 26660 30608
rect 26476 30280 26556 30308
rect 26424 30262 26476 30268
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 26332 29708 26384 29714
rect 26332 29650 26384 29656
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 26148 28076 26200 28082
rect 26148 28018 26200 28024
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26160 27606 26188 27814
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27334 26188 27406
rect 26148 27328 26200 27334
rect 26148 27270 26200 27276
rect 26068 26880 26188 26908
rect 25964 26852 26016 26858
rect 25964 26794 26016 26800
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 25976 21418 26004 25230
rect 25964 21412 26016 21418
rect 25964 21354 26016 21360
rect 26068 18222 26096 25298
rect 26160 24834 26188 26880
rect 26252 26450 26280 29446
rect 26344 28762 26372 29650
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26344 27538 26372 27950
rect 26332 27532 26384 27538
rect 26332 27474 26384 27480
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 26160 24806 26280 24834
rect 26252 20262 26280 24806
rect 26436 22094 26464 30262
rect 26516 29776 26568 29782
rect 26516 29718 26568 29724
rect 26528 29646 26556 29718
rect 26516 29640 26568 29646
rect 26516 29582 26568 29588
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26528 26314 26556 29242
rect 26620 28529 26648 30602
rect 26712 30598 26740 33934
rect 26804 31521 26832 34002
rect 26896 33454 26924 34167
rect 26884 33448 26936 33454
rect 26884 33390 26936 33396
rect 26884 33312 26936 33318
rect 26884 33254 26936 33260
rect 26896 33114 26924 33254
rect 26884 33108 26936 33114
rect 26884 33050 26936 33056
rect 26882 33008 26938 33017
rect 26882 32943 26938 32952
rect 26896 31890 26924 32943
rect 26988 32774 27016 35498
rect 27080 33930 27108 42298
rect 27172 41546 27200 50782
rect 27160 41540 27212 41546
rect 27160 41482 27212 41488
rect 27158 41440 27214 41449
rect 27158 41375 27214 41384
rect 27172 38214 27200 41375
rect 27160 38208 27212 38214
rect 27160 38150 27212 38156
rect 27160 36372 27212 36378
rect 27160 36314 27212 36320
rect 27172 35834 27200 36314
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 27068 33924 27120 33930
rect 27068 33866 27120 33872
rect 27068 33380 27120 33386
rect 27068 33322 27120 33328
rect 26976 32768 27028 32774
rect 26976 32710 27028 32716
rect 26974 32600 27030 32609
rect 26974 32535 26976 32544
rect 27028 32535 27030 32544
rect 26976 32506 27028 32512
rect 26974 32464 27030 32473
rect 26974 32399 26976 32408
rect 27028 32399 27030 32408
rect 26976 32370 27028 32376
rect 26974 32328 27030 32337
rect 26974 32263 27030 32272
rect 26988 32065 27016 32263
rect 26974 32056 27030 32065
rect 26974 31991 27030 32000
rect 26884 31884 26936 31890
rect 26884 31826 26936 31832
rect 26976 31748 27028 31754
rect 26976 31690 27028 31696
rect 26790 31512 26846 31521
rect 26790 31447 26846 31456
rect 26884 31408 26936 31414
rect 26882 31376 26884 31385
rect 26936 31376 26938 31385
rect 26792 31340 26844 31346
rect 26882 31311 26938 31320
rect 26792 31282 26844 31288
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26606 28520 26662 28529
rect 26606 28455 26662 28464
rect 26608 28416 26660 28422
rect 26608 28358 26660 28364
rect 26516 26308 26568 26314
rect 26516 26250 26568 26256
rect 26344 22066 26464 22094
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 25964 17808 26016 17814
rect 25964 17750 26016 17756
rect 25872 14476 25924 14482
rect 25872 14418 25924 14424
rect 25976 14006 26004 17750
rect 25964 14000 26016 14006
rect 25964 13942 26016 13948
rect 26344 13530 26372 22066
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25780 4072 25832 4078
rect 25780 4014 25832 4020
rect 25688 2576 25740 2582
rect 25688 2518 25740 2524
rect 25792 800 25820 4014
rect 25884 3398 25912 9114
rect 25976 4758 26004 11018
rect 26528 7002 26556 26250
rect 26620 7546 26648 28358
rect 26712 9722 26740 30534
rect 26804 26042 26832 31282
rect 26884 31272 26936 31278
rect 26884 31214 26936 31220
rect 26896 30598 26924 31214
rect 26988 30666 27016 31690
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 26884 30592 26936 30598
rect 26884 30534 26936 30540
rect 26896 29714 26924 30534
rect 26884 29708 26936 29714
rect 26884 29650 26936 29656
rect 26896 28014 26924 29650
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 26988 29306 27016 29582
rect 26976 29300 27028 29306
rect 26976 29242 27028 29248
rect 26976 29164 27028 29170
rect 26976 29106 27028 29112
rect 26884 28008 26936 28014
rect 26884 27950 26936 27956
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 26896 27470 26924 27814
rect 26884 27464 26936 27470
rect 26884 27406 26936 27412
rect 26884 27328 26936 27334
rect 26884 27270 26936 27276
rect 26896 26926 26924 27270
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26792 26036 26844 26042
rect 26792 25978 26844 25984
rect 26896 25362 26924 26862
rect 26988 25770 27016 29106
rect 27080 29034 27108 33322
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 27066 28248 27122 28257
rect 27066 28183 27122 28192
rect 27080 27928 27108 28183
rect 27172 28150 27200 28698
rect 27160 28144 27212 28150
rect 27160 28086 27212 28092
rect 27264 28014 27292 81670
rect 27356 81190 27384 87314
rect 27448 81433 27476 88402
rect 27620 88256 27672 88262
rect 27620 88198 27672 88204
rect 27528 87848 27580 87854
rect 27526 87816 27528 87825
rect 27580 87816 27582 87825
rect 27632 87786 27660 88198
rect 27526 87751 27582 87760
rect 27620 87780 27672 87786
rect 27620 87722 27672 87728
rect 27620 86964 27672 86970
rect 27620 86906 27672 86912
rect 27528 86828 27580 86834
rect 27528 86770 27580 86776
rect 27540 84726 27568 86770
rect 27632 86737 27660 86906
rect 27618 86728 27674 86737
rect 27618 86663 27674 86672
rect 27618 86320 27674 86329
rect 27618 86255 27674 86264
rect 27528 84720 27580 84726
rect 27526 84688 27528 84697
rect 27580 84688 27582 84697
rect 27526 84623 27582 84632
rect 27528 82476 27580 82482
rect 27528 82418 27580 82424
rect 27434 81424 27490 81433
rect 27434 81359 27490 81368
rect 27540 81274 27568 82418
rect 27448 81246 27568 81274
rect 27344 81184 27396 81190
rect 27344 81126 27396 81132
rect 27342 80880 27398 80889
rect 27342 80815 27398 80824
rect 27356 47802 27384 80815
rect 27448 79801 27476 81246
rect 27528 81184 27580 81190
rect 27528 81126 27580 81132
rect 27434 79792 27490 79801
rect 27434 79727 27490 79736
rect 27434 79656 27490 79665
rect 27434 79591 27490 79600
rect 27448 79150 27476 79591
rect 27436 79144 27488 79150
rect 27436 79086 27488 79092
rect 27436 78464 27488 78470
rect 27436 78406 27488 78412
rect 27448 74254 27476 78406
rect 27436 74248 27488 74254
rect 27436 74190 27488 74196
rect 27436 60036 27488 60042
rect 27436 59978 27488 59984
rect 27448 58041 27476 59978
rect 27434 58032 27490 58041
rect 27434 57967 27490 57976
rect 27436 57860 27488 57866
rect 27436 57802 27488 57808
rect 27448 57594 27476 57802
rect 27436 57588 27488 57594
rect 27436 57530 27488 57536
rect 27434 57216 27490 57225
rect 27434 57151 27490 57160
rect 27344 47796 27396 47802
rect 27344 47738 27396 47744
rect 27344 47660 27396 47666
rect 27344 47602 27396 47608
rect 27356 45898 27384 47602
rect 27344 45892 27396 45898
rect 27344 45834 27396 45840
rect 27448 45354 27476 57151
rect 27540 57050 27568 81126
rect 27528 57044 27580 57050
rect 27528 56986 27580 56992
rect 27528 56908 27580 56914
rect 27528 56850 27580 56856
rect 27540 56817 27568 56850
rect 27526 56808 27582 56817
rect 27526 56743 27582 56752
rect 27632 56506 27660 86255
rect 27620 56500 27672 56506
rect 27620 56442 27672 56448
rect 27528 56432 27580 56438
rect 27528 56374 27580 56380
rect 27540 52086 27568 56374
rect 27620 56228 27672 56234
rect 27620 56170 27672 56176
rect 27528 52080 27580 52086
rect 27528 52022 27580 52028
rect 27528 51604 27580 51610
rect 27528 51546 27580 51552
rect 27540 50726 27568 51546
rect 27528 50720 27580 50726
rect 27528 50662 27580 50668
rect 27540 49774 27568 50662
rect 27528 49768 27580 49774
rect 27528 49710 27580 49716
rect 27436 45348 27488 45354
rect 27436 45290 27488 45296
rect 27436 45076 27488 45082
rect 27436 45018 27488 45024
rect 27344 43376 27396 43382
rect 27344 43318 27396 43324
rect 27356 42906 27384 43318
rect 27344 42900 27396 42906
rect 27344 42842 27396 42848
rect 27344 42696 27396 42702
rect 27342 42664 27344 42673
rect 27396 42664 27398 42673
rect 27342 42599 27398 42608
rect 27344 42288 27396 42294
rect 27344 42230 27396 42236
rect 27356 41818 27384 42230
rect 27344 41812 27396 41818
rect 27344 41754 27396 41760
rect 27448 41274 27476 45018
rect 27540 45014 27568 49710
rect 27528 45008 27580 45014
rect 27528 44950 27580 44956
rect 27528 44736 27580 44742
rect 27528 44678 27580 44684
rect 27540 43178 27568 44678
rect 27528 43172 27580 43178
rect 27528 43114 27580 43120
rect 27540 42838 27568 43114
rect 27528 42832 27580 42838
rect 27528 42774 27580 42780
rect 27540 42226 27568 42774
rect 27528 42220 27580 42226
rect 27528 42162 27580 42168
rect 27528 42084 27580 42090
rect 27528 42026 27580 42032
rect 27540 41478 27568 42026
rect 27528 41472 27580 41478
rect 27528 41414 27580 41420
rect 27436 41268 27488 41274
rect 27436 41210 27488 41216
rect 27436 40520 27488 40526
rect 27436 40462 27488 40468
rect 27448 39982 27476 40462
rect 27436 39976 27488 39982
rect 27436 39918 27488 39924
rect 27540 38654 27568 41414
rect 27448 38626 27568 38654
rect 27344 38480 27396 38486
rect 27342 38448 27344 38457
rect 27396 38448 27398 38457
rect 27342 38383 27398 38392
rect 27344 37120 27396 37126
rect 27344 37062 27396 37068
rect 27356 36310 27384 37062
rect 27344 36304 27396 36310
rect 27344 36246 27396 36252
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27356 32609 27384 36110
rect 27448 34184 27476 38626
rect 27528 36032 27580 36038
rect 27528 35974 27580 35980
rect 27540 35154 27568 35974
rect 27528 35148 27580 35154
rect 27528 35090 27580 35096
rect 27448 34156 27568 34184
rect 27434 34096 27490 34105
rect 27434 34031 27490 34040
rect 27342 32600 27398 32609
rect 27342 32535 27398 32544
rect 27448 32434 27476 34031
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27344 32224 27396 32230
rect 27344 32166 27396 32172
rect 27356 31754 27384 32166
rect 27448 31958 27476 32370
rect 27540 32026 27568 34156
rect 27632 33425 27660 56170
rect 27724 51066 27752 89490
rect 27896 88936 27948 88942
rect 27896 88878 27948 88884
rect 27804 88868 27856 88874
rect 27804 88810 27856 88816
rect 27816 86426 27844 88810
rect 27804 86420 27856 86426
rect 27804 86362 27856 86368
rect 27804 85536 27856 85542
rect 27804 85478 27856 85484
rect 27816 85338 27844 85478
rect 27804 85332 27856 85338
rect 27804 85274 27856 85280
rect 27804 84108 27856 84114
rect 27804 84050 27856 84056
rect 27712 51060 27764 51066
rect 27712 51002 27764 51008
rect 27712 50720 27764 50726
rect 27712 50662 27764 50668
rect 27724 49366 27752 50662
rect 27712 49360 27764 49366
rect 27712 49302 27764 49308
rect 27712 48816 27764 48822
rect 27712 48758 27764 48764
rect 27724 41750 27752 48758
rect 27712 41744 27764 41750
rect 27712 41686 27764 41692
rect 27710 41576 27766 41585
rect 27710 41511 27766 41520
rect 27724 37194 27752 41511
rect 27816 40118 27844 84050
rect 27908 49978 27936 88878
rect 28000 51270 28028 89686
rect 28172 88596 28224 88602
rect 28172 88538 28224 88544
rect 28184 88466 28212 88538
rect 28172 88460 28224 88466
rect 28172 88402 28224 88408
rect 28172 87984 28224 87990
rect 28170 87952 28172 87961
rect 28224 87952 28226 87961
rect 28170 87887 28226 87896
rect 28080 87848 28132 87854
rect 28080 87790 28132 87796
rect 28170 87816 28226 87825
rect 27988 51264 28040 51270
rect 27988 51206 28040 51212
rect 27988 50788 28040 50794
rect 27988 50730 28040 50736
rect 28000 50318 28028 50730
rect 27988 50312 28040 50318
rect 27988 50254 28040 50260
rect 27896 49972 27948 49978
rect 27896 49914 27948 49920
rect 27896 48000 27948 48006
rect 27896 47942 27948 47948
rect 27908 47666 27936 47942
rect 27896 47660 27948 47666
rect 27896 47602 27948 47608
rect 27896 47456 27948 47462
rect 27896 47398 27948 47404
rect 27908 42634 27936 47398
rect 28092 46986 28120 87790
rect 28170 87751 28226 87760
rect 28184 87718 28212 87751
rect 28172 87712 28224 87718
rect 28172 87654 28224 87660
rect 28172 87440 28224 87446
rect 28172 87382 28224 87388
rect 28184 86902 28212 87382
rect 28276 87174 28304 94726
rect 28460 91118 28488 95882
rect 28920 93854 28948 96358
rect 28552 93826 28948 93854
rect 28356 91112 28408 91118
rect 28356 91054 28408 91060
rect 28448 91112 28500 91118
rect 28448 91054 28500 91060
rect 28264 87168 28316 87174
rect 28264 87110 28316 87116
rect 28172 86896 28224 86902
rect 28172 86838 28224 86844
rect 28184 85610 28212 86838
rect 28264 86828 28316 86834
rect 28264 86770 28316 86776
rect 28276 86329 28304 86770
rect 28262 86320 28318 86329
rect 28262 86255 28318 86264
rect 28264 86148 28316 86154
rect 28264 86090 28316 86096
rect 28172 85604 28224 85610
rect 28172 85546 28224 85552
rect 28184 85202 28212 85546
rect 28172 85196 28224 85202
rect 28172 85138 28224 85144
rect 28172 84992 28224 84998
rect 28172 84934 28224 84940
rect 28184 83722 28212 84934
rect 28276 84017 28304 86090
rect 28368 85338 28396 91054
rect 28448 89888 28500 89894
rect 28448 89830 28500 89836
rect 28460 89554 28488 89830
rect 28448 89548 28500 89554
rect 28448 89490 28500 89496
rect 28460 88874 28488 89490
rect 28448 88868 28500 88874
rect 28448 88810 28500 88816
rect 28448 88460 28500 88466
rect 28448 88402 28500 88408
rect 28460 88262 28488 88402
rect 28448 88256 28500 88262
rect 28448 88198 28500 88204
rect 28460 87786 28488 88198
rect 28448 87780 28500 87786
rect 28448 87722 28500 87728
rect 28552 87394 28580 93826
rect 29184 92200 29236 92206
rect 29184 92142 29236 92148
rect 28632 91112 28684 91118
rect 28632 91054 28684 91060
rect 28644 90710 28672 91054
rect 28724 91044 28776 91050
rect 28724 90986 28776 90992
rect 28632 90704 28684 90710
rect 28632 90646 28684 90652
rect 28644 90030 28672 90646
rect 28736 90642 28764 90986
rect 28724 90636 28776 90642
rect 28724 90578 28776 90584
rect 28632 90024 28684 90030
rect 28632 89966 28684 89972
rect 28736 89962 28764 90578
rect 29092 90568 29144 90574
rect 29092 90510 29144 90516
rect 29000 90432 29052 90438
rect 29000 90374 29052 90380
rect 29012 90030 29040 90374
rect 29000 90024 29052 90030
rect 29000 89966 29052 89972
rect 28724 89956 28776 89962
rect 28724 89898 28776 89904
rect 28736 89714 28764 89898
rect 28644 89686 28764 89714
rect 29104 89690 29132 90510
rect 28644 89554 28672 89686
rect 29092 89684 29144 89690
rect 29092 89626 29144 89632
rect 28632 89548 28684 89554
rect 28632 89490 28684 89496
rect 28816 89548 28868 89554
rect 28816 89490 28868 89496
rect 28908 89548 28960 89554
rect 28908 89490 28960 89496
rect 28644 88874 28672 89490
rect 28828 89078 28856 89490
rect 28920 89146 28948 89490
rect 28908 89140 28960 89146
rect 28908 89082 28960 89088
rect 29000 89140 29052 89146
rect 29000 89082 29052 89088
rect 28816 89072 28868 89078
rect 29012 89026 29040 89082
rect 28816 89014 28868 89020
rect 28920 88998 29040 89026
rect 28632 88868 28684 88874
rect 28632 88810 28684 88816
rect 28460 87366 28580 87394
rect 28356 85332 28408 85338
rect 28356 85274 28408 85280
rect 28460 85202 28488 87366
rect 28540 87168 28592 87174
rect 28540 87110 28592 87116
rect 28552 86766 28580 87110
rect 28540 86760 28592 86766
rect 28540 86702 28592 86708
rect 28540 86624 28592 86630
rect 28540 86566 28592 86572
rect 28552 85882 28580 86566
rect 28540 85876 28592 85882
rect 28540 85818 28592 85824
rect 28540 85672 28592 85678
rect 28540 85614 28592 85620
rect 28448 85196 28500 85202
rect 28448 85138 28500 85144
rect 28356 85060 28408 85066
rect 28356 85002 28408 85008
rect 28262 84008 28318 84017
rect 28262 83943 28318 83952
rect 28184 83694 28304 83722
rect 28172 83564 28224 83570
rect 28172 83506 28224 83512
rect 28184 83162 28212 83506
rect 28276 83473 28304 83694
rect 28262 83464 28318 83473
rect 28262 83399 28318 83408
rect 28172 83156 28224 83162
rect 28172 83098 28224 83104
rect 28264 82884 28316 82890
rect 28264 82826 28316 82832
rect 28172 82408 28224 82414
rect 28172 82350 28224 82356
rect 28184 82249 28212 82350
rect 28170 82240 28226 82249
rect 28170 82175 28226 82184
rect 28172 81388 28224 81394
rect 28172 81330 28224 81336
rect 28184 80442 28212 81330
rect 28172 80436 28224 80442
rect 28172 80378 28224 80384
rect 28276 80374 28304 82826
rect 28264 80368 28316 80374
rect 28264 80310 28316 80316
rect 28264 80232 28316 80238
rect 28264 80174 28316 80180
rect 28172 80096 28224 80102
rect 28170 80064 28172 80073
rect 28224 80064 28226 80073
rect 28170 79999 28226 80008
rect 28184 79830 28212 79999
rect 28172 79824 28224 79830
rect 28172 79766 28224 79772
rect 28184 79665 28212 79766
rect 28170 79656 28226 79665
rect 28170 79591 28226 79600
rect 28172 79552 28224 79558
rect 28172 79494 28224 79500
rect 28184 79257 28212 79494
rect 28170 79248 28226 79257
rect 28170 79183 28226 79192
rect 28170 79112 28226 79121
rect 28170 79047 28226 79056
rect 28184 79014 28212 79047
rect 28172 79008 28224 79014
rect 28172 78950 28224 78956
rect 28172 78804 28224 78810
rect 28172 78746 28224 78752
rect 28184 78674 28212 78746
rect 28172 78668 28224 78674
rect 28172 78610 28224 78616
rect 28172 74248 28224 74254
rect 28172 74190 28224 74196
rect 28080 46980 28132 46986
rect 28080 46922 28132 46928
rect 27988 46912 28040 46918
rect 27988 46854 28040 46860
rect 28000 46510 28028 46854
rect 27988 46504 28040 46510
rect 27988 46446 28040 46452
rect 27988 44192 28040 44198
rect 27988 44134 28040 44140
rect 28000 43110 28028 44134
rect 28080 43240 28132 43246
rect 28080 43182 28132 43188
rect 27988 43104 28040 43110
rect 27988 43046 28040 43052
rect 27896 42628 27948 42634
rect 27896 42570 27948 42576
rect 28000 42158 28028 43046
rect 27988 42152 28040 42158
rect 27988 42094 28040 42100
rect 27988 41744 28040 41750
rect 27988 41686 28040 41692
rect 27896 41540 27948 41546
rect 27896 41482 27948 41488
rect 27908 41313 27936 41482
rect 27894 41304 27950 41313
rect 27894 41239 27950 41248
rect 27896 40928 27948 40934
rect 27896 40870 27948 40876
rect 27804 40112 27856 40118
rect 27804 40054 27856 40060
rect 27804 39976 27856 39982
rect 27804 39918 27856 39924
rect 27816 39438 27844 39918
rect 27804 39432 27856 39438
rect 27804 39374 27856 39380
rect 27712 37188 27764 37194
rect 27712 37130 27764 37136
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 27724 34542 27752 36518
rect 27816 36038 27844 39374
rect 27908 38418 27936 40870
rect 27896 38412 27948 38418
rect 27896 38354 27948 38360
rect 27896 38208 27948 38214
rect 27896 38150 27948 38156
rect 27804 36032 27856 36038
rect 27804 35974 27856 35980
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27712 34536 27764 34542
rect 27712 34478 27764 34484
rect 27712 34400 27764 34406
rect 27712 34342 27764 34348
rect 27724 34066 27752 34342
rect 27712 34060 27764 34066
rect 27712 34002 27764 34008
rect 27712 33856 27764 33862
rect 27712 33798 27764 33804
rect 27618 33416 27674 33425
rect 27618 33351 27674 33360
rect 27620 33312 27672 33318
rect 27620 33254 27672 33260
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27436 31952 27488 31958
rect 27436 31894 27488 31900
rect 27344 31748 27396 31754
rect 27344 31690 27396 31696
rect 27448 31634 27476 31894
rect 27356 31606 27476 31634
rect 27356 31346 27384 31606
rect 27434 31512 27490 31521
rect 27434 31447 27490 31456
rect 27344 31340 27396 31346
rect 27344 31282 27396 31288
rect 27344 31204 27396 31210
rect 27344 31146 27396 31152
rect 27356 30394 27384 31146
rect 27344 30388 27396 30394
rect 27344 30330 27396 30336
rect 27344 29028 27396 29034
rect 27344 28970 27396 28976
rect 27252 28008 27304 28014
rect 27252 27950 27304 27956
rect 27080 27900 27200 27928
rect 27066 27840 27122 27849
rect 27066 27775 27122 27784
rect 27080 27674 27108 27775
rect 27068 27668 27120 27674
rect 27068 27610 27120 27616
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 26976 25764 27028 25770
rect 26976 25706 27028 25712
rect 26884 25356 26936 25362
rect 26884 25298 26936 25304
rect 26896 24750 26924 25298
rect 26884 24744 26936 24750
rect 26884 24686 26936 24692
rect 27080 23186 27108 27406
rect 27172 23866 27200 27900
rect 27356 26194 27384 28970
rect 27448 27826 27476 31447
rect 27540 31278 27568 31962
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27540 29238 27568 29650
rect 27632 29345 27660 33254
rect 27724 32881 27752 33798
rect 27710 32872 27766 32881
rect 27710 32807 27712 32816
rect 27764 32807 27766 32816
rect 27712 32778 27764 32784
rect 27724 32570 27752 32778
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27816 32450 27844 35770
rect 27908 33046 27936 38150
rect 28000 36786 28028 41686
rect 28092 39030 28120 43182
rect 28080 39024 28132 39030
rect 28080 38966 28132 38972
rect 28080 37460 28132 37466
rect 28080 37402 28132 37408
rect 27988 36780 28040 36786
rect 27988 36722 28040 36728
rect 27988 36644 28040 36650
rect 27988 36586 28040 36592
rect 28000 34678 28028 36586
rect 27988 34672 28040 34678
rect 27988 34614 28040 34620
rect 28000 33946 28028 34614
rect 28092 34066 28120 37402
rect 28080 34060 28132 34066
rect 28080 34002 28132 34008
rect 28000 33918 28120 33946
rect 27988 33584 28040 33590
rect 27988 33526 28040 33532
rect 28000 33289 28028 33526
rect 27986 33280 28042 33289
rect 27986 33215 28042 33224
rect 27986 33144 28042 33153
rect 27986 33079 28042 33088
rect 27896 33040 27948 33046
rect 27896 32982 27948 32988
rect 28000 32892 28028 33079
rect 27908 32864 28028 32892
rect 27908 32502 27936 32864
rect 27988 32768 28040 32774
rect 27986 32736 27988 32745
rect 28040 32736 28042 32745
rect 27986 32671 28042 32680
rect 27724 32422 27844 32450
rect 27896 32496 27948 32502
rect 27896 32438 27948 32444
rect 27724 31482 27752 32422
rect 27988 32360 28040 32366
rect 27986 32328 27988 32337
rect 28040 32328 28042 32337
rect 27896 32292 27948 32298
rect 27986 32263 28042 32272
rect 27896 32234 27948 32240
rect 27908 32026 27936 32234
rect 27988 32224 28040 32230
rect 27988 32166 28040 32172
rect 27896 32020 27948 32026
rect 27896 31962 27948 31968
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 27712 31476 27764 31482
rect 27712 31418 27764 31424
rect 27618 29336 27674 29345
rect 27618 29271 27674 29280
rect 27528 29232 27580 29238
rect 27816 29209 27844 31826
rect 27908 31657 27936 31826
rect 27894 31648 27950 31657
rect 27894 31583 27950 31592
rect 27896 31408 27948 31414
rect 27894 31376 27896 31385
rect 27948 31376 27950 31385
rect 27894 31311 27950 31320
rect 27896 31272 27948 31278
rect 27896 31214 27948 31220
rect 27908 30938 27936 31214
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 27896 30660 27948 30666
rect 27896 30602 27948 30608
rect 27528 29174 27580 29180
rect 27802 29200 27858 29209
rect 27802 29135 27858 29144
rect 27528 29096 27580 29102
rect 27580 29056 27752 29084
rect 27528 29038 27580 29044
rect 27724 28966 27752 29056
rect 27712 28960 27764 28966
rect 27712 28902 27764 28908
rect 27802 28928 27858 28937
rect 27802 28863 27858 28872
rect 27618 28656 27674 28665
rect 27618 28591 27674 28600
rect 27528 28484 27580 28490
rect 27528 28426 27580 28432
rect 27540 28014 27568 28426
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 27448 27798 27568 27826
rect 27434 27024 27490 27033
rect 27434 26959 27490 26968
rect 27264 26166 27384 26194
rect 27264 24274 27292 26166
rect 27344 26036 27396 26042
rect 27344 25978 27396 25984
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 27068 23180 27120 23186
rect 27068 23122 27120 23128
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26896 12434 26924 19246
rect 26804 12406 26924 12434
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 25964 4752 26016 4758
rect 25964 4694 26016 4700
rect 26608 4684 26660 4690
rect 26608 4626 26660 4632
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 26160 3602 26188 3674
rect 26056 3596 26108 3602
rect 26056 3538 26108 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 26068 800 26096 3538
rect 26148 3188 26200 3194
rect 26148 3130 26200 3136
rect 26160 3097 26188 3130
rect 26146 3088 26202 3097
rect 26146 3023 26202 3032
rect 26252 2990 26280 4422
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 26528 3058 26556 3878
rect 26516 3052 26568 3058
rect 26516 2994 26568 3000
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26332 2916 26384 2922
rect 26332 2858 26384 2864
rect 26344 800 26372 2858
rect 26620 800 26648 4626
rect 26804 3738 26832 12406
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26896 9110 26924 9318
rect 26884 9104 26936 9110
rect 26884 9046 26936 9052
rect 27356 6390 27384 25978
rect 27448 24138 27476 26959
rect 27540 25974 27568 27798
rect 27528 25968 27580 25974
rect 27528 25910 27580 25916
rect 27528 25832 27580 25838
rect 27528 25774 27580 25780
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27540 23594 27568 25774
rect 27528 23588 27580 23594
rect 27528 23530 27580 23536
rect 27632 22094 27660 28591
rect 27712 27940 27764 27946
rect 27712 27882 27764 27888
rect 27724 27849 27752 27882
rect 27710 27840 27766 27849
rect 27710 27775 27766 27784
rect 27712 27668 27764 27674
rect 27712 27610 27764 27616
rect 27724 25294 27752 27610
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27632 22066 27752 22094
rect 27724 18086 27752 22066
rect 27816 19990 27844 28863
rect 27908 25838 27936 30602
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 27804 19984 27856 19990
rect 27804 19926 27856 19932
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27908 5522 27936 23258
rect 28000 18766 28028 32166
rect 27988 18760 28040 18766
rect 27988 18702 28040 18708
rect 28092 18154 28120 33918
rect 28184 32570 28212 74190
rect 28276 37806 28304 80174
rect 28368 79257 28396 85002
rect 28448 84652 28500 84658
rect 28448 84594 28500 84600
rect 28460 84289 28488 84594
rect 28446 84280 28502 84289
rect 28446 84215 28502 84224
rect 28448 84108 28500 84114
rect 28448 84050 28500 84056
rect 28460 79937 28488 84050
rect 28446 79928 28502 79937
rect 28446 79863 28502 79872
rect 28354 79248 28410 79257
rect 28354 79183 28410 79192
rect 28356 79144 28408 79150
rect 28460 79132 28488 79863
rect 28408 79104 28488 79132
rect 28356 79086 28408 79092
rect 28356 79008 28408 79014
rect 28356 78950 28408 78956
rect 28264 37800 28316 37806
rect 28264 37742 28316 37748
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 28276 34241 28304 37062
rect 28262 34232 28318 34241
rect 28262 34167 28318 34176
rect 28368 34082 28396 78950
rect 28460 78674 28488 79104
rect 28448 78668 28500 78674
rect 28448 78610 28500 78616
rect 28460 78266 28488 78610
rect 28448 78260 28500 78266
rect 28448 78202 28500 78208
rect 28552 60734 28580 85614
rect 28644 84726 28672 88810
rect 28816 88528 28868 88534
rect 28816 88470 28868 88476
rect 28828 88398 28856 88470
rect 28920 88466 28948 88998
rect 29000 88528 29052 88534
rect 29000 88470 29052 88476
rect 28908 88460 28960 88466
rect 28908 88402 28960 88408
rect 28816 88392 28868 88398
rect 28816 88334 28868 88340
rect 29012 88058 29040 88470
rect 29092 88460 29144 88466
rect 29092 88402 29144 88408
rect 29000 88052 29052 88058
rect 29000 87994 29052 88000
rect 28816 87984 28868 87990
rect 28814 87952 28816 87961
rect 28868 87952 28870 87961
rect 28814 87887 28870 87896
rect 29000 87916 29052 87922
rect 29000 87858 29052 87864
rect 28816 87780 28868 87786
rect 28816 87722 28868 87728
rect 28724 87236 28776 87242
rect 28724 87178 28776 87184
rect 28632 84720 28684 84726
rect 28632 84662 28684 84668
rect 28632 84584 28684 84590
rect 28632 84526 28684 84532
rect 28644 84114 28672 84526
rect 28736 84182 28764 87178
rect 28828 86358 28856 87722
rect 28908 87304 28960 87310
rect 28908 87246 28960 87252
rect 28920 86834 28948 87246
rect 28908 86828 28960 86834
rect 28908 86770 28960 86776
rect 28906 86728 28962 86737
rect 28906 86663 28908 86672
rect 28960 86663 28962 86672
rect 28908 86634 28960 86640
rect 28816 86352 28868 86358
rect 28816 86294 28868 86300
rect 28816 86216 28868 86222
rect 28816 86158 28868 86164
rect 28906 86184 28962 86193
rect 28828 85882 28856 86158
rect 28906 86119 28962 86128
rect 28816 85876 28868 85882
rect 28816 85818 28868 85824
rect 28920 85626 28948 86119
rect 28828 85610 28948 85626
rect 28816 85604 28948 85610
rect 28868 85598 28948 85604
rect 28816 85546 28868 85552
rect 28828 85513 28856 85546
rect 28908 85536 28960 85542
rect 28814 85504 28870 85513
rect 28908 85478 28960 85484
rect 28814 85439 28870 85448
rect 28920 85338 28948 85478
rect 28816 85332 28868 85338
rect 28816 85274 28868 85280
rect 28908 85332 28960 85338
rect 28908 85274 28960 85280
rect 28724 84176 28776 84182
rect 28724 84118 28776 84124
rect 28632 84108 28684 84114
rect 28632 84050 28684 84056
rect 28736 83570 28764 84118
rect 28724 83564 28776 83570
rect 28724 83506 28776 83512
rect 28630 83464 28686 83473
rect 28630 83399 28686 83408
rect 28644 83366 28672 83399
rect 28632 83360 28684 83366
rect 28632 83302 28684 83308
rect 28630 83192 28686 83201
rect 28630 83127 28686 83136
rect 28644 82074 28672 83127
rect 28736 82414 28764 83506
rect 28724 82408 28776 82414
rect 28724 82350 28776 82356
rect 28724 82272 28776 82278
rect 28722 82240 28724 82249
rect 28776 82240 28778 82249
rect 28722 82175 28778 82184
rect 28632 82068 28684 82074
rect 28632 82010 28684 82016
rect 28724 81932 28776 81938
rect 28724 81874 28776 81880
rect 28632 81864 28684 81870
rect 28632 81806 28684 81812
rect 28644 81258 28672 81806
rect 28632 81252 28684 81258
rect 28632 81194 28684 81200
rect 28632 80640 28684 80646
rect 28632 80582 28684 80588
rect 28644 80306 28672 80582
rect 28632 80300 28684 80306
rect 28632 80242 28684 80248
rect 28632 80164 28684 80170
rect 28632 80106 28684 80112
rect 28644 80073 28672 80106
rect 28630 80064 28686 80073
rect 28630 79999 28686 80008
rect 28632 79892 28684 79898
rect 28632 79834 28684 79840
rect 28644 79626 28672 79834
rect 28632 79620 28684 79626
rect 28632 79562 28684 79568
rect 28630 79520 28686 79529
rect 28630 79455 28686 79464
rect 28644 79354 28672 79455
rect 28632 79348 28684 79354
rect 28632 79290 28684 79296
rect 28736 79286 28764 81874
rect 28724 79280 28776 79286
rect 28630 79248 28686 79257
rect 28724 79222 28776 79228
rect 28630 79183 28686 79192
rect 28644 73914 28672 79183
rect 28724 79008 28776 79014
rect 28724 78950 28776 78956
rect 28736 78606 28764 78950
rect 28724 78600 28776 78606
rect 28724 78542 28776 78548
rect 28724 78464 28776 78470
rect 28724 78406 28776 78412
rect 28632 73908 28684 73914
rect 28632 73850 28684 73856
rect 28644 60858 28672 73850
rect 28632 60852 28684 60858
rect 28632 60794 28684 60800
rect 28460 60706 28580 60734
rect 28460 42362 28488 60706
rect 28540 57928 28592 57934
rect 28540 57870 28592 57876
rect 28552 56930 28580 57870
rect 28632 57452 28684 57458
rect 28632 57394 28684 57400
rect 28644 57089 28672 57394
rect 28630 57080 28686 57089
rect 28630 57015 28686 57024
rect 28552 56902 28672 56930
rect 28540 56840 28592 56846
rect 28540 56782 28592 56788
rect 28552 52562 28580 56782
rect 28644 56302 28672 56902
rect 28632 56296 28684 56302
rect 28632 56238 28684 56244
rect 28632 55956 28684 55962
rect 28632 55898 28684 55904
rect 28644 55418 28672 55898
rect 28632 55412 28684 55418
rect 28632 55354 28684 55360
rect 28540 52556 28592 52562
rect 28540 52498 28592 52504
rect 28540 51468 28592 51474
rect 28540 51410 28592 51416
rect 28552 49910 28580 51410
rect 28644 50862 28672 55354
rect 28632 50856 28684 50862
rect 28632 50798 28684 50804
rect 28540 49904 28592 49910
rect 28540 49846 28592 49852
rect 28540 48068 28592 48074
rect 28540 48010 28592 48016
rect 28552 45558 28580 48010
rect 28632 46912 28684 46918
rect 28632 46854 28684 46860
rect 28540 45552 28592 45558
rect 28540 45494 28592 45500
rect 28540 45416 28592 45422
rect 28540 45358 28592 45364
rect 28448 42356 28500 42362
rect 28448 42298 28500 42304
rect 28552 42242 28580 45358
rect 28644 43450 28672 46854
rect 28632 43444 28684 43450
rect 28632 43386 28684 43392
rect 28630 43344 28686 43353
rect 28630 43279 28686 43288
rect 28460 42214 28580 42242
rect 28460 38010 28488 42214
rect 28540 42152 28592 42158
rect 28540 42094 28592 42100
rect 28448 38004 28500 38010
rect 28448 37946 28500 37952
rect 28448 37868 28500 37874
rect 28448 37810 28500 37816
rect 28460 37777 28488 37810
rect 28446 37768 28502 37777
rect 28446 37703 28502 37712
rect 28448 37664 28500 37670
rect 28448 37606 28500 37612
rect 28460 35154 28488 37606
rect 28448 35148 28500 35154
rect 28448 35090 28500 35096
rect 28448 34196 28500 34202
rect 28448 34138 28500 34144
rect 28276 34054 28396 34082
rect 28460 34066 28488 34138
rect 28448 34060 28500 34066
rect 28276 33266 28304 34054
rect 28448 34002 28500 34008
rect 28448 33584 28500 33590
rect 28552 33572 28580 42094
rect 28644 41857 28672 43279
rect 28630 41848 28686 41857
rect 28630 41783 28686 41792
rect 28632 41744 28684 41750
rect 28632 41686 28684 41692
rect 28644 38894 28672 41686
rect 28632 38888 28684 38894
rect 28632 38830 28684 38836
rect 28630 38584 28686 38593
rect 28630 38519 28686 38528
rect 28644 37942 28672 38519
rect 28632 37936 28684 37942
rect 28632 37878 28684 37884
rect 28632 37800 28684 37806
rect 28632 37742 28684 37748
rect 28644 35290 28672 37742
rect 28736 35834 28764 78406
rect 28828 56438 28856 85274
rect 29012 85202 29040 87858
rect 28908 85196 28960 85202
rect 28908 85138 28960 85144
rect 29000 85196 29052 85202
rect 29000 85138 29052 85144
rect 28816 56432 28868 56438
rect 28816 56374 28868 56380
rect 28816 52148 28868 52154
rect 28816 52090 28868 52096
rect 28828 51542 28856 52090
rect 28816 51536 28868 51542
rect 28816 51478 28868 51484
rect 28920 51074 28948 85138
rect 28998 84552 29054 84561
rect 28998 84487 29054 84496
rect 29012 84454 29040 84487
rect 29000 84448 29052 84454
rect 29000 84390 29052 84396
rect 29104 84182 29132 88402
rect 29196 85746 29224 92142
rect 29368 88868 29420 88874
rect 29368 88810 29420 88816
rect 29276 87168 29328 87174
rect 29276 87110 29328 87116
rect 29288 86426 29316 87110
rect 29276 86420 29328 86426
rect 29276 86362 29328 86368
rect 29274 86320 29330 86329
rect 29274 86255 29277 86264
rect 29329 86255 29330 86264
rect 29277 86226 29329 86232
rect 29274 86184 29330 86193
rect 29274 86119 29276 86128
rect 29328 86119 29330 86128
rect 29276 86090 29328 86096
rect 29380 85762 29408 88810
rect 29184 85740 29236 85746
rect 29184 85682 29236 85688
rect 29288 85734 29408 85762
rect 29288 85626 29316 85734
rect 29196 85598 29316 85626
rect 29092 84176 29144 84182
rect 29092 84118 29144 84124
rect 29092 84040 29144 84046
rect 29090 84008 29092 84017
rect 29144 84008 29146 84017
rect 29090 83943 29146 83952
rect 29000 83904 29052 83910
rect 29052 83864 29132 83892
rect 29000 83846 29052 83852
rect 29000 83564 29052 83570
rect 29000 83506 29052 83512
rect 29012 82618 29040 83506
rect 29104 83434 29132 83864
rect 29092 83428 29144 83434
rect 29092 83370 29144 83376
rect 29104 82822 29132 83370
rect 29092 82816 29144 82822
rect 29092 82758 29144 82764
rect 29000 82612 29052 82618
rect 29000 82554 29052 82560
rect 29104 82346 29132 82758
rect 29092 82340 29144 82346
rect 29092 82282 29144 82288
rect 29196 81938 29224 85598
rect 29368 85536 29420 85542
rect 29274 85504 29330 85513
rect 29368 85478 29420 85484
rect 29274 85439 29330 85448
rect 29288 85338 29316 85439
rect 29276 85332 29328 85338
rect 29276 85274 29328 85280
rect 29288 84522 29316 85274
rect 29380 85066 29408 85478
rect 29368 85060 29420 85066
rect 29368 85002 29420 85008
rect 29380 84697 29408 85002
rect 29366 84688 29422 84697
rect 29366 84623 29422 84632
rect 29276 84516 29328 84522
rect 29276 84458 29328 84464
rect 29380 84289 29408 84623
rect 29366 84280 29422 84289
rect 29366 84215 29422 84224
rect 29368 84176 29420 84182
rect 29368 84118 29420 84124
rect 29276 84108 29328 84114
rect 29276 84050 29328 84056
rect 29288 83502 29316 84050
rect 29276 83496 29328 83502
rect 29276 83438 29328 83444
rect 29184 81932 29236 81938
rect 29184 81874 29236 81880
rect 29182 81560 29238 81569
rect 29182 81495 29238 81504
rect 29196 81394 29224 81495
rect 29184 81388 29236 81394
rect 29184 81330 29236 81336
rect 29000 81320 29052 81326
rect 29000 81262 29052 81268
rect 29012 80730 29040 81262
rect 29184 80844 29236 80850
rect 29184 80786 29236 80792
rect 29012 80702 29132 80730
rect 29000 80300 29052 80306
rect 29000 80242 29052 80248
rect 29012 79830 29040 80242
rect 29000 79824 29052 79830
rect 29000 79766 29052 79772
rect 29000 79688 29052 79694
rect 28998 79656 29000 79665
rect 29052 79656 29054 79665
rect 28998 79591 29054 79600
rect 29104 79121 29132 80702
rect 29196 79898 29224 80786
rect 29288 80345 29316 83438
rect 29274 80336 29330 80345
rect 29274 80271 29330 80280
rect 29276 80096 29328 80102
rect 29276 80038 29328 80044
rect 29184 79892 29236 79898
rect 29184 79834 29236 79840
rect 29288 79676 29316 80038
rect 29196 79648 29316 79676
rect 29090 79112 29146 79121
rect 29090 79047 29146 79056
rect 29196 78996 29224 79648
rect 29276 79076 29328 79082
rect 29276 79018 29328 79024
rect 28998 78976 29054 78985
rect 28998 78911 29054 78920
rect 29104 78968 29224 78996
rect 29012 78062 29040 78911
rect 29000 78056 29052 78062
rect 29000 77998 29052 78004
rect 29012 77110 29040 77998
rect 29104 77926 29132 78968
rect 29288 78606 29316 79018
rect 29276 78600 29328 78606
rect 29276 78542 29328 78548
rect 29184 78464 29236 78470
rect 29184 78406 29236 78412
rect 29092 77920 29144 77926
rect 29092 77862 29144 77868
rect 29000 77104 29052 77110
rect 29000 77046 29052 77052
rect 29196 75274 29224 78406
rect 29288 77994 29316 78542
rect 29276 77988 29328 77994
rect 29276 77930 29328 77936
rect 29288 76906 29316 77930
rect 29276 76900 29328 76906
rect 29276 76842 29328 76848
rect 29184 75268 29236 75274
rect 29184 75210 29236 75216
rect 29288 73710 29316 76842
rect 29276 73704 29328 73710
rect 29276 73646 29328 73652
rect 29184 68944 29236 68950
rect 29184 68886 29236 68892
rect 29092 63028 29144 63034
rect 29092 62970 29144 62976
rect 29000 55684 29052 55690
rect 29000 55626 29052 55632
rect 29012 51490 29040 55626
rect 29104 55214 29132 62970
rect 29092 55208 29144 55214
rect 29092 55150 29144 55156
rect 29104 51610 29132 55150
rect 29196 51610 29224 68886
rect 29092 51604 29144 51610
rect 29092 51546 29144 51552
rect 29184 51604 29236 51610
rect 29184 51546 29236 51552
rect 29012 51462 29224 51490
rect 29092 51400 29144 51406
rect 28998 51368 29054 51377
rect 29092 51342 29144 51348
rect 28998 51303 29054 51312
rect 28828 51046 28948 51074
rect 28828 45082 28856 51046
rect 28908 48884 28960 48890
rect 28908 48826 28960 48832
rect 28920 46714 28948 48826
rect 28908 46708 28960 46714
rect 28908 46650 28960 46656
rect 28908 46572 28960 46578
rect 28908 46514 28960 46520
rect 28816 45076 28868 45082
rect 28816 45018 28868 45024
rect 28816 44804 28868 44810
rect 28816 44746 28868 44752
rect 28828 42158 28856 44746
rect 28920 43353 28948 46514
rect 29012 45014 29040 51303
rect 29104 45082 29132 51342
rect 29092 45076 29144 45082
rect 29092 45018 29144 45024
rect 29000 45008 29052 45014
rect 29000 44950 29052 44956
rect 29012 44282 29040 44950
rect 29104 44418 29132 45018
rect 29196 44878 29224 51462
rect 29184 44872 29236 44878
rect 29184 44814 29236 44820
rect 29104 44390 29224 44418
rect 29012 44254 29132 44282
rect 29196 44266 29224 44390
rect 29000 44192 29052 44198
rect 29000 44134 29052 44140
rect 28906 43344 28962 43353
rect 28906 43279 28962 43288
rect 28908 43104 28960 43110
rect 28908 43046 28960 43052
rect 28816 42152 28868 42158
rect 28816 42094 28868 42100
rect 28816 42016 28868 42022
rect 28816 41958 28868 41964
rect 28828 40594 28856 41958
rect 28816 40588 28868 40594
rect 28816 40530 28868 40536
rect 28816 39908 28868 39914
rect 28816 39850 28868 39856
rect 28828 38593 28856 39850
rect 28920 39574 28948 43046
rect 29012 40662 29040 44134
rect 29104 42158 29132 44254
rect 29184 44260 29236 44266
rect 29184 44202 29236 44208
rect 29184 43852 29236 43858
rect 29184 43794 29236 43800
rect 29092 42152 29144 42158
rect 29092 42094 29144 42100
rect 29104 41750 29132 42094
rect 29092 41744 29144 41750
rect 29092 41686 29144 41692
rect 29092 41608 29144 41614
rect 29196 41585 29224 43794
rect 29288 42838 29316 73646
rect 29380 70394 29408 84118
rect 29472 81394 29500 97990
rect 29644 91316 29696 91322
rect 29644 91258 29696 91264
rect 29552 87372 29604 87378
rect 29552 87314 29604 87320
rect 29564 85542 29592 87314
rect 29656 86290 29684 91258
rect 29644 86284 29696 86290
rect 29644 86226 29696 86232
rect 29644 85876 29696 85882
rect 29644 85818 29696 85824
rect 29552 85536 29604 85542
rect 29552 85478 29604 85484
rect 29656 84674 29684 85818
rect 29564 84646 29684 84674
rect 29460 81388 29512 81394
rect 29460 81330 29512 81336
rect 29460 81252 29512 81258
rect 29460 81194 29512 81200
rect 29472 80918 29500 81194
rect 29460 80912 29512 80918
rect 29460 80854 29512 80860
rect 29460 80776 29512 80782
rect 29460 80718 29512 80724
rect 29472 80170 29500 80718
rect 29460 80164 29512 80170
rect 29460 80106 29512 80112
rect 29472 77110 29500 80106
rect 29460 77104 29512 77110
rect 29460 77046 29512 77052
rect 29564 75410 29592 84646
rect 29644 84584 29696 84590
rect 29644 84526 29696 84532
rect 29656 83745 29684 84526
rect 29642 83736 29698 83745
rect 29642 83671 29698 83680
rect 29642 83600 29698 83609
rect 29642 83535 29698 83544
rect 29656 81433 29684 83535
rect 29642 81424 29698 81433
rect 29642 81359 29698 81368
rect 29644 81184 29696 81190
rect 29644 81126 29696 81132
rect 29656 80782 29684 81126
rect 29644 80776 29696 80782
rect 29644 80718 29696 80724
rect 29644 80640 29696 80646
rect 29644 80582 29696 80588
rect 29552 75404 29604 75410
rect 29552 75346 29604 75352
rect 29552 75268 29604 75274
rect 29552 75210 29604 75216
rect 29380 70366 29500 70394
rect 29368 57316 29420 57322
rect 29368 57258 29420 57264
rect 29380 51649 29408 57258
rect 29366 51640 29422 51649
rect 29366 51575 29422 51584
rect 29368 51468 29420 51474
rect 29368 51410 29420 51416
rect 29380 50182 29408 51410
rect 29368 50176 29420 50182
rect 29368 50118 29420 50124
rect 29368 49700 29420 49706
rect 29368 49642 29420 49648
rect 29380 46578 29408 49642
rect 29472 48890 29500 70366
rect 29564 60586 29592 75210
rect 29552 60580 29604 60586
rect 29552 60522 29604 60528
rect 29552 51400 29604 51406
rect 29552 51342 29604 51348
rect 29460 48884 29512 48890
rect 29460 48826 29512 48832
rect 29564 48314 29592 51342
rect 29472 48286 29592 48314
rect 29368 46572 29420 46578
rect 29368 46514 29420 46520
rect 29472 43466 29500 48286
rect 29552 44736 29604 44742
rect 29552 44678 29604 44684
rect 29380 43438 29500 43466
rect 29276 42832 29328 42838
rect 29276 42774 29328 42780
rect 29276 42696 29328 42702
rect 29276 42638 29328 42644
rect 29092 41550 29144 41556
rect 29182 41576 29238 41585
rect 29104 41002 29132 41550
rect 29182 41511 29238 41520
rect 29184 41472 29236 41478
rect 29184 41414 29236 41420
rect 29092 40996 29144 41002
rect 29092 40938 29144 40944
rect 29000 40656 29052 40662
rect 29000 40598 29052 40604
rect 28908 39568 28960 39574
rect 28908 39510 28960 39516
rect 28908 39296 28960 39302
rect 28908 39238 28960 39244
rect 28920 38865 28948 39238
rect 29104 38894 29132 40938
rect 29092 38888 29144 38894
rect 28906 38856 28962 38865
rect 29092 38830 29144 38836
rect 28906 38791 28962 38800
rect 28814 38584 28870 38593
rect 28814 38519 28870 38528
rect 29196 38434 29224 41414
rect 29288 40594 29316 42638
rect 29276 40588 29328 40594
rect 29276 40530 29328 40536
rect 29276 40112 29328 40118
rect 29276 40054 29328 40060
rect 28816 38412 28868 38418
rect 28816 38354 28868 38360
rect 29012 38406 29224 38434
rect 29288 38418 29316 40054
rect 29276 38412 29328 38418
rect 28724 35828 28776 35834
rect 28724 35770 28776 35776
rect 28632 35284 28684 35290
rect 28632 35226 28684 35232
rect 28724 34604 28776 34610
rect 28724 34546 28776 34552
rect 28632 34400 28684 34406
rect 28632 34342 28684 34348
rect 28644 33697 28672 34342
rect 28630 33688 28686 33697
rect 28630 33623 28686 33632
rect 28500 33544 28580 33572
rect 28448 33526 28500 33532
rect 28356 33448 28408 33454
rect 28408 33408 28488 33436
rect 28356 33390 28408 33396
rect 28276 33238 28396 33266
rect 28262 33144 28318 33153
rect 28262 33079 28318 33088
rect 28172 32564 28224 32570
rect 28172 32506 28224 32512
rect 28276 32450 28304 33079
rect 28184 32422 28304 32450
rect 28184 29288 28212 32422
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28276 30190 28304 32302
rect 28368 32026 28396 33238
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 28354 31920 28410 31929
rect 28354 31855 28410 31864
rect 28368 30190 28396 31855
rect 28460 31226 28488 33408
rect 28630 33416 28686 33425
rect 28540 33380 28592 33386
rect 28630 33351 28686 33360
rect 28540 33322 28592 33328
rect 28552 33289 28580 33322
rect 28538 33280 28594 33289
rect 28538 33215 28594 33224
rect 28538 32872 28594 32881
rect 28538 32807 28594 32816
rect 28552 31482 28580 32807
rect 28644 32366 28672 33351
rect 28632 32360 28684 32366
rect 28632 32302 28684 32308
rect 28632 32224 28684 32230
rect 28630 32192 28632 32201
rect 28684 32192 28686 32201
rect 28630 32127 28686 32136
rect 28540 31476 28592 31482
rect 28540 31418 28592 31424
rect 28460 31198 28580 31226
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28356 30184 28408 30190
rect 28356 30126 28408 30132
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28184 29260 28304 29288
rect 28276 28490 28304 29260
rect 28356 29028 28408 29034
rect 28356 28970 28408 28976
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 28368 28234 28396 28970
rect 28184 28206 28396 28234
rect 28184 21146 28212 28206
rect 28264 28076 28316 28082
rect 28264 28018 28316 28024
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28276 19718 28304 28018
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28172 18896 28224 18902
rect 28172 18838 28224 18844
rect 28080 18148 28132 18154
rect 28080 18090 28132 18096
rect 27540 5494 27936 5522
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27160 4004 27212 4010
rect 27160 3946 27212 3952
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 26792 3392 26844 3398
rect 26792 3334 26844 3340
rect 26804 3126 26832 3334
rect 27172 3126 27200 3946
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 27356 3466 27384 3878
rect 27344 3460 27396 3466
rect 27344 3402 27396 3408
rect 26792 3120 26844 3126
rect 26792 3062 26844 3068
rect 27160 3120 27212 3126
rect 27160 3062 27212 3068
rect 27448 2774 27476 4014
rect 27540 2990 27568 5494
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 27908 3194 27936 3878
rect 28000 3670 28028 3878
rect 27988 3664 28040 3670
rect 27988 3606 28040 3612
rect 28080 3392 28132 3398
rect 28080 3334 28132 3340
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27448 2746 27568 2774
rect 26976 2508 27028 2514
rect 26976 2450 27028 2456
rect 26988 800 27016 2450
rect 27252 1488 27304 1494
rect 27252 1430 27304 1436
rect 27264 800 27292 1430
rect 27540 800 27568 2746
rect 27804 2508 27856 2514
rect 27804 2450 27856 2456
rect 27816 800 27844 2450
rect 28092 800 28120 3334
rect 28184 2990 28212 18838
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28276 3670 28304 17818
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28368 5846 28396 16730
rect 28460 16658 28488 29990
rect 28552 23730 28580 31198
rect 28632 30592 28684 30598
rect 28632 30534 28684 30540
rect 28644 29102 28672 30534
rect 28736 30054 28764 34546
rect 28828 34513 28856 38354
rect 28906 38312 28962 38321
rect 28906 38247 28962 38256
rect 28920 37670 28948 38247
rect 28908 37664 28960 37670
rect 28908 37606 28960 37612
rect 28908 37324 28960 37330
rect 28908 37266 28960 37272
rect 28814 34504 28870 34513
rect 28814 34439 28870 34448
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 28828 25702 28856 34342
rect 28920 34202 28948 37266
rect 29012 34678 29040 38406
rect 29276 38354 29328 38360
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 29104 37330 29132 37742
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 29104 36718 29132 37266
rect 29092 36712 29144 36718
rect 29092 36654 29144 36660
rect 29000 34672 29052 34678
rect 29000 34614 29052 34620
rect 29092 34468 29144 34474
rect 29092 34410 29144 34416
rect 28908 34196 28960 34202
rect 28908 34138 28960 34144
rect 28816 25696 28868 25702
rect 28816 25638 28868 25644
rect 28632 24880 28684 24886
rect 28632 24822 28684 24828
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28540 23248 28592 23254
rect 28540 23190 28592 23196
rect 28552 21894 28580 23190
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 28356 5840 28408 5846
rect 28356 5782 28408 5788
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28264 2848 28316 2854
rect 28264 2790 28316 2796
rect 28276 1494 28304 2790
rect 28264 1488 28316 1494
rect 28264 1430 28316 1436
rect 28368 800 28396 4014
rect 28552 4010 28580 4150
rect 28540 4004 28592 4010
rect 28540 3946 28592 3952
rect 28446 3088 28502 3097
rect 28446 3023 28502 3032
rect 28460 2854 28488 3023
rect 28448 2848 28500 2854
rect 28448 2790 28500 2796
rect 28644 2774 28672 24822
rect 28920 23322 28948 34138
rect 29104 33862 29132 34410
rect 29092 33856 29144 33862
rect 29092 33798 29144 33804
rect 29000 33516 29052 33522
rect 29000 33458 29052 33464
rect 29012 28422 29040 33458
rect 29104 33386 29132 33798
rect 29092 33380 29144 33386
rect 29092 33322 29144 33328
rect 29196 33114 29224 38286
rect 29276 37868 29328 37874
rect 29276 37810 29328 37816
rect 29288 34950 29316 37810
rect 29276 34944 29328 34950
rect 29276 34886 29328 34892
rect 29184 33108 29236 33114
rect 29184 33050 29236 33056
rect 29196 32994 29224 33050
rect 29104 32966 29224 32994
rect 29000 28416 29052 28422
rect 29000 28358 29052 28364
rect 28908 23316 28960 23322
rect 28908 23258 28960 23264
rect 29104 17882 29132 32966
rect 29288 32858 29316 34886
rect 29196 32830 29316 32858
rect 29196 18902 29224 32830
rect 29276 32768 29328 32774
rect 29276 32710 29328 32716
rect 29288 29646 29316 32710
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 29184 18896 29236 18902
rect 29184 18838 29236 18844
rect 29092 17876 29144 17882
rect 29092 17818 29144 17824
rect 28908 5364 28960 5370
rect 28908 5306 28960 5312
rect 28920 3670 28948 5306
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 28552 2746 28672 2774
rect 28552 2446 28580 2746
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28736 800 28764 2450
rect 29012 800 29040 3334
rect 29288 800 29316 4014
rect 29380 3194 29408 43438
rect 29460 43240 29512 43246
rect 29460 43182 29512 43188
rect 29472 39386 29500 43182
rect 29564 39982 29592 44678
rect 29552 39976 29604 39982
rect 29552 39918 29604 39924
rect 29552 39840 29604 39846
rect 29552 39782 29604 39788
rect 29564 39574 29592 39782
rect 29552 39568 29604 39574
rect 29552 39510 29604 39516
rect 29472 39358 29592 39386
rect 29564 39302 29592 39358
rect 29552 39296 29604 39302
rect 29552 39238 29604 39244
rect 29460 38412 29512 38418
rect 29460 38354 29512 38360
rect 29472 37806 29500 38354
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29460 37460 29512 37466
rect 29460 37402 29512 37408
rect 29472 37330 29500 37402
rect 29460 37324 29512 37330
rect 29460 37266 29512 37272
rect 29460 36916 29512 36922
rect 29460 36858 29512 36864
rect 29472 34610 29500 36858
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29458 32600 29514 32609
rect 29458 32535 29514 32544
rect 29472 24410 29500 32535
rect 29460 24404 29512 24410
rect 29460 24346 29512 24352
rect 29564 5370 29592 39238
rect 29656 20466 29684 80582
rect 29748 51270 29776 115398
rect 29840 112878 29868 115942
rect 29932 114646 29960 119200
rect 30012 116884 30064 116890
rect 30012 116826 30064 116832
rect 29920 114640 29972 114646
rect 29920 114582 29972 114588
rect 30024 114578 30052 116826
rect 30012 114572 30064 114578
rect 30012 114514 30064 114520
rect 30116 113966 30144 119200
rect 30196 116748 30248 116754
rect 30196 116690 30248 116696
rect 30208 114442 30236 116690
rect 30392 116498 30420 119200
rect 30300 116470 30420 116498
rect 30300 114578 30328 116470
rect 30576 116362 30604 119200
rect 30656 117156 30708 117162
rect 30656 117098 30708 117104
rect 30392 116334 30604 116362
rect 30288 114572 30340 114578
rect 30288 114514 30340 114520
rect 30196 114436 30248 114442
rect 30196 114378 30248 114384
rect 30288 114368 30340 114374
rect 30288 114310 30340 114316
rect 30104 113960 30156 113966
rect 30104 113902 30156 113908
rect 29828 112872 29880 112878
rect 29828 112814 29880 112820
rect 30300 111794 30328 114310
rect 30392 114034 30420 116334
rect 30668 116249 30696 117098
rect 30760 116362 30788 119200
rect 31036 116822 31064 119200
rect 31116 117972 31168 117978
rect 31116 117914 31168 117920
rect 31128 117434 31156 117914
rect 31116 117428 31168 117434
rect 31116 117370 31168 117376
rect 31024 116816 31076 116822
rect 31024 116758 31076 116764
rect 31024 116680 31076 116686
rect 31024 116622 31076 116628
rect 31220 116634 31248 119200
rect 30932 116544 30984 116550
rect 30932 116486 30984 116492
rect 30760 116334 30880 116362
rect 30748 116272 30800 116278
rect 30654 116240 30710 116249
rect 30564 116204 30616 116210
rect 30748 116214 30800 116220
rect 30654 116175 30710 116184
rect 30564 116146 30616 116152
rect 30472 114912 30524 114918
rect 30472 114854 30524 114860
rect 30484 114510 30512 114854
rect 30472 114504 30524 114510
rect 30472 114446 30524 114452
rect 30380 114028 30432 114034
rect 30380 113970 30432 113976
rect 30576 113082 30604 116146
rect 30656 116068 30708 116074
rect 30656 116010 30708 116016
rect 30668 113354 30696 116010
rect 30760 113626 30788 116214
rect 30748 113620 30800 113626
rect 30748 113562 30800 113568
rect 30852 113490 30880 116334
rect 30944 114714 30972 116486
rect 31036 115802 31064 116622
rect 31220 116606 31340 116634
rect 31208 116544 31260 116550
rect 31208 116486 31260 116492
rect 31116 116204 31168 116210
rect 31116 116146 31168 116152
rect 31024 115796 31076 115802
rect 31024 115738 31076 115744
rect 31128 115258 31156 116146
rect 31220 115802 31248 116486
rect 31208 115796 31260 115802
rect 31208 115738 31260 115744
rect 31116 115252 31168 115258
rect 31116 115194 31168 115200
rect 30932 114708 30984 114714
rect 30932 114650 30984 114656
rect 31206 114064 31262 114073
rect 31206 113999 31262 114008
rect 30840 113484 30892 113490
rect 30840 113426 30892 113432
rect 30656 113348 30708 113354
rect 30656 113290 30708 113296
rect 30564 113076 30616 113082
rect 30564 113018 30616 113024
rect 31024 112940 31076 112946
rect 31024 112882 31076 112888
rect 30208 111766 30328 111794
rect 29920 99408 29972 99414
rect 29920 99350 29972 99356
rect 29828 89412 29880 89418
rect 29828 89354 29880 89360
rect 29840 88398 29868 89354
rect 29828 88392 29880 88398
rect 29828 88334 29880 88340
rect 29828 86760 29880 86766
rect 29828 86702 29880 86708
rect 29840 86426 29868 86702
rect 29828 86420 29880 86426
rect 29828 86362 29880 86368
rect 29828 86216 29880 86222
rect 29828 86158 29880 86164
rect 29840 85746 29868 86158
rect 29828 85740 29880 85746
rect 29828 85682 29880 85688
rect 29828 85060 29880 85066
rect 29828 85002 29880 85008
rect 29840 84658 29868 85002
rect 29828 84652 29880 84658
rect 29828 84594 29880 84600
rect 29828 84516 29880 84522
rect 29828 84458 29880 84464
rect 29840 82890 29868 84458
rect 29828 82884 29880 82890
rect 29828 82826 29880 82832
rect 29828 82544 29880 82550
rect 29828 82486 29880 82492
rect 29736 51264 29788 51270
rect 29736 51206 29788 51212
rect 29736 45076 29788 45082
rect 29736 45018 29788 45024
rect 29748 41682 29776 45018
rect 29736 41676 29788 41682
rect 29736 41618 29788 41624
rect 29736 40452 29788 40458
rect 29736 40394 29788 40400
rect 29748 38282 29776 40394
rect 29736 38276 29788 38282
rect 29736 38218 29788 38224
rect 29734 38176 29790 38185
rect 29734 38111 29790 38120
rect 29748 37262 29776 38111
rect 29840 37330 29868 82486
rect 29932 62354 29960 99350
rect 30104 87304 30156 87310
rect 30104 87246 30156 87252
rect 30116 86902 30144 87246
rect 30104 86896 30156 86902
rect 30104 86838 30156 86844
rect 30012 86216 30064 86222
rect 30012 86158 30064 86164
rect 30024 85184 30052 86158
rect 30104 85196 30156 85202
rect 30024 85156 30104 85184
rect 30024 84114 30052 85156
rect 30104 85138 30156 85144
rect 30012 84108 30064 84114
rect 30012 84050 30064 84056
rect 30104 83428 30156 83434
rect 30104 83370 30156 83376
rect 30012 82340 30064 82346
rect 30012 82282 30064 82288
rect 30024 78674 30052 82282
rect 30116 80986 30144 83370
rect 30104 80980 30156 80986
rect 30104 80922 30156 80928
rect 30104 80776 30156 80782
rect 30104 80718 30156 80724
rect 30116 80481 30144 80718
rect 30102 80472 30158 80481
rect 30102 80407 30158 80416
rect 30104 79756 30156 79762
rect 30104 79698 30156 79704
rect 30116 78742 30144 79698
rect 30104 78736 30156 78742
rect 30104 78678 30156 78684
rect 30012 78668 30064 78674
rect 30012 78610 30064 78616
rect 30012 77376 30064 77382
rect 30012 77318 30064 77324
rect 29920 62348 29972 62354
rect 29920 62290 29972 62296
rect 29920 56364 29972 56370
rect 29920 56306 29972 56312
rect 29932 50318 29960 56306
rect 29920 50312 29972 50318
rect 29920 50254 29972 50260
rect 29920 46096 29972 46102
rect 29920 46038 29972 46044
rect 29932 41478 29960 46038
rect 30024 45014 30052 77318
rect 30104 60648 30156 60654
rect 30104 60590 30156 60596
rect 30012 45008 30064 45014
rect 30012 44950 30064 44956
rect 30012 43240 30064 43246
rect 30012 43182 30064 43188
rect 29920 41472 29972 41478
rect 29920 41414 29972 41420
rect 30024 41290 30052 43182
rect 29932 41262 30052 41290
rect 29932 38049 29960 41262
rect 30012 40588 30064 40594
rect 30012 40530 30064 40536
rect 29918 38040 29974 38049
rect 29918 37975 29974 37984
rect 29920 37868 29972 37874
rect 29920 37810 29972 37816
rect 29828 37324 29880 37330
rect 29828 37266 29880 37272
rect 29736 37256 29788 37262
rect 29736 37198 29788 37204
rect 29826 37224 29882 37233
rect 29826 37159 29882 37168
rect 29736 37120 29788 37126
rect 29736 37062 29788 37068
rect 29748 33318 29776 37062
rect 29840 34678 29868 37159
rect 29932 36786 29960 37810
rect 30024 37505 30052 40530
rect 30010 37496 30066 37505
rect 30010 37431 30066 37440
rect 30012 37324 30064 37330
rect 30012 37266 30064 37272
rect 29920 36780 29972 36786
rect 29920 36722 29972 36728
rect 30024 36718 30052 37266
rect 30012 36712 30064 36718
rect 30012 36654 30064 36660
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29828 34672 29880 34678
rect 29828 34614 29880 34620
rect 29828 34060 29880 34066
rect 29828 34002 29880 34008
rect 29736 33312 29788 33318
rect 29736 33254 29788 33260
rect 29840 31278 29868 34002
rect 29932 32842 29960 35022
rect 30024 34202 30052 36654
rect 30012 34196 30064 34202
rect 30012 34138 30064 34144
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 29920 32836 29972 32842
rect 29920 32778 29972 32784
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 29734 31104 29790 31113
rect 29734 31039 29790 31048
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29644 17740 29696 17746
rect 29644 17682 29696 17688
rect 29552 5364 29604 5370
rect 29552 5306 29604 5312
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29564 3602 29592 3878
rect 29552 3596 29604 3602
rect 29552 3538 29604 3544
rect 29368 3188 29420 3194
rect 29368 3130 29420 3136
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29564 800 29592 2926
rect 29656 2446 29684 17682
rect 29748 12986 29776 31039
rect 30024 24818 30052 33866
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 30116 12434 30144 60590
rect 30208 51542 30236 111766
rect 30472 101856 30524 101862
rect 30472 101798 30524 101804
rect 30288 92064 30340 92070
rect 30288 92006 30340 92012
rect 30300 87854 30328 92006
rect 30380 89344 30432 89350
rect 30380 89286 30432 89292
rect 30288 87848 30340 87854
rect 30288 87790 30340 87796
rect 30288 86692 30340 86698
rect 30288 86634 30340 86640
rect 30300 86290 30328 86634
rect 30288 86284 30340 86290
rect 30288 86226 30340 86232
rect 30392 85626 30420 89286
rect 30300 85598 30420 85626
rect 30300 82550 30328 85598
rect 30380 85536 30432 85542
rect 30380 85478 30432 85484
rect 30392 84561 30420 85478
rect 30484 84658 30512 101798
rect 31036 99754 31064 112882
rect 31116 111240 31168 111246
rect 31116 111182 31168 111188
rect 31128 101454 31156 111182
rect 31220 104894 31248 113999
rect 31312 113490 31340 116606
rect 31300 113484 31352 113490
rect 31300 113426 31352 113432
rect 31404 112878 31432 119200
rect 31484 116272 31536 116278
rect 31484 116214 31536 116220
rect 31496 114170 31524 116214
rect 31588 115666 31616 119200
rect 31760 117156 31812 117162
rect 31760 117098 31812 117104
rect 31668 116748 31720 116754
rect 31668 116690 31720 116696
rect 31576 115660 31628 115666
rect 31576 115602 31628 115608
rect 31680 115258 31708 116690
rect 31668 115252 31720 115258
rect 31668 115194 31720 115200
rect 31484 114164 31536 114170
rect 31484 114106 31536 114112
rect 31576 113892 31628 113898
rect 31576 113834 31628 113840
rect 31392 112872 31444 112878
rect 31392 112814 31444 112820
rect 31588 111466 31616 113834
rect 31404 111438 31616 111466
rect 31220 104866 31340 104894
rect 31208 103624 31260 103630
rect 31208 103566 31260 103572
rect 31116 101448 31168 101454
rect 31116 101390 31168 101396
rect 31116 100224 31168 100230
rect 31116 100166 31168 100172
rect 31024 99748 31076 99754
rect 31024 99690 31076 99696
rect 30932 95328 30984 95334
rect 30932 95270 30984 95276
rect 30564 90432 30616 90438
rect 30564 90374 30616 90380
rect 30472 84652 30524 84658
rect 30472 84594 30524 84600
rect 30378 84552 30434 84561
rect 30378 84487 30434 84496
rect 30472 84516 30524 84522
rect 30472 84458 30524 84464
rect 30380 84244 30432 84250
rect 30380 84186 30432 84192
rect 30392 83910 30420 84186
rect 30380 83904 30432 83910
rect 30380 83846 30432 83852
rect 30378 83736 30434 83745
rect 30484 83706 30512 84458
rect 30378 83671 30434 83680
rect 30472 83700 30524 83706
rect 30392 83094 30420 83671
rect 30472 83642 30524 83648
rect 30380 83088 30432 83094
rect 30380 83030 30432 83036
rect 30288 82544 30340 82550
rect 30288 82486 30340 82492
rect 30472 82340 30524 82346
rect 30472 82282 30524 82288
rect 30288 82068 30340 82074
rect 30288 82010 30340 82016
rect 30300 80238 30328 82010
rect 30380 81252 30432 81258
rect 30380 81194 30432 81200
rect 30288 80232 30340 80238
rect 30288 80174 30340 80180
rect 30286 80068 30342 80077
rect 30286 80003 30342 80012
rect 30300 79286 30328 80003
rect 30392 79665 30420 81194
rect 30378 79656 30434 79665
rect 30378 79591 30434 79600
rect 30380 79552 30432 79558
rect 30380 79494 30432 79500
rect 30288 79280 30340 79286
rect 30288 79222 30340 79228
rect 30392 79098 30420 79494
rect 30300 79070 30420 79098
rect 30300 77450 30328 79070
rect 30378 78976 30434 78985
rect 30378 78911 30434 78920
rect 30392 77518 30420 78911
rect 30380 77512 30432 77518
rect 30380 77454 30432 77460
rect 30288 77444 30340 77450
rect 30288 77386 30340 77392
rect 30288 75404 30340 75410
rect 30288 75346 30340 75352
rect 30196 51536 30248 51542
rect 30196 51478 30248 51484
rect 30300 46918 30328 75346
rect 30288 46912 30340 46918
rect 30288 46854 30340 46860
rect 30380 46640 30432 46646
rect 30380 46582 30432 46588
rect 30288 44940 30340 44946
rect 30288 44882 30340 44888
rect 30196 44804 30248 44810
rect 30196 44746 30248 44752
rect 30208 39574 30236 44746
rect 30300 44334 30328 44882
rect 30288 44328 30340 44334
rect 30288 44270 30340 44276
rect 30300 43858 30328 44270
rect 30392 43858 30420 46582
rect 30288 43852 30340 43858
rect 30288 43794 30340 43800
rect 30380 43852 30432 43858
rect 30380 43794 30432 43800
rect 30300 43246 30328 43794
rect 30380 43648 30432 43654
rect 30380 43590 30432 43596
rect 30288 43240 30340 43246
rect 30288 43182 30340 43188
rect 30288 42764 30340 42770
rect 30288 42706 30340 42712
rect 30300 41478 30328 42706
rect 30288 41472 30340 41478
rect 30288 41414 30340 41420
rect 30392 39574 30420 43590
rect 30196 39568 30248 39574
rect 30196 39510 30248 39516
rect 30380 39568 30432 39574
rect 30380 39510 30432 39516
rect 30208 37210 30236 39510
rect 30378 39400 30434 39409
rect 30378 39335 30434 39344
rect 30392 38978 30420 39335
rect 30300 38950 30420 38978
rect 30300 37874 30328 38950
rect 30380 38752 30432 38758
rect 30380 38694 30432 38700
rect 30392 37942 30420 38694
rect 30380 37936 30432 37942
rect 30380 37878 30432 37884
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30288 37732 30340 37738
rect 30288 37674 30340 37680
rect 30300 37398 30328 37674
rect 30380 37664 30432 37670
rect 30380 37606 30432 37612
rect 30392 37466 30420 37606
rect 30380 37460 30432 37466
rect 30380 37402 30432 37408
rect 30288 37392 30340 37398
rect 30288 37334 30340 37340
rect 30208 37182 30420 37210
rect 30194 37088 30250 37097
rect 30194 37023 30250 37032
rect 30208 33998 30236 37023
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30300 29714 30328 35974
rect 30288 29708 30340 29714
rect 30288 29650 30340 29656
rect 30392 16574 30420 37182
rect 30484 22030 30512 82282
rect 30576 39409 30604 90374
rect 30748 88800 30800 88806
rect 30748 88742 30800 88748
rect 30760 88466 30788 88742
rect 30748 88460 30800 88466
rect 30748 88402 30800 88408
rect 30840 88392 30892 88398
rect 30840 88334 30892 88340
rect 30656 87984 30708 87990
rect 30656 87926 30708 87932
rect 30668 84726 30696 87926
rect 30852 87378 30880 88334
rect 30944 87446 30972 95270
rect 31024 88324 31076 88330
rect 31024 88266 31076 88272
rect 30932 87440 30984 87446
rect 30932 87382 30984 87388
rect 30840 87372 30892 87378
rect 30840 87314 30892 87320
rect 31036 87310 31064 88266
rect 30748 87304 30800 87310
rect 30748 87246 30800 87252
rect 31024 87304 31076 87310
rect 31024 87246 31076 87252
rect 30760 87174 30788 87246
rect 30748 87168 30800 87174
rect 30748 87110 30800 87116
rect 30840 87168 30892 87174
rect 30840 87110 30892 87116
rect 30748 86352 30800 86358
rect 30748 86294 30800 86300
rect 30760 85814 30788 86294
rect 30748 85808 30800 85814
rect 30748 85750 30800 85756
rect 30748 85604 30800 85610
rect 30748 85546 30800 85552
rect 30656 84720 30708 84726
rect 30656 84662 30708 84668
rect 30656 84040 30708 84046
rect 30656 83982 30708 83988
rect 30668 83638 30696 83982
rect 30656 83632 30708 83638
rect 30656 83574 30708 83580
rect 30656 83020 30708 83026
rect 30656 82962 30708 82968
rect 30668 82618 30696 82962
rect 30656 82612 30708 82618
rect 30656 82554 30708 82560
rect 30656 81932 30708 81938
rect 30656 81874 30708 81880
rect 30668 80646 30696 81874
rect 30656 80640 30708 80646
rect 30656 80582 30708 80588
rect 30654 80472 30710 80481
rect 30654 80407 30710 80416
rect 30668 46186 30696 80407
rect 30760 46374 30788 85546
rect 30748 46368 30800 46374
rect 30748 46310 30800 46316
rect 30668 46158 30788 46186
rect 30656 44260 30708 44266
rect 30656 44202 30708 44208
rect 30668 40390 30696 44202
rect 30760 41002 30788 46158
rect 30748 40996 30800 41002
rect 30748 40938 30800 40944
rect 30746 40896 30802 40905
rect 30746 40831 30802 40840
rect 30656 40384 30708 40390
rect 30656 40326 30708 40332
rect 30562 39400 30618 39409
rect 30562 39335 30618 39344
rect 30564 39092 30616 39098
rect 30564 39034 30616 39040
rect 30576 31754 30604 39034
rect 30668 37913 30696 40326
rect 30654 37904 30710 37913
rect 30654 37839 30710 37848
rect 30656 37732 30708 37738
rect 30656 37674 30708 37680
rect 30668 35086 30696 37674
rect 30656 35080 30708 35086
rect 30656 35022 30708 35028
rect 30760 34354 30788 40831
rect 30852 38010 30880 87110
rect 31036 86902 31064 87246
rect 31024 86896 31076 86902
rect 31024 86838 31076 86844
rect 30932 86692 30984 86698
rect 30932 86634 30984 86640
rect 30944 40905 30972 86634
rect 31024 86080 31076 86086
rect 31024 86022 31076 86028
rect 30930 40896 30986 40905
rect 30930 40831 30986 40840
rect 30930 40760 30986 40769
rect 30930 40695 30986 40704
rect 30840 38004 30892 38010
rect 30840 37946 30892 37952
rect 30838 37904 30894 37913
rect 30838 37839 30894 37848
rect 30668 34326 30788 34354
rect 30668 32774 30696 34326
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30656 32768 30708 32774
rect 30656 32710 30708 32716
rect 30576 31726 30696 31754
rect 30472 22024 30524 22030
rect 30472 21966 30524 21972
rect 30392 16546 30512 16574
rect 29840 12406 30144 12434
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 29748 3602 29776 4422
rect 29736 3596 29788 3602
rect 29736 3538 29788 3544
rect 29840 2650 29868 12406
rect 30196 4684 30248 4690
rect 30196 4626 30248 4632
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29932 1442 29960 3130
rect 29840 1414 29960 1442
rect 29840 800 29868 1414
rect 30208 800 30236 4626
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 30300 3398 30328 4082
rect 30392 3670 30420 4082
rect 30484 4010 30512 16546
rect 30564 5772 30616 5778
rect 30564 5714 30616 5720
rect 30576 4078 30604 5714
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 30472 4004 30524 4010
rect 30472 3946 30524 3952
rect 30668 3670 30696 31726
rect 30760 26994 30788 34138
rect 30748 26988 30800 26994
rect 30748 26930 30800 26936
rect 30852 4078 30880 37839
rect 30944 32026 30972 40695
rect 30932 32020 30984 32026
rect 30932 31962 30984 31968
rect 31036 31414 31064 86022
rect 31128 83026 31156 100166
rect 31220 88398 31248 103566
rect 31312 103222 31340 104866
rect 31404 104242 31432 111438
rect 31484 111308 31536 111314
rect 31484 111250 31536 111256
rect 31392 104236 31444 104242
rect 31392 104178 31444 104184
rect 31300 103216 31352 103222
rect 31300 103158 31352 103164
rect 31496 98666 31524 111250
rect 31576 99136 31628 99142
rect 31576 99078 31628 99084
rect 31484 98660 31536 98666
rect 31484 98602 31536 98608
rect 31300 96960 31352 96966
rect 31300 96902 31352 96908
rect 31312 88874 31340 96902
rect 31392 90500 31444 90506
rect 31392 90442 31444 90448
rect 31404 89714 31432 90442
rect 31404 89686 31524 89714
rect 31496 89486 31524 89686
rect 31484 89480 31536 89486
rect 31484 89422 31536 89428
rect 31496 89078 31524 89422
rect 31484 89072 31536 89078
rect 31484 89014 31536 89020
rect 31300 88868 31352 88874
rect 31300 88810 31352 88816
rect 31392 88460 31444 88466
rect 31392 88402 31444 88408
rect 31208 88392 31260 88398
rect 31208 88334 31260 88340
rect 31300 87780 31352 87786
rect 31300 87722 31352 87728
rect 31208 87508 31260 87514
rect 31208 87450 31260 87456
rect 31220 86698 31248 87450
rect 31208 86692 31260 86698
rect 31208 86634 31260 86640
rect 31208 86080 31260 86086
rect 31208 86022 31260 86028
rect 31220 85678 31248 86022
rect 31208 85672 31260 85678
rect 31208 85614 31260 85620
rect 31208 85060 31260 85066
rect 31208 85002 31260 85008
rect 31220 84590 31248 85002
rect 31208 84584 31260 84590
rect 31208 84526 31260 84532
rect 31220 84046 31248 84526
rect 31208 84040 31260 84046
rect 31208 83982 31260 83988
rect 31206 83872 31262 83881
rect 31206 83807 31262 83816
rect 31220 83638 31248 83807
rect 31208 83632 31260 83638
rect 31208 83574 31260 83580
rect 31208 83496 31260 83502
rect 31208 83438 31260 83444
rect 31116 83020 31168 83026
rect 31116 82962 31168 82968
rect 31220 82958 31248 83438
rect 31208 82952 31260 82958
rect 31208 82894 31260 82900
rect 31220 82414 31248 82894
rect 31116 82408 31168 82414
rect 31116 82350 31168 82356
rect 31208 82408 31260 82414
rect 31208 82350 31260 82356
rect 31128 81569 31156 82350
rect 31220 81802 31248 82350
rect 31208 81796 31260 81802
rect 31208 81738 31260 81744
rect 31114 81560 31170 81569
rect 31114 81495 31170 81504
rect 31220 81326 31248 81738
rect 31116 81320 31168 81326
rect 31116 81262 31168 81268
rect 31208 81320 31260 81326
rect 31208 81262 31260 81268
rect 31128 80306 31156 81262
rect 31206 81016 31262 81025
rect 31206 80951 31208 80960
rect 31260 80951 31262 80960
rect 31208 80922 31260 80928
rect 31208 80844 31260 80850
rect 31208 80786 31260 80792
rect 31116 80300 31168 80306
rect 31116 80242 31168 80248
rect 31116 80096 31168 80102
rect 31116 80038 31168 80044
rect 31128 51074 31156 80038
rect 31220 77382 31248 80786
rect 31208 77376 31260 77382
rect 31208 77318 31260 77324
rect 31312 51074 31340 87722
rect 31404 80481 31432 88402
rect 31496 88398 31524 89014
rect 31484 88392 31536 88398
rect 31484 88334 31536 88340
rect 31496 87922 31524 88334
rect 31484 87916 31536 87922
rect 31484 87858 31536 87864
rect 31496 86154 31524 87858
rect 31484 86148 31536 86154
rect 31484 86090 31536 86096
rect 31484 85672 31536 85678
rect 31484 85614 31536 85620
rect 31496 85134 31524 85614
rect 31484 85128 31536 85134
rect 31484 85070 31536 85076
rect 31484 84720 31536 84726
rect 31484 84662 31536 84668
rect 31496 84590 31524 84662
rect 31484 84584 31536 84590
rect 31484 84526 31536 84532
rect 31496 84114 31524 84526
rect 31484 84108 31536 84114
rect 31484 84050 31536 84056
rect 31496 84017 31524 84050
rect 31482 84008 31538 84017
rect 31482 83943 31538 83952
rect 31484 83904 31536 83910
rect 31484 83846 31536 83852
rect 31390 80472 31446 80481
rect 31390 80407 31446 80416
rect 31392 80368 31444 80374
rect 31390 80336 31392 80345
rect 31444 80336 31446 80345
rect 31390 80271 31446 80280
rect 31392 79620 31444 79626
rect 31392 79562 31444 79568
rect 31404 78198 31432 79562
rect 31392 78192 31444 78198
rect 31392 78134 31444 78140
rect 31496 60734 31524 83846
rect 31588 82482 31616 99078
rect 31668 88596 31720 88602
rect 31668 88538 31720 88544
rect 31680 87854 31708 88538
rect 31668 87848 31720 87854
rect 31668 87790 31720 87796
rect 31668 86896 31720 86902
rect 31668 86838 31720 86844
rect 31680 86154 31708 86838
rect 31668 86148 31720 86154
rect 31668 86090 31720 86096
rect 31680 84250 31708 86090
rect 31668 84244 31720 84250
rect 31668 84186 31720 84192
rect 31668 83700 31720 83706
rect 31668 83642 31720 83648
rect 31576 82476 31628 82482
rect 31576 82418 31628 82424
rect 31576 82340 31628 82346
rect 31576 82282 31628 82288
rect 31588 81938 31616 82282
rect 31576 81932 31628 81938
rect 31576 81874 31628 81880
rect 31588 81530 31616 81874
rect 31576 81524 31628 81530
rect 31576 81466 31628 81472
rect 31576 81252 31628 81258
rect 31576 81194 31628 81200
rect 31588 76294 31616 81194
rect 31576 76288 31628 76294
rect 31576 76230 31628 76236
rect 31404 60706 31524 60734
rect 31404 54126 31432 60706
rect 31392 54120 31444 54126
rect 31392 54062 31444 54068
rect 31128 51046 31248 51074
rect 31312 51046 31432 51074
rect 31220 46458 31248 51046
rect 31220 46430 31340 46458
rect 31208 46368 31260 46374
rect 31208 46310 31260 46316
rect 31116 45892 31168 45898
rect 31116 45834 31168 45840
rect 31128 43722 31156 45834
rect 31116 43716 31168 43722
rect 31116 43658 31168 43664
rect 31116 41812 31168 41818
rect 31116 41754 31168 41760
rect 31128 40769 31156 41754
rect 31114 40760 31170 40769
rect 31114 40695 31170 40704
rect 31114 40080 31170 40089
rect 31114 40015 31170 40024
rect 31024 31408 31076 31414
rect 31024 31350 31076 31356
rect 31128 31346 31156 40015
rect 31116 31340 31168 31346
rect 31116 31282 31168 31288
rect 31116 29572 31168 29578
rect 31116 29514 31168 29520
rect 31024 27600 31076 27606
rect 31024 27542 31076 27548
rect 31036 4842 31064 27542
rect 31128 11898 31156 29514
rect 31220 29170 31248 46310
rect 31312 44198 31340 46430
rect 31300 44192 31352 44198
rect 31300 44134 31352 44140
rect 31300 43852 31352 43858
rect 31300 43794 31352 43800
rect 31312 39846 31340 43794
rect 31300 39840 31352 39846
rect 31300 39782 31352 39788
rect 31300 39568 31352 39574
rect 31300 39510 31352 39516
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31312 24614 31340 39510
rect 31404 36922 31432 51046
rect 31576 45348 31628 45354
rect 31576 45290 31628 45296
rect 31484 43784 31536 43790
rect 31484 43726 31536 43732
rect 31496 39370 31524 43726
rect 31588 42294 31616 45290
rect 31576 42288 31628 42294
rect 31576 42230 31628 42236
rect 31576 40996 31628 41002
rect 31576 40938 31628 40944
rect 31484 39364 31536 39370
rect 31484 39306 31536 39312
rect 31496 39098 31524 39306
rect 31484 39092 31536 39098
rect 31484 39034 31536 39040
rect 31484 38480 31536 38486
rect 31484 38422 31536 38428
rect 31496 37874 31524 38422
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 31392 36916 31444 36922
rect 31392 36858 31444 36864
rect 31588 35494 31616 40938
rect 31576 35488 31628 35494
rect 31576 35430 31628 35436
rect 31392 35284 31444 35290
rect 31392 35226 31444 35232
rect 31404 25498 31432 35226
rect 31576 32292 31628 32298
rect 31576 32234 31628 32240
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31208 24064 31260 24070
rect 31208 24006 31260 24012
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31220 9178 31248 24006
rect 31588 22094 31616 32234
rect 31680 27674 31708 83642
rect 31772 62966 31800 117098
rect 31864 115734 31892 119200
rect 31944 116272 31996 116278
rect 31944 116214 31996 116220
rect 31852 115728 31904 115734
rect 31852 115670 31904 115676
rect 31956 114170 31984 116214
rect 32048 115054 32076 119200
rect 32128 116136 32180 116142
rect 32128 116078 32180 116084
rect 32036 115048 32088 115054
rect 32036 114990 32088 114996
rect 31944 114164 31996 114170
rect 31944 114106 31996 114112
rect 32140 113354 32168 116078
rect 32232 114578 32260 119200
rect 32312 117156 32364 117162
rect 32312 117098 32364 117104
rect 32220 114572 32272 114578
rect 32220 114514 32272 114520
rect 32128 113348 32180 113354
rect 32128 113290 32180 113296
rect 31944 112804 31996 112810
rect 31944 112746 31996 112752
rect 31956 108390 31984 112746
rect 32324 109034 32352 117098
rect 32404 116136 32456 116142
rect 32404 116078 32456 116084
rect 32416 115258 32444 116078
rect 32404 115252 32456 115258
rect 32404 115194 32456 115200
rect 32404 114980 32456 114986
rect 32404 114922 32456 114928
rect 32232 109006 32352 109034
rect 31944 108384 31996 108390
rect 31944 108326 31996 108332
rect 32036 105256 32088 105262
rect 32036 105198 32088 105204
rect 31944 91044 31996 91050
rect 31944 90986 31996 90992
rect 31852 90636 31904 90642
rect 31852 90578 31904 90584
rect 31864 89554 31892 90578
rect 31852 89548 31904 89554
rect 31852 89490 31904 89496
rect 31864 89350 31892 89490
rect 31852 89344 31904 89350
rect 31852 89286 31904 89292
rect 31852 88868 31904 88874
rect 31852 88810 31904 88816
rect 31760 62960 31812 62966
rect 31760 62902 31812 62908
rect 31758 62520 31814 62529
rect 31758 62455 31814 62464
rect 31772 62422 31800 62455
rect 31760 62416 31812 62422
rect 31760 62358 31812 62364
rect 31760 53780 31812 53786
rect 31760 53722 31812 53728
rect 31772 51066 31800 53722
rect 31760 51060 31812 51066
rect 31760 51002 31812 51008
rect 31758 43208 31814 43217
rect 31758 43143 31814 43152
rect 31772 32434 31800 43143
rect 31864 37262 31892 88810
rect 31956 80866 31984 90986
rect 32048 81002 32076 105198
rect 32128 100972 32180 100978
rect 32128 100914 32180 100920
rect 32140 86834 32168 100914
rect 32232 100026 32260 109006
rect 32416 106962 32444 114922
rect 32508 113966 32536 119200
rect 32692 116192 32720 119200
rect 32772 116748 32824 116754
rect 32772 116690 32824 116696
rect 32600 116164 32720 116192
rect 32600 115190 32628 116164
rect 32680 116068 32732 116074
rect 32680 116010 32732 116016
rect 32588 115184 32640 115190
rect 32588 115126 32640 115132
rect 32496 113960 32548 113966
rect 32496 113902 32548 113908
rect 32692 113626 32720 116010
rect 32784 114646 32812 116690
rect 32876 116192 32904 119200
rect 33048 116816 33100 116822
rect 33048 116758 33100 116764
rect 32876 116164 32996 116192
rect 32864 116068 32916 116074
rect 32864 116010 32916 116016
rect 32772 114640 32824 114646
rect 32772 114582 32824 114588
rect 32772 114504 32824 114510
rect 32772 114446 32824 114452
rect 32680 113620 32732 113626
rect 32680 113562 32732 113568
rect 32784 110090 32812 114446
rect 32876 114170 32904 116010
rect 32864 114164 32916 114170
rect 32864 114106 32916 114112
rect 32968 113490 32996 116164
rect 33060 114034 33088 116758
rect 33152 116550 33180 119200
rect 33140 116544 33192 116550
rect 33140 116486 33192 116492
rect 33140 116272 33192 116278
rect 33140 116214 33192 116220
rect 33048 114028 33100 114034
rect 33048 113970 33100 113976
rect 32956 113484 33008 113490
rect 32956 113426 33008 113432
rect 33152 113082 33180 116214
rect 33232 114572 33284 114578
rect 33232 114514 33284 114520
rect 33140 113076 33192 113082
rect 33140 113018 33192 113024
rect 33140 112736 33192 112742
rect 33140 112678 33192 112684
rect 32772 110084 32824 110090
rect 32772 110026 32824 110032
rect 32680 109064 32732 109070
rect 32680 109006 32732 109012
rect 32404 106956 32456 106962
rect 32404 106898 32456 106904
rect 32312 103556 32364 103562
rect 32312 103498 32364 103504
rect 32220 100020 32272 100026
rect 32220 99962 32272 99968
rect 32324 90642 32352 103498
rect 32496 102196 32548 102202
rect 32496 102138 32548 102144
rect 32404 98116 32456 98122
rect 32404 98058 32456 98064
rect 32312 90636 32364 90642
rect 32312 90578 32364 90584
rect 32220 89956 32272 89962
rect 32220 89898 32272 89904
rect 32128 86828 32180 86834
rect 32128 86770 32180 86776
rect 32128 86284 32180 86290
rect 32128 86226 32180 86232
rect 32140 85746 32168 86226
rect 32128 85740 32180 85746
rect 32128 85682 32180 85688
rect 32140 85202 32168 85682
rect 32128 85196 32180 85202
rect 32128 85138 32180 85144
rect 32048 80974 32168 81002
rect 31956 80838 32076 80866
rect 31944 80776 31996 80782
rect 31944 80718 31996 80724
rect 31956 80442 31984 80718
rect 31944 80436 31996 80442
rect 31944 80378 31996 80384
rect 32048 80186 32076 80838
rect 31956 80158 32076 80186
rect 31956 38758 31984 80158
rect 32140 80054 32168 80974
rect 32048 80026 32168 80054
rect 31944 38752 31996 38758
rect 31944 38694 31996 38700
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 31852 36304 31904 36310
rect 31852 36246 31904 36252
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31864 29238 31892 36246
rect 31944 35692 31996 35698
rect 31944 35634 31996 35640
rect 31852 29232 31904 29238
rect 31956 29209 31984 35634
rect 31852 29174 31904 29180
rect 31942 29200 31998 29209
rect 31942 29135 31998 29144
rect 31944 28484 31996 28490
rect 31944 28426 31996 28432
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31956 23526 31984 28426
rect 32048 24886 32076 80026
rect 32128 62756 32180 62762
rect 32128 62698 32180 62704
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 31944 23520 31996 23526
rect 31944 23462 31996 23468
rect 31404 22066 31616 22094
rect 31404 19174 31432 22066
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31208 9172 31260 9178
rect 31208 9114 31260 9120
rect 31300 5160 31352 5166
rect 31300 5102 31352 5108
rect 31036 4814 31156 4842
rect 31024 4684 31076 4690
rect 31024 4626 31076 4632
rect 30840 4072 30892 4078
rect 30840 4014 30892 4020
rect 30748 3936 30800 3942
rect 30748 3878 30800 3884
rect 30380 3664 30432 3670
rect 30380 3606 30432 3612
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30656 3664 30708 3670
rect 30656 3606 30708 3612
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 30484 2922 30512 3606
rect 30564 3596 30616 3602
rect 30564 3538 30616 3544
rect 30576 3194 30604 3538
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30472 2916 30524 2922
rect 30472 2858 30524 2864
rect 30472 2508 30524 2514
rect 30472 2450 30524 2456
rect 30484 800 30512 2450
rect 30760 800 30788 3878
rect 31036 800 31064 4626
rect 31128 2922 31156 4814
rect 31116 2916 31168 2922
rect 31116 2858 31168 2864
rect 31312 800 31340 5102
rect 31760 5092 31812 5098
rect 31760 5034 31812 5040
rect 31392 4480 31444 4486
rect 31392 4422 31444 4428
rect 31404 3466 31432 4422
rect 31576 3936 31628 3942
rect 31576 3878 31628 3884
rect 31484 3664 31536 3670
rect 31484 3606 31536 3612
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 31496 3058 31524 3606
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 31588 800 31616 3878
rect 31668 3188 31720 3194
rect 31668 3130 31720 3136
rect 31680 3040 31708 3130
rect 31772 3040 31800 5034
rect 31680 3012 31800 3040
rect 32140 2650 32168 62698
rect 32232 40118 32260 89898
rect 32312 89684 32364 89690
rect 32312 89626 32364 89632
rect 32324 88602 32352 89626
rect 32312 88596 32364 88602
rect 32312 88538 32364 88544
rect 32416 88466 32444 98058
rect 32404 88460 32456 88466
rect 32404 88402 32456 88408
rect 32312 88392 32364 88398
rect 32312 88334 32364 88340
rect 32324 87854 32352 88334
rect 32404 88324 32456 88330
rect 32404 88266 32456 88272
rect 32416 87990 32444 88266
rect 32508 87990 32536 102138
rect 32588 89888 32640 89894
rect 32588 89830 32640 89836
rect 32600 88942 32628 89830
rect 32588 88936 32640 88942
rect 32588 88878 32640 88884
rect 32588 88460 32640 88466
rect 32588 88402 32640 88408
rect 32404 87984 32456 87990
rect 32404 87926 32456 87932
rect 32496 87984 32548 87990
rect 32496 87926 32548 87932
rect 32312 87848 32364 87854
rect 32312 87790 32364 87796
rect 32324 87378 32352 87790
rect 32600 87786 32628 88402
rect 32588 87780 32640 87786
rect 32588 87722 32640 87728
rect 32404 87712 32456 87718
rect 32404 87654 32456 87660
rect 32496 87712 32548 87718
rect 32496 87654 32548 87660
rect 32416 87446 32444 87654
rect 32404 87440 32456 87446
rect 32404 87382 32456 87388
rect 32508 87378 32536 87654
rect 32312 87372 32364 87378
rect 32312 87314 32364 87320
rect 32496 87372 32548 87378
rect 32496 87314 32548 87320
rect 32324 86426 32352 87314
rect 32404 87168 32456 87174
rect 32404 87110 32456 87116
rect 32416 86766 32444 87110
rect 32494 87000 32550 87009
rect 32600 86970 32628 87722
rect 32494 86935 32496 86944
rect 32548 86935 32550 86944
rect 32588 86964 32640 86970
rect 32496 86906 32548 86912
rect 32588 86906 32640 86912
rect 32404 86760 32456 86766
rect 32456 86720 32536 86748
rect 32404 86702 32456 86708
rect 32404 86624 32456 86630
rect 32404 86566 32456 86572
rect 32312 86420 32364 86426
rect 32312 86362 32364 86368
rect 32416 85746 32444 86566
rect 32508 86290 32536 86720
rect 32588 86692 32640 86698
rect 32588 86634 32640 86640
rect 32496 86284 32548 86290
rect 32496 86226 32548 86232
rect 32404 85740 32456 85746
rect 32404 85682 32456 85688
rect 32600 85610 32628 86634
rect 32692 85678 32720 109006
rect 32772 108520 32824 108526
rect 32772 108462 32824 108468
rect 32784 94586 32812 108462
rect 32956 107636 33008 107642
rect 32956 107578 33008 107584
rect 32864 106344 32916 106350
rect 32864 106286 32916 106292
rect 32772 94580 32824 94586
rect 32772 94522 32824 94528
rect 32876 91186 32904 106286
rect 32864 91180 32916 91186
rect 32864 91122 32916 91128
rect 32772 91112 32824 91118
rect 32968 91066 32996 107578
rect 33048 94580 33100 94586
rect 33048 94522 33100 94528
rect 32772 91054 32824 91060
rect 32784 90098 32812 91054
rect 32876 91038 32996 91066
rect 32876 90642 32904 91038
rect 32956 90976 33008 90982
rect 32956 90918 33008 90924
rect 32864 90636 32916 90642
rect 32864 90578 32916 90584
rect 32864 90432 32916 90438
rect 32864 90374 32916 90380
rect 32772 90092 32824 90098
rect 32772 90034 32824 90040
rect 32784 89690 32812 90034
rect 32772 89684 32824 89690
rect 32772 89626 32824 89632
rect 32772 89480 32824 89486
rect 32772 89422 32824 89428
rect 32784 89078 32812 89422
rect 32772 89072 32824 89078
rect 32772 89014 32824 89020
rect 32772 88936 32824 88942
rect 32772 88878 32824 88884
rect 32784 88602 32812 88878
rect 32772 88596 32824 88602
rect 32772 88538 32824 88544
rect 32784 86902 32812 88538
rect 32876 87174 32904 90374
rect 32968 90030 32996 90918
rect 33060 90166 33088 94522
rect 33048 90160 33100 90166
rect 33048 90102 33100 90108
rect 32956 90024 33008 90030
rect 32956 89966 33008 89972
rect 32968 89350 32996 89966
rect 32956 89344 33008 89350
rect 32956 89286 33008 89292
rect 32968 88942 32996 89286
rect 32956 88936 33008 88942
rect 32956 88878 33008 88884
rect 32968 87514 32996 88878
rect 33048 88596 33100 88602
rect 33048 88538 33100 88544
rect 32956 87508 33008 87514
rect 32956 87450 33008 87456
rect 32956 87372 33008 87378
rect 32956 87314 33008 87320
rect 32864 87168 32916 87174
rect 32864 87110 32916 87116
rect 32968 86986 32996 87314
rect 32876 86958 32996 86986
rect 32772 86896 32824 86902
rect 32772 86838 32824 86844
rect 32772 86760 32824 86766
rect 32770 86728 32772 86737
rect 32824 86728 32826 86737
rect 32770 86663 32826 86672
rect 32772 86624 32824 86630
rect 32772 86566 32824 86572
rect 32680 85672 32732 85678
rect 32680 85614 32732 85620
rect 32588 85604 32640 85610
rect 32588 85546 32640 85552
rect 32496 85536 32548 85542
rect 32496 85478 32548 85484
rect 32312 84516 32364 84522
rect 32312 84458 32364 84464
rect 32220 40112 32272 40118
rect 32220 40054 32272 40060
rect 32220 39908 32272 39914
rect 32220 39850 32272 39856
rect 32232 16182 32260 39850
rect 32324 39574 32352 84458
rect 32404 81320 32456 81326
rect 32404 81262 32456 81268
rect 32416 78849 32444 81262
rect 32402 78840 32458 78849
rect 32402 78775 32458 78784
rect 32404 63232 32456 63238
rect 32404 63174 32456 63180
rect 32416 63034 32444 63174
rect 32404 63028 32456 63034
rect 32404 62970 32456 62976
rect 32404 62688 32456 62694
rect 32404 62630 32456 62636
rect 32312 39568 32364 39574
rect 32312 39510 32364 39516
rect 32312 37460 32364 37466
rect 32312 37402 32364 37408
rect 32324 29510 32352 37402
rect 32312 29504 32364 29510
rect 32312 29446 32364 29452
rect 32312 28688 32364 28694
rect 32310 28656 32312 28665
rect 32364 28656 32366 28665
rect 32310 28591 32366 28600
rect 32220 16176 32272 16182
rect 32220 16118 32272 16124
rect 32416 3194 32444 62630
rect 32508 43178 32536 85478
rect 32600 80714 32628 85546
rect 32680 81252 32732 81258
rect 32680 81194 32732 81200
rect 32588 80708 32640 80714
rect 32588 80650 32640 80656
rect 32600 80170 32628 80650
rect 32588 80164 32640 80170
rect 32588 80106 32640 80112
rect 32600 78470 32628 80106
rect 32588 78464 32640 78470
rect 32588 78406 32640 78412
rect 32588 75948 32640 75954
rect 32588 75890 32640 75896
rect 32600 57390 32628 75890
rect 32588 57384 32640 57390
rect 32588 57326 32640 57332
rect 32692 54534 32720 81194
rect 32680 54528 32732 54534
rect 32680 54470 32732 54476
rect 32784 51074 32812 86566
rect 32876 86290 32904 86958
rect 32956 86896 33008 86902
rect 32956 86838 33008 86844
rect 32864 86284 32916 86290
rect 32864 86226 32916 86232
rect 32876 85082 32904 86226
rect 32968 85678 32996 86838
rect 32956 85672 33008 85678
rect 32956 85614 33008 85620
rect 32968 85338 32996 85614
rect 32956 85332 33008 85338
rect 32956 85274 33008 85280
rect 33060 85270 33088 88538
rect 33048 85264 33100 85270
rect 33048 85206 33100 85212
rect 32876 85054 33088 85082
rect 32956 84992 33008 84998
rect 32956 84934 33008 84940
rect 32864 81728 32916 81734
rect 32864 81670 32916 81676
rect 32876 80850 32904 81670
rect 32864 80844 32916 80850
rect 32864 80786 32916 80792
rect 32968 80238 32996 84934
rect 33060 82006 33088 85054
rect 33048 82000 33100 82006
rect 33048 81942 33100 81948
rect 33060 81326 33088 81942
rect 33048 81320 33100 81326
rect 33048 81262 33100 81268
rect 32956 80232 33008 80238
rect 32956 80174 33008 80180
rect 33060 79694 33088 81262
rect 33048 79688 33100 79694
rect 33048 79630 33100 79636
rect 32864 65476 32916 65482
rect 32864 65418 32916 65424
rect 32692 51046 32812 51074
rect 32876 51066 32904 65418
rect 33152 63594 33180 112678
rect 33244 108458 33272 114514
rect 33336 112878 33364 119200
rect 33416 116680 33468 116686
rect 33416 116622 33468 116628
rect 33428 115462 33456 116622
rect 33416 115456 33468 115462
rect 33416 115398 33468 115404
rect 33416 114980 33468 114986
rect 33416 114922 33468 114928
rect 33324 112872 33376 112878
rect 33324 112814 33376 112820
rect 33232 108452 33284 108458
rect 33232 108394 33284 108400
rect 33232 107840 33284 107846
rect 33232 107782 33284 107788
rect 33244 106350 33272 107782
rect 33232 106344 33284 106350
rect 33232 106286 33284 106292
rect 33324 105664 33376 105670
rect 33324 105606 33376 105612
rect 33336 98122 33364 105606
rect 33324 98116 33376 98122
rect 33324 98058 33376 98064
rect 33232 90636 33284 90642
rect 33232 90578 33284 90584
rect 33244 88466 33272 90578
rect 33324 90160 33376 90166
rect 33324 90102 33376 90108
rect 33336 89690 33364 90102
rect 33324 89684 33376 89690
rect 33324 89626 33376 89632
rect 33324 89344 33376 89350
rect 33324 89286 33376 89292
rect 33232 88460 33284 88466
rect 33232 88402 33284 88408
rect 33232 88256 33284 88262
rect 33232 88198 33284 88204
rect 33060 63566 33180 63594
rect 32956 63504 33008 63510
rect 32956 63446 33008 63452
rect 32968 62830 32996 63446
rect 33060 63034 33088 63566
rect 33140 63436 33192 63442
rect 33140 63378 33192 63384
rect 33048 63028 33100 63034
rect 33048 62970 33100 62976
rect 33048 62892 33100 62898
rect 33048 62834 33100 62840
rect 32956 62824 33008 62830
rect 32956 62766 33008 62772
rect 32968 62490 32996 62766
rect 32956 62484 33008 62490
rect 32956 62426 33008 62432
rect 33060 62354 33088 62834
rect 33048 62348 33100 62354
rect 33048 62290 33100 62296
rect 32956 56500 33008 56506
rect 32956 56442 33008 56448
rect 32864 51060 32916 51066
rect 32588 50176 32640 50182
rect 32588 50118 32640 50124
rect 32600 45778 32628 50118
rect 32692 45898 32720 51046
rect 32864 51002 32916 51008
rect 32772 50788 32824 50794
rect 32772 50730 32824 50736
rect 32680 45892 32732 45898
rect 32680 45834 32732 45840
rect 32600 45750 32720 45778
rect 32496 43172 32548 43178
rect 32496 43114 32548 43120
rect 32588 41472 32640 41478
rect 32588 41414 32640 41420
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32508 14074 32536 31078
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32496 4276 32548 4282
rect 32496 4218 32548 4224
rect 32508 4078 32536 4218
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32404 3188 32456 3194
rect 32404 3130 32456 3136
rect 32220 2984 32272 2990
rect 32220 2926 32272 2932
rect 32496 2984 32548 2990
rect 32496 2926 32548 2932
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31956 800 31984 2450
rect 32232 800 32260 2926
rect 32508 800 32536 2926
rect 32600 2446 32628 41414
rect 32692 40050 32720 45750
rect 32680 40044 32732 40050
rect 32680 39986 32732 39992
rect 32680 39568 32732 39574
rect 32680 39510 32732 39516
rect 32692 27878 32720 39510
rect 32680 27872 32732 27878
rect 32680 27814 32732 27820
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32692 2582 32720 21354
rect 32784 19310 32812 50730
rect 32864 46164 32916 46170
rect 32864 46106 32916 46112
rect 32876 39098 32904 46106
rect 32968 44538 32996 56442
rect 33048 54528 33100 54534
rect 33048 54470 33100 54476
rect 32956 44532 33008 44538
rect 32956 44474 33008 44480
rect 33060 43110 33088 54470
rect 33048 43104 33100 43110
rect 33048 43046 33100 43052
rect 33048 42288 33100 42294
rect 33048 42230 33100 42236
rect 32956 40384 33008 40390
rect 32956 40326 33008 40332
rect 32864 39092 32916 39098
rect 32864 39034 32916 39040
rect 32864 33108 32916 33114
rect 32864 33050 32916 33056
rect 32772 19304 32824 19310
rect 32772 19246 32824 19252
rect 32876 17882 32904 33050
rect 32968 29782 32996 40326
rect 33060 36378 33088 42230
rect 33048 36372 33100 36378
rect 33048 36314 33100 36320
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 32956 29776 33008 29782
rect 32956 29718 33008 29724
rect 33060 28762 33088 35430
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 33048 4208 33100 4214
rect 33048 4150 33100 4156
rect 33060 3534 33088 4150
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33152 3194 33180 63378
rect 33244 35714 33272 88198
rect 33336 65550 33364 89286
rect 33428 85338 33456 114922
rect 33520 112962 33548 119200
rect 33600 116544 33652 116550
rect 33600 116486 33652 116492
rect 33612 113490 33640 116486
rect 33704 113966 33732 119200
rect 33876 116204 33928 116210
rect 33876 116146 33928 116152
rect 33784 115660 33836 115666
rect 33784 115602 33836 115608
rect 33692 113960 33744 113966
rect 33692 113902 33744 113908
rect 33600 113484 33652 113490
rect 33600 113426 33652 113432
rect 33520 112934 33640 112962
rect 33612 112878 33640 112934
rect 33600 112872 33652 112878
rect 33600 112814 33652 112820
rect 33796 111450 33824 115602
rect 33888 113082 33916 116146
rect 33980 115054 34008 119200
rect 34164 117434 34192 119200
rect 34152 117428 34204 117434
rect 34152 117370 34204 117376
rect 34348 117298 34376 119200
rect 34518 118008 34574 118017
rect 34518 117943 34574 117952
rect 34336 117292 34388 117298
rect 34336 117234 34388 117240
rect 34244 117156 34296 117162
rect 34244 117098 34296 117104
rect 34060 116068 34112 116074
rect 34060 116010 34112 116016
rect 33968 115048 34020 115054
rect 33968 114990 34020 114996
rect 33968 114028 34020 114034
rect 33968 113970 34020 113976
rect 33876 113076 33928 113082
rect 33876 113018 33928 113024
rect 33980 111794 34008 113970
rect 34072 113830 34100 116010
rect 34152 114640 34204 114646
rect 34152 114582 34204 114588
rect 34060 113824 34112 113830
rect 34060 113766 34112 113772
rect 33888 111766 34008 111794
rect 33784 111444 33836 111450
rect 33784 111386 33836 111392
rect 33888 109034 33916 111766
rect 33796 109006 33916 109034
rect 33600 99748 33652 99754
rect 33600 99690 33652 99696
rect 33508 97504 33560 97510
rect 33508 97446 33560 97452
rect 33416 85332 33468 85338
rect 33416 85274 33468 85280
rect 33416 85196 33468 85202
rect 33416 85138 33468 85144
rect 33324 65544 33376 65550
rect 33324 65486 33376 65492
rect 33324 63844 33376 63850
rect 33324 63786 33376 63792
rect 33336 55894 33364 63786
rect 33324 55888 33376 55894
rect 33324 55830 33376 55836
rect 33324 51264 33376 51270
rect 33324 51206 33376 51212
rect 33336 47258 33364 51206
rect 33324 47252 33376 47258
rect 33324 47194 33376 47200
rect 33324 47116 33376 47122
rect 33324 47058 33376 47064
rect 33336 45626 33364 47058
rect 33324 45620 33376 45626
rect 33324 45562 33376 45568
rect 33322 44432 33378 44441
rect 33322 44367 33324 44376
rect 33376 44367 33378 44376
rect 33324 44338 33376 44344
rect 33324 42220 33376 42226
rect 33324 42162 33376 42168
rect 33336 35834 33364 42162
rect 33324 35828 33376 35834
rect 33324 35770 33376 35776
rect 33244 35686 33364 35714
rect 33232 35624 33284 35630
rect 33232 35566 33284 35572
rect 33244 25974 33272 35566
rect 33336 35562 33364 35686
rect 33324 35556 33376 35562
rect 33324 35498 33376 35504
rect 33322 35456 33378 35465
rect 33322 35391 33378 35400
rect 33336 31822 33364 35391
rect 33324 31816 33376 31822
rect 33324 31758 33376 31764
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 33428 21418 33456 85138
rect 33520 81326 33548 97446
rect 33508 81320 33560 81326
rect 33508 81262 33560 81268
rect 33508 67652 33560 67658
rect 33508 67594 33560 67600
rect 33520 63442 33548 67594
rect 33508 63436 33560 63442
rect 33508 63378 33560 63384
rect 33508 55888 33560 55894
rect 33508 55830 33560 55836
rect 33416 21412 33468 21418
rect 33416 21354 33468 21360
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 33244 4078 33272 4626
rect 33324 4548 33376 4554
rect 33324 4490 33376 4496
rect 33232 4072 33284 4078
rect 33232 4014 33284 4020
rect 33336 4010 33364 4490
rect 33324 4004 33376 4010
rect 33324 3946 33376 3952
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33244 3534 33272 3878
rect 33520 3738 33548 55830
rect 33612 30394 33640 99690
rect 33692 89684 33744 89690
rect 33692 89626 33744 89632
rect 33704 86086 33732 89626
rect 33692 86080 33744 86086
rect 33692 86022 33744 86028
rect 33692 84040 33744 84046
rect 33692 83982 33744 83988
rect 33704 81025 33732 83982
rect 33690 81016 33746 81025
rect 33690 80951 33746 80960
rect 33692 71528 33744 71534
rect 33692 71470 33744 71476
rect 33600 30388 33652 30394
rect 33600 30330 33652 30336
rect 33704 17746 33732 71470
rect 33796 62422 33824 109006
rect 34164 108338 34192 114582
rect 34256 112742 34284 117098
rect 34532 115734 34560 117943
rect 34624 116890 34652 119200
rect 34702 118824 34758 118833
rect 34702 118759 34758 118768
rect 34612 116884 34664 116890
rect 34716 116872 34744 118759
rect 34808 117178 34836 119200
rect 34992 117858 35020 119200
rect 35268 117978 35296 119200
rect 35256 117972 35308 117978
rect 35256 117914 35308 117920
rect 34992 117830 35388 117858
rect 35256 117700 35308 117706
rect 35256 117642 35308 117648
rect 34940 117532 35236 117552
rect 34996 117530 35020 117532
rect 35076 117530 35100 117532
rect 35156 117530 35180 117532
rect 35018 117478 35020 117530
rect 35082 117478 35094 117530
rect 35156 117478 35158 117530
rect 34996 117476 35020 117478
rect 35076 117476 35100 117478
rect 35156 117476 35180 117478
rect 34940 117456 35236 117476
rect 34980 117224 35032 117230
rect 34808 117150 34928 117178
rect 34980 117166 35032 117172
rect 34900 116890 34928 117150
rect 34888 116884 34940 116890
rect 34716 116844 34836 116872
rect 34612 116826 34664 116832
rect 34704 116748 34756 116754
rect 34704 116690 34756 116696
rect 34612 116680 34664 116686
rect 34612 116622 34664 116628
rect 34520 115728 34572 115734
rect 34520 115670 34572 115676
rect 34336 115660 34388 115666
rect 34336 115602 34388 115608
rect 34244 112736 34296 112742
rect 34244 112678 34296 112684
rect 34072 108310 34192 108338
rect 33968 89548 34020 89554
rect 33968 89490 34020 89496
rect 33980 88466 34008 89490
rect 33968 88460 34020 88466
rect 33968 88402 34020 88408
rect 33980 87854 34008 88402
rect 33968 87848 34020 87854
rect 33968 87790 34020 87796
rect 33968 87508 34020 87514
rect 33968 87450 34020 87456
rect 33980 87310 34008 87450
rect 33968 87304 34020 87310
rect 33968 87246 34020 87252
rect 33966 87000 34022 87009
rect 33966 86935 33968 86944
rect 34020 86935 34022 86944
rect 33968 86906 34020 86912
rect 33968 86760 34020 86766
rect 33968 86702 34020 86708
rect 33980 85678 34008 86702
rect 33968 85672 34020 85678
rect 33968 85614 34020 85620
rect 33876 85536 33928 85542
rect 33876 85478 33928 85484
rect 33888 82074 33916 85478
rect 33968 84720 34020 84726
rect 33968 84662 34020 84668
rect 33876 82068 33928 82074
rect 33876 82010 33928 82016
rect 33980 81705 34008 84662
rect 33966 81696 34022 81705
rect 33966 81631 34022 81640
rect 33968 75744 34020 75750
rect 33968 75686 34020 75692
rect 33980 71738 34008 75686
rect 33968 71732 34020 71738
rect 33968 71674 34020 71680
rect 34072 68950 34100 108310
rect 34152 105120 34204 105126
rect 34152 105062 34204 105068
rect 34164 89554 34192 105062
rect 34244 104168 34296 104174
rect 34244 104110 34296 104116
rect 34152 89548 34204 89554
rect 34152 89490 34204 89496
rect 34256 88466 34284 104110
rect 34244 88460 34296 88466
rect 34244 88402 34296 88408
rect 34152 87848 34204 87854
rect 34152 87790 34204 87796
rect 34164 85814 34192 87790
rect 34244 86624 34296 86630
rect 34244 86566 34296 86572
rect 34152 85808 34204 85814
rect 34152 85750 34204 85756
rect 34256 84640 34284 86566
rect 34164 84612 34284 84640
rect 34164 82414 34192 84612
rect 34244 84516 34296 84522
rect 34244 84458 34296 84464
rect 34256 83502 34284 84458
rect 34244 83496 34296 83502
rect 34244 83438 34296 83444
rect 34152 82408 34204 82414
rect 34152 82350 34204 82356
rect 34060 68944 34112 68950
rect 34060 68886 34112 68892
rect 34060 65544 34112 65550
rect 34060 65486 34112 65492
rect 33876 65136 33928 65142
rect 33876 65078 33928 65084
rect 33888 63594 33916 65078
rect 33968 64456 34020 64462
rect 33968 64398 34020 64404
rect 33980 63986 34008 64398
rect 33968 63980 34020 63986
rect 33968 63922 34020 63928
rect 33888 63566 34008 63594
rect 33876 63436 33928 63442
rect 33876 63378 33928 63384
rect 33784 62416 33836 62422
rect 33784 62358 33836 62364
rect 33888 62234 33916 63378
rect 33980 62694 34008 63566
rect 33968 62688 34020 62694
rect 33968 62630 34020 62636
rect 33796 62206 33916 62234
rect 33692 17740 33744 17746
rect 33692 17682 33744 17688
rect 33600 5024 33652 5030
rect 33600 4966 33652 4972
rect 33612 4010 33640 4966
rect 33600 4004 33652 4010
rect 33600 3946 33652 3952
rect 33508 3732 33560 3738
rect 33508 3674 33560 3680
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 33140 3188 33192 3194
rect 33140 3130 33192 3136
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 32772 2508 32824 2514
rect 32772 2450 32824 2456
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 32784 800 32812 2450
rect 33060 800 33088 2926
rect 33336 800 33364 3538
rect 33690 2816 33746 2825
rect 33690 2751 33746 2760
rect 33704 800 33732 2751
rect 33796 2650 33824 62206
rect 33876 62144 33928 62150
rect 33876 62086 33928 62092
rect 33888 3194 33916 62086
rect 33968 58948 34020 58954
rect 33968 58890 34020 58896
rect 33980 53786 34008 58890
rect 34072 56234 34100 65486
rect 34152 65000 34204 65006
rect 34152 64942 34204 64948
rect 34164 64122 34192 64942
rect 34244 64524 34296 64530
rect 34244 64466 34296 64472
rect 34152 64116 34204 64122
rect 34152 64058 34204 64064
rect 34152 63912 34204 63918
rect 34152 63854 34204 63860
rect 34164 62898 34192 63854
rect 34152 62892 34204 62898
rect 34152 62834 34204 62840
rect 34152 62688 34204 62694
rect 34152 62630 34204 62636
rect 34060 56228 34112 56234
rect 34060 56170 34112 56176
rect 34060 55888 34112 55894
rect 34060 55830 34112 55836
rect 33968 53780 34020 53786
rect 33968 53722 34020 53728
rect 34072 53038 34100 55830
rect 34060 53032 34112 53038
rect 34060 52974 34112 52980
rect 34164 51074 34192 62630
rect 33980 51046 34192 51074
rect 33980 45830 34008 51046
rect 34060 49836 34112 49842
rect 34060 49778 34112 49784
rect 34072 47190 34100 49778
rect 34152 49632 34204 49638
rect 34152 49574 34204 49580
rect 34060 47184 34112 47190
rect 34060 47126 34112 47132
rect 34060 47048 34112 47054
rect 34060 46990 34112 46996
rect 33968 45824 34020 45830
rect 33968 45766 34020 45772
rect 33968 45620 34020 45626
rect 33968 45562 34020 45568
rect 33980 40458 34008 45562
rect 34072 41274 34100 46990
rect 34164 43994 34192 49574
rect 34152 43988 34204 43994
rect 34152 43930 34204 43936
rect 34152 42900 34204 42906
rect 34152 42842 34204 42848
rect 34060 41268 34112 41274
rect 34060 41210 34112 41216
rect 34164 41002 34192 42842
rect 34152 40996 34204 41002
rect 34152 40938 34204 40944
rect 34060 40724 34112 40730
rect 34060 40666 34112 40672
rect 33968 40452 34020 40458
rect 33968 40394 34020 40400
rect 33968 35828 34020 35834
rect 33968 35770 34020 35776
rect 33980 33114 34008 35770
rect 33968 33108 34020 33114
rect 33968 33050 34020 33056
rect 33968 32972 34020 32978
rect 33968 32914 34020 32920
rect 33980 27402 34008 32914
rect 34072 30938 34100 40666
rect 34150 39536 34206 39545
rect 34150 39471 34206 39480
rect 34164 32978 34192 39471
rect 34152 32972 34204 32978
rect 34152 32914 34204 32920
rect 34152 31884 34204 31890
rect 34152 31826 34204 31832
rect 34164 31754 34192 31826
rect 34152 31748 34204 31754
rect 34152 31690 34204 31696
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 34060 30660 34112 30666
rect 34060 30602 34112 30608
rect 33968 27396 34020 27402
rect 33968 27338 34020 27344
rect 34072 22506 34100 30602
rect 34152 26852 34204 26858
rect 34152 26794 34204 26800
rect 34164 23322 34192 26794
rect 34152 23316 34204 23322
rect 34152 23258 34204 23264
rect 34060 22500 34112 22506
rect 34060 22442 34112 22448
rect 34256 3738 34284 64466
rect 34348 58954 34376 115602
rect 34520 115592 34572 115598
rect 34520 115534 34572 115540
rect 34532 115190 34560 115534
rect 34520 115184 34572 115190
rect 34520 115126 34572 115132
rect 34520 114980 34572 114986
rect 34520 114922 34572 114928
rect 34532 113608 34560 114922
rect 34440 113580 34560 113608
rect 34440 112266 34468 113580
rect 34520 113484 34572 113490
rect 34520 113426 34572 113432
rect 34428 112260 34480 112266
rect 34428 112202 34480 112208
rect 34532 111382 34560 113426
rect 34520 111376 34572 111382
rect 34520 111318 34572 111324
rect 34624 111194 34652 116622
rect 34532 111166 34652 111194
rect 34428 99748 34480 99754
rect 34428 99690 34480 99696
rect 34336 58948 34388 58954
rect 34336 58890 34388 58896
rect 34336 58608 34388 58614
rect 34336 58550 34388 58556
rect 34348 54874 34376 58550
rect 34336 54868 34388 54874
rect 34336 54810 34388 54816
rect 34336 52012 34388 52018
rect 34336 51954 34388 51960
rect 34348 50998 34376 51954
rect 34336 50992 34388 50998
rect 34336 50934 34388 50940
rect 34336 49904 34388 49910
rect 34336 49846 34388 49852
rect 34348 43994 34376 49846
rect 34336 43988 34388 43994
rect 34336 43930 34388 43936
rect 34336 40928 34388 40934
rect 34336 40870 34388 40876
rect 34348 39001 34376 40870
rect 34334 38992 34390 39001
rect 34334 38927 34390 38936
rect 34334 38720 34390 38729
rect 34334 38655 34390 38664
rect 34348 35465 34376 38655
rect 34334 35456 34390 35465
rect 34334 35391 34390 35400
rect 34336 31816 34388 31822
rect 34336 31758 34388 31764
rect 34348 17270 34376 31758
rect 34440 18086 34468 99690
rect 34532 63510 34560 111166
rect 34612 111104 34664 111110
rect 34612 111046 34664 111052
rect 34624 87378 34652 111046
rect 34612 87372 34664 87378
rect 34612 87314 34664 87320
rect 34716 87281 34744 116690
rect 34808 116192 34836 116844
rect 34888 116826 34940 116832
rect 34992 116822 35020 117166
rect 34980 116816 35032 116822
rect 34980 116758 35032 116764
rect 34940 116444 35236 116464
rect 34996 116442 35020 116444
rect 35076 116442 35100 116444
rect 35156 116442 35180 116444
rect 35018 116390 35020 116442
rect 35082 116390 35094 116442
rect 35156 116390 35158 116442
rect 34996 116388 35020 116390
rect 35076 116388 35100 116390
rect 35156 116388 35180 116390
rect 34940 116368 35236 116388
rect 35268 116346 35296 117642
rect 35360 116822 35388 117830
rect 35348 116816 35400 116822
rect 35348 116758 35400 116764
rect 35452 116550 35480 119200
rect 35636 117314 35664 119200
rect 35636 117286 35756 117314
rect 35624 117156 35676 117162
rect 35624 117098 35676 117104
rect 35532 116680 35584 116686
rect 35532 116622 35584 116628
rect 35440 116544 35492 116550
rect 35440 116486 35492 116492
rect 35256 116340 35308 116346
rect 35256 116282 35308 116288
rect 35346 116240 35402 116249
rect 34808 116164 34928 116192
rect 35346 116175 35402 116184
rect 34900 115598 34928 116164
rect 35256 116068 35308 116074
rect 35256 116010 35308 116016
rect 34888 115592 34940 115598
rect 34888 115534 34940 115540
rect 34940 115356 35236 115376
rect 34996 115354 35020 115356
rect 35076 115354 35100 115356
rect 35156 115354 35180 115356
rect 35018 115302 35020 115354
rect 35082 115302 35094 115354
rect 35156 115302 35158 115354
rect 34996 115300 35020 115302
rect 35076 115300 35100 115302
rect 35156 115300 35180 115302
rect 34940 115280 35236 115300
rect 35072 115048 35124 115054
rect 35072 114990 35124 114996
rect 34796 114572 34848 114578
rect 34796 114514 34848 114520
rect 34702 87272 34758 87281
rect 34612 87236 34664 87242
rect 34702 87207 34758 87216
rect 34612 87178 34664 87184
rect 34624 64666 34652 87178
rect 34702 87000 34758 87009
rect 34702 86935 34758 86944
rect 34716 67658 34744 86935
rect 34704 67652 34756 67658
rect 34704 67594 34756 67600
rect 34704 65612 34756 65618
rect 34704 65554 34756 65560
rect 34612 64660 34664 64666
rect 34612 64602 34664 64608
rect 34612 63776 34664 63782
rect 34612 63718 34664 63724
rect 34520 63504 34572 63510
rect 34520 63446 34572 63452
rect 34520 56976 34572 56982
rect 34520 56918 34572 56924
rect 34532 52426 34560 56918
rect 34520 52420 34572 52426
rect 34520 52362 34572 52368
rect 34520 50244 34572 50250
rect 34520 50186 34572 50192
rect 34532 45082 34560 50186
rect 34624 48754 34652 63718
rect 34716 63238 34744 65554
rect 34808 65482 34836 114514
rect 35084 114510 35112 114990
rect 35072 114504 35124 114510
rect 35072 114446 35124 114452
rect 34940 114268 35236 114288
rect 34996 114266 35020 114268
rect 35076 114266 35100 114268
rect 35156 114266 35180 114268
rect 35018 114214 35020 114266
rect 35082 114214 35094 114266
rect 35156 114214 35158 114266
rect 34996 114212 35020 114214
rect 35076 114212 35100 114214
rect 35156 114212 35180 114214
rect 34940 114192 35236 114212
rect 34940 113180 35236 113200
rect 34996 113178 35020 113180
rect 35076 113178 35100 113180
rect 35156 113178 35180 113180
rect 35018 113126 35020 113178
rect 35082 113126 35094 113178
rect 35156 113126 35158 113178
rect 34996 113124 35020 113126
rect 35076 113124 35100 113126
rect 35156 113124 35180 113126
rect 34940 113104 35236 113124
rect 34940 112092 35236 112112
rect 34996 112090 35020 112092
rect 35076 112090 35100 112092
rect 35156 112090 35180 112092
rect 35018 112038 35020 112090
rect 35082 112038 35094 112090
rect 35156 112038 35158 112090
rect 34996 112036 35020 112038
rect 35076 112036 35100 112038
rect 35156 112036 35180 112038
rect 34940 112016 35236 112036
rect 34940 111004 35236 111024
rect 34996 111002 35020 111004
rect 35076 111002 35100 111004
rect 35156 111002 35180 111004
rect 35018 110950 35020 111002
rect 35082 110950 35094 111002
rect 35156 110950 35158 111002
rect 34996 110948 35020 110950
rect 35076 110948 35100 110950
rect 35156 110948 35180 110950
rect 34940 110928 35236 110948
rect 34940 109916 35236 109936
rect 34996 109914 35020 109916
rect 35076 109914 35100 109916
rect 35156 109914 35180 109916
rect 35018 109862 35020 109914
rect 35082 109862 35094 109914
rect 35156 109862 35158 109914
rect 34996 109860 35020 109862
rect 35076 109860 35100 109862
rect 35156 109860 35180 109862
rect 34940 109840 35236 109860
rect 34940 108828 35236 108848
rect 34996 108826 35020 108828
rect 35076 108826 35100 108828
rect 35156 108826 35180 108828
rect 35018 108774 35020 108826
rect 35082 108774 35094 108826
rect 35156 108774 35158 108826
rect 34996 108772 35020 108774
rect 35076 108772 35100 108774
rect 35156 108772 35180 108774
rect 34940 108752 35236 108772
rect 34940 107740 35236 107760
rect 34996 107738 35020 107740
rect 35076 107738 35100 107740
rect 35156 107738 35180 107740
rect 35018 107686 35020 107738
rect 35082 107686 35094 107738
rect 35156 107686 35158 107738
rect 34996 107684 35020 107686
rect 35076 107684 35100 107686
rect 35156 107684 35180 107686
rect 34940 107664 35236 107684
rect 34940 106652 35236 106672
rect 34996 106650 35020 106652
rect 35076 106650 35100 106652
rect 35156 106650 35180 106652
rect 35018 106598 35020 106650
rect 35082 106598 35094 106650
rect 35156 106598 35158 106650
rect 34996 106596 35020 106598
rect 35076 106596 35100 106598
rect 35156 106596 35180 106598
rect 34940 106576 35236 106596
rect 34940 105564 35236 105584
rect 34996 105562 35020 105564
rect 35076 105562 35100 105564
rect 35156 105562 35180 105564
rect 35018 105510 35020 105562
rect 35082 105510 35094 105562
rect 35156 105510 35158 105562
rect 34996 105508 35020 105510
rect 35076 105508 35100 105510
rect 35156 105508 35180 105510
rect 34940 105488 35236 105508
rect 34940 104476 35236 104496
rect 34996 104474 35020 104476
rect 35076 104474 35100 104476
rect 35156 104474 35180 104476
rect 35018 104422 35020 104474
rect 35082 104422 35094 104474
rect 35156 104422 35158 104474
rect 34996 104420 35020 104422
rect 35076 104420 35100 104422
rect 35156 104420 35180 104422
rect 34940 104400 35236 104420
rect 34940 103388 35236 103408
rect 34996 103386 35020 103388
rect 35076 103386 35100 103388
rect 35156 103386 35180 103388
rect 35018 103334 35020 103386
rect 35082 103334 35094 103386
rect 35156 103334 35158 103386
rect 34996 103332 35020 103334
rect 35076 103332 35100 103334
rect 35156 103332 35180 103334
rect 34940 103312 35236 103332
rect 34940 102300 35236 102320
rect 34996 102298 35020 102300
rect 35076 102298 35100 102300
rect 35156 102298 35180 102300
rect 35018 102246 35020 102298
rect 35082 102246 35094 102298
rect 35156 102246 35158 102298
rect 34996 102244 35020 102246
rect 35076 102244 35100 102246
rect 35156 102244 35180 102246
rect 34940 102224 35236 102244
rect 34940 101212 35236 101232
rect 34996 101210 35020 101212
rect 35076 101210 35100 101212
rect 35156 101210 35180 101212
rect 35018 101158 35020 101210
rect 35082 101158 35094 101210
rect 35156 101158 35158 101210
rect 34996 101156 35020 101158
rect 35076 101156 35100 101158
rect 35156 101156 35180 101158
rect 34940 101136 35236 101156
rect 34940 100124 35236 100144
rect 34996 100122 35020 100124
rect 35076 100122 35100 100124
rect 35156 100122 35180 100124
rect 35018 100070 35020 100122
rect 35082 100070 35094 100122
rect 35156 100070 35158 100122
rect 34996 100068 35020 100070
rect 35076 100068 35100 100070
rect 35156 100068 35180 100070
rect 34940 100048 35236 100068
rect 34940 99036 35236 99056
rect 34996 99034 35020 99036
rect 35076 99034 35100 99036
rect 35156 99034 35180 99036
rect 35018 98982 35020 99034
rect 35082 98982 35094 99034
rect 35156 98982 35158 99034
rect 34996 98980 35020 98982
rect 35076 98980 35100 98982
rect 35156 98980 35180 98982
rect 34940 98960 35236 98980
rect 34940 97948 35236 97968
rect 34996 97946 35020 97948
rect 35076 97946 35100 97948
rect 35156 97946 35180 97948
rect 35018 97894 35020 97946
rect 35082 97894 35094 97946
rect 35156 97894 35158 97946
rect 34996 97892 35020 97894
rect 35076 97892 35100 97894
rect 35156 97892 35180 97894
rect 34940 97872 35236 97892
rect 34940 96860 35236 96880
rect 34996 96858 35020 96860
rect 35076 96858 35100 96860
rect 35156 96858 35180 96860
rect 35018 96806 35020 96858
rect 35082 96806 35094 96858
rect 35156 96806 35158 96858
rect 34996 96804 35020 96806
rect 35076 96804 35100 96806
rect 35156 96804 35180 96806
rect 34940 96784 35236 96804
rect 34940 95772 35236 95792
rect 34996 95770 35020 95772
rect 35076 95770 35100 95772
rect 35156 95770 35180 95772
rect 35018 95718 35020 95770
rect 35082 95718 35094 95770
rect 35156 95718 35158 95770
rect 34996 95716 35020 95718
rect 35076 95716 35100 95718
rect 35156 95716 35180 95718
rect 34940 95696 35236 95716
rect 34940 94684 35236 94704
rect 34996 94682 35020 94684
rect 35076 94682 35100 94684
rect 35156 94682 35180 94684
rect 35018 94630 35020 94682
rect 35082 94630 35094 94682
rect 35156 94630 35158 94682
rect 34996 94628 35020 94630
rect 35076 94628 35100 94630
rect 35156 94628 35180 94630
rect 34940 94608 35236 94628
rect 34940 93596 35236 93616
rect 34996 93594 35020 93596
rect 35076 93594 35100 93596
rect 35156 93594 35180 93596
rect 35018 93542 35020 93594
rect 35082 93542 35094 93594
rect 35156 93542 35158 93594
rect 34996 93540 35020 93542
rect 35076 93540 35100 93542
rect 35156 93540 35180 93542
rect 34940 93520 35236 93540
rect 34940 92508 35236 92528
rect 34996 92506 35020 92508
rect 35076 92506 35100 92508
rect 35156 92506 35180 92508
rect 35018 92454 35020 92506
rect 35082 92454 35094 92506
rect 35156 92454 35158 92506
rect 34996 92452 35020 92454
rect 35076 92452 35100 92454
rect 35156 92452 35180 92454
rect 34940 92432 35236 92452
rect 34940 91420 35236 91440
rect 34996 91418 35020 91420
rect 35076 91418 35100 91420
rect 35156 91418 35180 91420
rect 35018 91366 35020 91418
rect 35082 91366 35094 91418
rect 35156 91366 35158 91418
rect 34996 91364 35020 91366
rect 35076 91364 35100 91366
rect 35156 91364 35180 91366
rect 34940 91344 35236 91364
rect 34940 90332 35236 90352
rect 34996 90330 35020 90332
rect 35076 90330 35100 90332
rect 35156 90330 35180 90332
rect 35018 90278 35020 90330
rect 35082 90278 35094 90330
rect 35156 90278 35158 90330
rect 34996 90276 35020 90278
rect 35076 90276 35100 90278
rect 35156 90276 35180 90278
rect 34940 90256 35236 90276
rect 34940 89244 35236 89264
rect 34996 89242 35020 89244
rect 35076 89242 35100 89244
rect 35156 89242 35180 89244
rect 35018 89190 35020 89242
rect 35082 89190 35094 89242
rect 35156 89190 35158 89242
rect 34996 89188 35020 89190
rect 35076 89188 35100 89190
rect 35156 89188 35180 89190
rect 34940 89168 35236 89188
rect 34940 88156 35236 88176
rect 34996 88154 35020 88156
rect 35076 88154 35100 88156
rect 35156 88154 35180 88156
rect 35018 88102 35020 88154
rect 35082 88102 35094 88154
rect 35156 88102 35158 88154
rect 34996 88100 35020 88102
rect 35076 88100 35100 88102
rect 35156 88100 35180 88102
rect 34940 88080 35236 88100
rect 35268 87768 35296 116010
rect 35360 115734 35388 116175
rect 35348 115728 35400 115734
rect 35348 115670 35400 115676
rect 35348 115592 35400 115598
rect 35348 115534 35400 115540
rect 35360 114073 35388 115534
rect 35346 114064 35402 114073
rect 35544 114050 35572 116622
rect 35346 113999 35402 114008
rect 35452 114022 35572 114050
rect 35348 113892 35400 113898
rect 35348 113834 35400 113840
rect 35360 104378 35388 113834
rect 35348 104372 35400 104378
rect 35348 104314 35400 104320
rect 35348 101448 35400 101454
rect 35348 101390 35400 101396
rect 35176 87740 35296 87768
rect 35176 87242 35204 87740
rect 35360 87666 35388 101390
rect 35268 87638 35388 87666
rect 35268 87378 35296 87638
rect 35452 87496 35480 114022
rect 35532 113960 35584 113966
rect 35532 113902 35584 113908
rect 35544 111858 35572 113902
rect 35532 111852 35584 111858
rect 35532 111794 35584 111800
rect 35532 111716 35584 111722
rect 35532 111658 35584 111664
rect 35360 87468 35480 87496
rect 35256 87372 35308 87378
rect 35256 87314 35308 87320
rect 35360 87281 35388 87468
rect 35440 87372 35492 87378
rect 35440 87314 35492 87320
rect 35346 87272 35402 87281
rect 35164 87236 35216 87242
rect 35346 87207 35402 87216
rect 35164 87178 35216 87184
rect 35256 87168 35308 87174
rect 35452 87122 35480 87314
rect 35256 87110 35308 87116
rect 34940 87068 35236 87088
rect 34996 87066 35020 87068
rect 35076 87066 35100 87068
rect 35156 87066 35180 87068
rect 35018 87014 35020 87066
rect 35082 87014 35094 87066
rect 35156 87014 35158 87066
rect 34996 87012 35020 87014
rect 35076 87012 35100 87014
rect 35156 87012 35180 87014
rect 34940 86992 35236 87012
rect 34940 85980 35236 86000
rect 34996 85978 35020 85980
rect 35076 85978 35100 85980
rect 35156 85978 35180 85980
rect 35018 85926 35020 85978
rect 35082 85926 35094 85978
rect 35156 85926 35158 85978
rect 34996 85924 35020 85926
rect 35076 85924 35100 85926
rect 35156 85924 35180 85926
rect 34940 85904 35236 85924
rect 34940 84892 35236 84912
rect 34996 84890 35020 84892
rect 35076 84890 35100 84892
rect 35156 84890 35180 84892
rect 35018 84838 35020 84890
rect 35082 84838 35094 84890
rect 35156 84838 35158 84890
rect 34996 84836 35020 84838
rect 35076 84836 35100 84838
rect 35156 84836 35180 84838
rect 34940 84816 35236 84836
rect 34940 83804 35236 83824
rect 34996 83802 35020 83804
rect 35076 83802 35100 83804
rect 35156 83802 35180 83804
rect 35018 83750 35020 83802
rect 35082 83750 35094 83802
rect 35156 83750 35158 83802
rect 34996 83748 35020 83750
rect 35076 83748 35100 83750
rect 35156 83748 35180 83750
rect 34940 83728 35236 83748
rect 34940 82716 35236 82736
rect 34996 82714 35020 82716
rect 35076 82714 35100 82716
rect 35156 82714 35180 82716
rect 35018 82662 35020 82714
rect 35082 82662 35094 82714
rect 35156 82662 35158 82714
rect 34996 82660 35020 82662
rect 35076 82660 35100 82662
rect 35156 82660 35180 82662
rect 34940 82640 35236 82660
rect 34940 81628 35236 81648
rect 34996 81626 35020 81628
rect 35076 81626 35100 81628
rect 35156 81626 35180 81628
rect 35018 81574 35020 81626
rect 35082 81574 35094 81626
rect 35156 81574 35158 81626
rect 34996 81572 35020 81574
rect 35076 81572 35100 81574
rect 35156 81572 35180 81574
rect 34940 81552 35236 81572
rect 34940 80540 35236 80560
rect 34996 80538 35020 80540
rect 35076 80538 35100 80540
rect 35156 80538 35180 80540
rect 35018 80486 35020 80538
rect 35082 80486 35094 80538
rect 35156 80486 35158 80538
rect 34996 80484 35020 80486
rect 35076 80484 35100 80486
rect 35156 80484 35180 80486
rect 34940 80464 35236 80484
rect 34940 79452 35236 79472
rect 34996 79450 35020 79452
rect 35076 79450 35100 79452
rect 35156 79450 35180 79452
rect 35018 79398 35020 79450
rect 35082 79398 35094 79450
rect 35156 79398 35158 79450
rect 34996 79396 35020 79398
rect 35076 79396 35100 79398
rect 35156 79396 35180 79398
rect 34940 79376 35236 79396
rect 34940 78364 35236 78384
rect 34996 78362 35020 78364
rect 35076 78362 35100 78364
rect 35156 78362 35180 78364
rect 35018 78310 35020 78362
rect 35082 78310 35094 78362
rect 35156 78310 35158 78362
rect 34996 78308 35020 78310
rect 35076 78308 35100 78310
rect 35156 78308 35180 78310
rect 34940 78288 35236 78308
rect 34940 77276 35236 77296
rect 34996 77274 35020 77276
rect 35076 77274 35100 77276
rect 35156 77274 35180 77276
rect 35018 77222 35020 77274
rect 35082 77222 35094 77274
rect 35156 77222 35158 77274
rect 34996 77220 35020 77222
rect 35076 77220 35100 77222
rect 35156 77220 35180 77222
rect 34940 77200 35236 77220
rect 34940 76188 35236 76208
rect 34996 76186 35020 76188
rect 35076 76186 35100 76188
rect 35156 76186 35180 76188
rect 35018 76134 35020 76186
rect 35082 76134 35094 76186
rect 35156 76134 35158 76186
rect 34996 76132 35020 76134
rect 35076 76132 35100 76134
rect 35156 76132 35180 76134
rect 34940 76112 35236 76132
rect 34940 75100 35236 75120
rect 34996 75098 35020 75100
rect 35076 75098 35100 75100
rect 35156 75098 35180 75100
rect 35018 75046 35020 75098
rect 35082 75046 35094 75098
rect 35156 75046 35158 75098
rect 34996 75044 35020 75046
rect 35076 75044 35100 75046
rect 35156 75044 35180 75046
rect 34940 75024 35236 75044
rect 34940 74012 35236 74032
rect 34996 74010 35020 74012
rect 35076 74010 35100 74012
rect 35156 74010 35180 74012
rect 35018 73958 35020 74010
rect 35082 73958 35094 74010
rect 35156 73958 35158 74010
rect 34996 73956 35020 73958
rect 35076 73956 35100 73958
rect 35156 73956 35180 73958
rect 34940 73936 35236 73956
rect 34940 72924 35236 72944
rect 34996 72922 35020 72924
rect 35076 72922 35100 72924
rect 35156 72922 35180 72924
rect 35018 72870 35020 72922
rect 35082 72870 35094 72922
rect 35156 72870 35158 72922
rect 34996 72868 35020 72870
rect 35076 72868 35100 72870
rect 35156 72868 35180 72870
rect 34940 72848 35236 72868
rect 34940 71836 35236 71856
rect 34996 71834 35020 71836
rect 35076 71834 35100 71836
rect 35156 71834 35180 71836
rect 35018 71782 35020 71834
rect 35082 71782 35094 71834
rect 35156 71782 35158 71834
rect 34996 71780 35020 71782
rect 35076 71780 35100 71782
rect 35156 71780 35180 71782
rect 34940 71760 35236 71780
rect 34940 70748 35236 70768
rect 34996 70746 35020 70748
rect 35076 70746 35100 70748
rect 35156 70746 35180 70748
rect 35018 70694 35020 70746
rect 35082 70694 35094 70746
rect 35156 70694 35158 70746
rect 34996 70692 35020 70694
rect 35076 70692 35100 70694
rect 35156 70692 35180 70694
rect 34940 70672 35236 70692
rect 34940 69660 35236 69680
rect 34996 69658 35020 69660
rect 35076 69658 35100 69660
rect 35156 69658 35180 69660
rect 35018 69606 35020 69658
rect 35082 69606 35094 69658
rect 35156 69606 35158 69658
rect 34996 69604 35020 69606
rect 35076 69604 35100 69606
rect 35156 69604 35180 69606
rect 34940 69584 35236 69604
rect 34940 68572 35236 68592
rect 34996 68570 35020 68572
rect 35076 68570 35100 68572
rect 35156 68570 35180 68572
rect 35018 68518 35020 68570
rect 35082 68518 35094 68570
rect 35156 68518 35158 68570
rect 34996 68516 35020 68518
rect 35076 68516 35100 68518
rect 35156 68516 35180 68518
rect 34940 68496 35236 68516
rect 34940 67484 35236 67504
rect 34996 67482 35020 67484
rect 35076 67482 35100 67484
rect 35156 67482 35180 67484
rect 35018 67430 35020 67482
rect 35082 67430 35094 67482
rect 35156 67430 35158 67482
rect 34996 67428 35020 67430
rect 35076 67428 35100 67430
rect 35156 67428 35180 67430
rect 34940 67408 35236 67428
rect 34940 66396 35236 66416
rect 34996 66394 35020 66396
rect 35076 66394 35100 66396
rect 35156 66394 35180 66396
rect 35018 66342 35020 66394
rect 35082 66342 35094 66394
rect 35156 66342 35158 66394
rect 34996 66340 35020 66342
rect 35076 66340 35100 66342
rect 35156 66340 35180 66342
rect 34940 66320 35236 66340
rect 34796 65476 34848 65482
rect 34796 65418 34848 65424
rect 34940 65308 35236 65328
rect 34996 65306 35020 65308
rect 35076 65306 35100 65308
rect 35156 65306 35180 65308
rect 35018 65254 35020 65306
rect 35082 65254 35094 65306
rect 35156 65254 35158 65306
rect 34996 65252 35020 65254
rect 35076 65252 35100 65254
rect 35156 65252 35180 65254
rect 34940 65232 35236 65252
rect 35268 65006 35296 87110
rect 35360 87094 35480 87122
rect 35256 65000 35308 65006
rect 35256 64942 35308 64948
rect 34940 64220 35236 64240
rect 34996 64218 35020 64220
rect 35076 64218 35100 64220
rect 35156 64218 35180 64220
rect 35018 64166 35020 64218
rect 35082 64166 35094 64218
rect 35156 64166 35158 64218
rect 34996 64164 35020 64166
rect 35076 64164 35100 64166
rect 35156 64164 35180 64166
rect 34940 64144 35236 64164
rect 34888 63844 34940 63850
rect 34888 63786 34940 63792
rect 34900 63578 34928 63786
rect 34888 63572 34940 63578
rect 34888 63514 34940 63520
rect 35256 63436 35308 63442
rect 35256 63378 35308 63384
rect 34704 63232 34756 63238
rect 34704 63174 34756 63180
rect 34940 63132 35236 63152
rect 34996 63130 35020 63132
rect 35076 63130 35100 63132
rect 35156 63130 35180 63132
rect 35018 63078 35020 63130
rect 35082 63078 35094 63130
rect 35156 63078 35158 63130
rect 34996 63076 35020 63078
rect 35076 63076 35100 63078
rect 35156 63076 35180 63078
rect 34940 63056 35236 63076
rect 35268 62898 35296 63378
rect 34980 62892 35032 62898
rect 34980 62834 35032 62840
rect 35256 62892 35308 62898
rect 35256 62834 35308 62840
rect 34992 62354 35020 62834
rect 35360 62354 35388 87094
rect 35438 87000 35494 87009
rect 35438 86935 35494 86944
rect 35452 63578 35480 86935
rect 35544 65618 35572 111658
rect 35636 99958 35664 117098
rect 35728 116278 35756 117286
rect 35716 116272 35768 116278
rect 35716 116214 35768 116220
rect 35716 116136 35768 116142
rect 35716 116078 35768 116084
rect 35728 113778 35756 116078
rect 35820 115802 35848 119200
rect 35900 116748 35952 116754
rect 35900 116690 35952 116696
rect 35808 115796 35860 115802
rect 35808 115738 35860 115744
rect 35912 115682 35940 116690
rect 36096 115802 36124 119200
rect 36280 117298 36308 119200
rect 36268 117292 36320 117298
rect 36268 117234 36320 117240
rect 36084 115796 36136 115802
rect 36084 115738 36136 115744
rect 35820 115654 35940 115682
rect 36268 115660 36320 115666
rect 35820 114034 35848 115654
rect 36268 115602 36320 115608
rect 35992 114980 36044 114986
rect 35992 114922 36044 114928
rect 35808 114028 35860 114034
rect 35808 113970 35860 113976
rect 35728 113750 35940 113778
rect 35806 113656 35862 113665
rect 35806 113591 35862 113600
rect 35716 113484 35768 113490
rect 35716 113426 35768 113432
rect 35624 99952 35676 99958
rect 35624 99894 35676 99900
rect 35624 98116 35676 98122
rect 35624 98058 35676 98064
rect 35636 87553 35664 98058
rect 35622 87544 35678 87553
rect 35622 87479 35678 87488
rect 35622 87000 35678 87009
rect 35622 86935 35678 86944
rect 35532 65612 35584 65618
rect 35532 65554 35584 65560
rect 35636 65498 35664 86935
rect 35544 65470 35664 65498
rect 35440 63572 35492 63578
rect 35440 63514 35492 63520
rect 34980 62348 35032 62354
rect 34980 62290 35032 62296
rect 35348 62348 35400 62354
rect 35348 62290 35400 62296
rect 34940 62044 35236 62064
rect 34996 62042 35020 62044
rect 35076 62042 35100 62044
rect 35156 62042 35180 62044
rect 35018 61990 35020 62042
rect 35082 61990 35094 62042
rect 35156 61990 35158 62042
rect 34996 61988 35020 61990
rect 35076 61988 35100 61990
rect 35156 61988 35180 61990
rect 34940 61968 35236 61988
rect 35348 61600 35400 61606
rect 35348 61542 35400 61548
rect 34796 61056 34848 61062
rect 34796 60998 34848 61004
rect 34704 57452 34756 57458
rect 34704 57394 34756 57400
rect 34716 53174 34744 57394
rect 34704 53168 34756 53174
rect 34704 53110 34756 53116
rect 34704 53032 34756 53038
rect 34704 52974 34756 52980
rect 34612 48748 34664 48754
rect 34612 48690 34664 48696
rect 34612 48612 34664 48618
rect 34612 48554 34664 48560
rect 34520 45076 34572 45082
rect 34520 45018 34572 45024
rect 34518 44976 34574 44985
rect 34518 44911 34520 44920
rect 34572 44911 34574 44920
rect 34520 44882 34572 44888
rect 34624 44538 34652 48554
rect 34612 44532 34664 44538
rect 34612 44474 34664 44480
rect 34520 43376 34572 43382
rect 34520 43318 34572 43324
rect 34532 39624 34560 43318
rect 34612 43172 34664 43178
rect 34612 43114 34664 43120
rect 34624 41818 34652 43114
rect 34612 41812 34664 41818
rect 34612 41754 34664 41760
rect 34610 41168 34666 41177
rect 34610 41103 34666 41112
rect 34624 41070 34652 41103
rect 34612 41064 34664 41070
rect 34612 41006 34664 41012
rect 34612 39976 34664 39982
rect 34612 39918 34664 39924
rect 34624 39817 34652 39918
rect 34610 39808 34666 39817
rect 34610 39743 34666 39752
rect 34532 39596 34652 39624
rect 34520 39500 34572 39506
rect 34520 39442 34572 39448
rect 34532 39409 34560 39442
rect 34518 39400 34574 39409
rect 34518 39335 34574 39344
rect 34520 38820 34572 38826
rect 34520 38762 34572 38768
rect 34532 36038 34560 38762
rect 34624 38554 34652 39596
rect 34612 38548 34664 38554
rect 34612 38490 34664 38496
rect 34612 38276 34664 38282
rect 34612 38218 34664 38224
rect 34624 36038 34652 38218
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34624 35222 34652 35974
rect 34612 35216 34664 35222
rect 34612 35158 34664 35164
rect 34520 35148 34572 35154
rect 34520 35090 34572 35096
rect 34532 31890 34560 35090
rect 34610 34640 34666 34649
rect 34610 34575 34666 34584
rect 34624 34542 34652 34575
rect 34612 34536 34664 34542
rect 34612 34478 34664 34484
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34520 30864 34572 30870
rect 34520 30806 34572 30812
rect 34532 29170 34560 30806
rect 34612 30388 34664 30394
rect 34612 30330 34664 30336
rect 34624 30138 34652 30330
rect 34716 30258 34744 52974
rect 34808 42276 34836 60998
rect 34940 60956 35236 60976
rect 34996 60954 35020 60956
rect 35076 60954 35100 60956
rect 35156 60954 35180 60956
rect 35018 60902 35020 60954
rect 35082 60902 35094 60954
rect 35156 60902 35158 60954
rect 34996 60900 35020 60902
rect 35076 60900 35100 60902
rect 35156 60900 35180 60902
rect 34940 60880 35236 60900
rect 34940 59868 35236 59888
rect 34996 59866 35020 59868
rect 35076 59866 35100 59868
rect 35156 59866 35180 59868
rect 35018 59814 35020 59866
rect 35082 59814 35094 59866
rect 35156 59814 35158 59866
rect 34996 59812 35020 59814
rect 35076 59812 35100 59814
rect 35156 59812 35180 59814
rect 34940 59792 35236 59812
rect 35256 58948 35308 58954
rect 35256 58890 35308 58896
rect 34940 58780 35236 58800
rect 34996 58778 35020 58780
rect 35076 58778 35100 58780
rect 35156 58778 35180 58780
rect 35018 58726 35020 58778
rect 35082 58726 35094 58778
rect 35156 58726 35158 58778
rect 34996 58724 35020 58726
rect 35076 58724 35100 58726
rect 35156 58724 35180 58726
rect 34940 58704 35236 58724
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 35268 55894 35296 58890
rect 35256 55888 35308 55894
rect 34886 55856 34942 55865
rect 35256 55830 35308 55836
rect 34886 55791 34888 55800
rect 34940 55791 34942 55800
rect 34888 55762 34940 55768
rect 35256 55616 35308 55622
rect 35256 55558 35308 55564
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 35164 55072 35216 55078
rect 35164 55014 35216 55020
rect 35176 54602 35204 55014
rect 35164 54596 35216 54602
rect 35164 54538 35216 54544
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 35164 48748 35216 48754
rect 35164 48690 35216 48696
rect 35176 48142 35204 48690
rect 35164 48136 35216 48142
rect 35164 48078 35216 48084
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 35268 47274 35296 55558
rect 35360 47410 35388 61542
rect 35438 55448 35494 55457
rect 35438 55383 35494 55392
rect 35452 55214 35480 55383
rect 35440 55208 35492 55214
rect 35440 55150 35492 55156
rect 35440 55072 35492 55078
rect 35440 55014 35492 55020
rect 35452 53990 35480 55014
rect 35440 53984 35492 53990
rect 35440 53926 35492 53932
rect 35440 53100 35492 53106
rect 35440 53042 35492 53048
rect 35452 48074 35480 53042
rect 35544 51542 35572 65470
rect 35728 60858 35756 113426
rect 35820 112538 35848 113591
rect 35808 112532 35860 112538
rect 35808 112474 35860 112480
rect 35808 111852 35860 111858
rect 35808 111794 35860 111800
rect 35820 105738 35848 111794
rect 35912 111110 35940 113750
rect 36004 112470 36032 114922
rect 36176 114572 36228 114578
rect 36176 114514 36228 114520
rect 36084 113484 36136 113490
rect 36084 113426 36136 113432
rect 35992 112464 36044 112470
rect 35992 112406 36044 112412
rect 35900 111104 35952 111110
rect 35900 111046 35952 111052
rect 35808 105732 35860 105738
rect 35808 105674 35860 105680
rect 36096 105466 36124 113426
rect 36188 109750 36216 114514
rect 36280 110770 36308 115602
rect 36372 113558 36400 119575
rect 36450 119200 36506 120800
rect 36634 119232 36690 119241
rect 36464 117094 36492 119200
rect 36726 119200 36782 120800
rect 36910 119200 36966 120800
rect 37094 119200 37150 120800
rect 37370 119200 37426 120800
rect 37554 119200 37610 120800
rect 37738 119200 37794 120800
rect 37922 119200 37978 120800
rect 38198 119200 38254 120800
rect 38382 119200 38438 120800
rect 38566 119200 38622 120800
rect 38842 119200 38898 120800
rect 39026 119200 39082 120800
rect 39210 119200 39266 120800
rect 39486 119200 39542 120800
rect 39670 119200 39726 120800
rect 39854 119200 39910 120800
rect 36634 119167 36690 119176
rect 36544 117292 36596 117298
rect 36544 117234 36596 117240
rect 36556 117201 36584 117234
rect 36542 117192 36598 117201
rect 36542 117127 36598 117136
rect 36452 117088 36504 117094
rect 36452 117030 36504 117036
rect 36648 115954 36676 119167
rect 36556 115926 36676 115954
rect 36360 113552 36412 113558
rect 36360 113494 36412 113500
rect 36556 113082 36584 115926
rect 36636 115660 36688 115666
rect 36636 115602 36688 115608
rect 36544 113076 36596 113082
rect 36544 113018 36596 113024
rect 36360 112804 36412 112810
rect 36360 112746 36412 112752
rect 36268 110764 36320 110770
rect 36268 110706 36320 110712
rect 36176 109744 36228 109750
rect 36176 109686 36228 109692
rect 36084 105460 36136 105466
rect 36084 105402 36136 105408
rect 36084 103148 36136 103154
rect 36084 103090 36136 103096
rect 35992 95600 36044 95606
rect 35992 95542 36044 95548
rect 35900 94512 35952 94518
rect 35900 94454 35952 94460
rect 35808 92336 35860 92342
rect 35808 92278 35860 92284
rect 35820 88806 35848 92278
rect 35912 90234 35940 94454
rect 36004 90710 36032 95542
rect 35992 90704 36044 90710
rect 35992 90646 36044 90652
rect 35900 90228 35952 90234
rect 35900 90170 35952 90176
rect 36096 89714 36124 103090
rect 36176 95872 36228 95878
rect 36176 95814 36228 95820
rect 35912 89686 36124 89714
rect 35808 88800 35860 88806
rect 35808 88742 35860 88748
rect 35808 88528 35860 88534
rect 35808 88470 35860 88476
rect 35820 83366 35848 88470
rect 35912 87854 35940 89686
rect 36188 89570 36216 95814
rect 36372 89714 36400 112746
rect 36542 111480 36598 111489
rect 36542 111415 36544 111424
rect 36596 111415 36598 111424
rect 36544 111386 36596 111392
rect 36452 111308 36504 111314
rect 36452 111250 36504 111256
rect 36464 110906 36492 111250
rect 36452 110900 36504 110906
rect 36452 110842 36504 110848
rect 36452 110764 36504 110770
rect 36452 110706 36504 110712
rect 36004 89542 36216 89570
rect 36280 89686 36400 89714
rect 35900 87848 35952 87854
rect 35900 87790 35952 87796
rect 35900 87712 35952 87718
rect 35900 87654 35952 87660
rect 35912 83978 35940 87654
rect 36004 86358 36032 89542
rect 36084 88800 36136 88806
rect 36084 88742 36136 88748
rect 35992 86352 36044 86358
rect 35992 86294 36044 86300
rect 36096 84794 36124 88742
rect 36176 87984 36228 87990
rect 36176 87926 36228 87932
rect 36084 84788 36136 84794
rect 36084 84730 36136 84736
rect 35900 83972 35952 83978
rect 35900 83914 35952 83920
rect 35808 83360 35860 83366
rect 35808 83302 35860 83308
rect 36188 83162 36216 87926
rect 36176 83156 36228 83162
rect 36176 83098 36228 83104
rect 36280 80054 36308 89686
rect 36360 89480 36412 89486
rect 36360 89422 36412 89428
rect 36372 84046 36400 89422
rect 36360 84040 36412 84046
rect 36360 83982 36412 83988
rect 36360 83904 36412 83910
rect 36360 83846 36412 83852
rect 36188 80026 36308 80054
rect 35900 78464 35952 78470
rect 35900 78406 35952 78412
rect 35912 74474 35940 78406
rect 35992 77988 36044 77994
rect 35992 77930 36044 77936
rect 35820 74446 35940 74474
rect 35716 60852 35768 60858
rect 35716 60794 35768 60800
rect 35820 60734 35848 74446
rect 35636 60706 35848 60734
rect 35532 51536 35584 51542
rect 35532 51478 35584 51484
rect 35532 50924 35584 50930
rect 35532 50866 35584 50872
rect 35544 49434 35572 50866
rect 35532 49428 35584 49434
rect 35532 49370 35584 49376
rect 35636 49298 35664 60706
rect 35900 58676 35952 58682
rect 35900 58618 35952 58624
rect 35808 57044 35860 57050
rect 35808 56986 35860 56992
rect 35820 56302 35848 56986
rect 35808 56296 35860 56302
rect 35808 56238 35860 56244
rect 35716 56228 35768 56234
rect 35716 56170 35768 56176
rect 35728 55282 35756 56170
rect 35716 55276 35768 55282
rect 35716 55218 35768 55224
rect 35806 54904 35862 54913
rect 35806 54839 35862 54848
rect 35716 54732 35768 54738
rect 35716 54674 35768 54680
rect 35728 54097 35756 54674
rect 35820 54126 35848 54839
rect 35912 54262 35940 58618
rect 36004 58478 36032 77930
rect 36084 75812 36136 75818
rect 36084 75754 36136 75760
rect 35992 58472 36044 58478
rect 35992 58414 36044 58420
rect 35992 58336 36044 58342
rect 35992 58278 36044 58284
rect 36004 55214 36032 58278
rect 35992 55208 36044 55214
rect 35992 55150 36044 55156
rect 35992 54664 36044 54670
rect 35992 54606 36044 54612
rect 35900 54256 35952 54262
rect 35900 54198 35952 54204
rect 35808 54120 35860 54126
rect 35714 54088 35770 54097
rect 35808 54062 35860 54068
rect 35714 54023 35770 54032
rect 35716 53984 35768 53990
rect 35716 53926 35768 53932
rect 35900 53984 35952 53990
rect 35900 53926 35952 53932
rect 35728 52714 35756 53926
rect 35808 53032 35860 53038
rect 35808 52974 35860 52980
rect 35820 52873 35848 52974
rect 35806 52864 35862 52873
rect 35806 52799 35862 52808
rect 35728 52686 35848 52714
rect 35820 51074 35848 52686
rect 35728 51046 35848 51074
rect 35912 51074 35940 53926
rect 36004 51610 36032 54606
rect 35992 51604 36044 51610
rect 35992 51546 36044 51552
rect 35912 51046 36032 51074
rect 35728 49638 35756 51046
rect 35900 50992 35952 50998
rect 35900 50934 35952 50940
rect 35808 50380 35860 50386
rect 35808 50322 35860 50328
rect 35820 50289 35848 50322
rect 35806 50280 35862 50289
rect 35806 50215 35862 50224
rect 35716 49632 35768 49638
rect 35716 49574 35768 49580
rect 35716 49360 35768 49366
rect 35716 49302 35768 49308
rect 35624 49292 35676 49298
rect 35624 49234 35676 49240
rect 35624 49156 35676 49162
rect 35624 49098 35676 49104
rect 35530 48920 35586 48929
rect 35530 48855 35586 48864
rect 35544 48210 35572 48855
rect 35532 48204 35584 48210
rect 35532 48146 35584 48152
rect 35440 48068 35492 48074
rect 35440 48010 35492 48016
rect 35360 47382 35572 47410
rect 35268 47246 35388 47274
rect 35256 47116 35308 47122
rect 35256 47058 35308 47064
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 35164 46436 35216 46442
rect 35164 46378 35216 46384
rect 35176 45812 35204 46378
rect 35268 46345 35296 47058
rect 35254 46336 35310 46345
rect 35254 46271 35310 46280
rect 35176 45784 35296 45812
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 35268 44946 35296 45784
rect 35256 44940 35308 44946
rect 35256 44882 35308 44888
rect 35360 44690 35388 47246
rect 35440 47048 35492 47054
rect 35440 46990 35492 46996
rect 35268 44662 35388 44690
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 35072 43852 35124 43858
rect 35072 43794 35124 43800
rect 35084 43761 35112 43794
rect 35070 43752 35126 43761
rect 35070 43687 35126 43696
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34978 43344 35034 43353
rect 34978 43279 35034 43288
rect 34992 43246 35020 43279
rect 34980 43240 35032 43246
rect 34980 43182 35032 43188
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34808 42248 34928 42276
rect 34796 42152 34848 42158
rect 34796 42094 34848 42100
rect 34808 41993 34836 42094
rect 34794 41984 34850 41993
rect 34794 41919 34850 41928
rect 34796 41676 34848 41682
rect 34796 41618 34848 41624
rect 34808 41585 34836 41618
rect 34900 41614 34928 42248
rect 34888 41608 34940 41614
rect 34794 41576 34850 41585
rect 34888 41550 34940 41556
rect 35268 41546 35296 44662
rect 35346 44568 35402 44577
rect 35346 44503 35402 44512
rect 35360 44334 35388 44503
rect 35348 44328 35400 44334
rect 35348 44270 35400 44276
rect 35346 44024 35402 44033
rect 35346 43959 35402 43968
rect 35360 43926 35388 43959
rect 35348 43920 35400 43926
rect 35348 43862 35400 43868
rect 35452 43330 35480 46990
rect 35360 43302 35480 43330
rect 35360 42906 35388 43302
rect 35440 43240 35492 43246
rect 35440 43182 35492 43188
rect 35348 42900 35400 42906
rect 35348 42842 35400 42848
rect 35348 42764 35400 42770
rect 35348 42706 35400 42712
rect 35360 42401 35388 42706
rect 35346 42392 35402 42401
rect 35346 42327 35402 42336
rect 35348 41608 35400 41614
rect 35348 41550 35400 41556
rect 34794 41511 34850 41520
rect 35256 41540 35308 41546
rect 35256 41482 35308 41488
rect 34796 41472 34848 41478
rect 34796 41414 34848 41420
rect 34808 41154 34836 41414
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34808 41126 34928 41154
rect 34796 40996 34848 41002
rect 34796 40938 34848 40944
rect 34808 38978 34836 40938
rect 34900 40526 34928 41126
rect 35360 41120 35388 41550
rect 35268 41092 35388 41120
rect 35162 40760 35218 40769
rect 35162 40695 35218 40704
rect 35176 40594 35204 40695
rect 35164 40588 35216 40594
rect 35164 40530 35216 40536
rect 34888 40520 34940 40526
rect 34888 40462 34940 40468
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34888 39840 34940 39846
rect 34888 39782 34940 39788
rect 34900 39642 34928 39782
rect 34888 39636 34940 39642
rect 34888 39578 34940 39584
rect 35268 39438 35296 41092
rect 35348 40996 35400 41002
rect 35348 40938 35400 40944
rect 35256 39432 35308 39438
rect 35256 39374 35308 39380
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 35256 39024 35308 39030
rect 34978 38992 35034 39001
rect 34808 38950 34928 38978
rect 34796 38888 34848 38894
rect 34796 38830 34848 38836
rect 34808 38593 34836 38830
rect 34794 38584 34850 38593
rect 34794 38519 34850 38528
rect 34900 38434 34928 38950
rect 35256 38966 35308 38972
rect 34978 38927 35034 38936
rect 34808 38406 34928 38434
rect 34808 36378 34836 38406
rect 34992 38282 35020 38927
rect 35268 38826 35296 38966
rect 35256 38820 35308 38826
rect 35256 38762 35308 38768
rect 35360 38570 35388 40938
rect 35452 40934 35480 43182
rect 35544 41614 35572 47382
rect 35636 42634 35664 49098
rect 35728 46170 35756 49302
rect 35808 49292 35860 49298
rect 35808 49234 35860 49240
rect 35820 48278 35848 49234
rect 35808 48272 35860 48278
rect 35808 48214 35860 48220
rect 35912 47802 35940 50934
rect 35900 47796 35952 47802
rect 35900 47738 35952 47744
rect 35898 47696 35954 47705
rect 35898 47631 35954 47640
rect 35808 47592 35860 47598
rect 35806 47560 35808 47569
rect 35860 47560 35862 47569
rect 35806 47495 35862 47504
rect 35806 47152 35862 47161
rect 35806 47087 35808 47096
rect 35860 47087 35862 47096
rect 35808 47058 35860 47064
rect 35716 46164 35768 46170
rect 35716 46106 35768 46112
rect 35716 46028 35768 46034
rect 35716 45970 35768 45976
rect 35808 46028 35860 46034
rect 35808 45970 35860 45976
rect 35728 45937 35756 45970
rect 35714 45928 35770 45937
rect 35714 45863 35770 45872
rect 35714 45792 35770 45801
rect 35714 45727 35770 45736
rect 35728 45558 35756 45727
rect 35716 45552 35768 45558
rect 35820 45529 35848 45970
rect 35716 45494 35768 45500
rect 35806 45520 35862 45529
rect 35806 45455 35862 45464
rect 35808 45416 35860 45422
rect 35806 45384 35808 45393
rect 35860 45384 35862 45393
rect 35806 45319 35862 45328
rect 35714 45248 35770 45257
rect 35714 45183 35770 45192
rect 35728 44878 35756 45183
rect 35808 44940 35860 44946
rect 35808 44882 35860 44888
rect 35716 44872 35768 44878
rect 35716 44814 35768 44820
rect 35820 44713 35848 44882
rect 35806 44704 35862 44713
rect 35806 44639 35862 44648
rect 35912 44305 35940 47631
rect 36004 47598 36032 51046
rect 35992 47592 36044 47598
rect 35992 47534 36044 47540
rect 35992 47456 36044 47462
rect 35992 47398 36044 47404
rect 36004 46714 36032 47398
rect 35992 46708 36044 46714
rect 35992 46650 36044 46656
rect 36004 44742 36032 46650
rect 36096 45898 36124 75754
rect 36188 75750 36216 80026
rect 36372 79218 36400 83846
rect 36360 79212 36412 79218
rect 36360 79154 36412 79160
rect 36176 75744 36228 75750
rect 36176 75686 36228 75692
rect 36360 75200 36412 75206
rect 36360 75142 36412 75148
rect 36372 60734 36400 75142
rect 36464 63578 36492 110706
rect 36544 106412 36596 106418
rect 36544 106354 36596 106360
rect 36556 102202 36584 106354
rect 36544 102196 36596 102202
rect 36544 102138 36596 102144
rect 36648 101454 36676 115602
rect 36740 115054 36768 119200
rect 36818 117464 36874 117473
rect 36818 117399 36874 117408
rect 36728 115048 36780 115054
rect 36728 114990 36780 114996
rect 36726 114880 36782 114889
rect 36726 114815 36782 114824
rect 36740 114510 36768 114815
rect 36728 114504 36780 114510
rect 36728 114446 36780 114452
rect 36832 114102 36860 117399
rect 36924 115258 36952 119200
rect 37002 118416 37058 118425
rect 37002 118351 37058 118360
rect 36912 115252 36964 115258
rect 36912 115194 36964 115200
rect 36912 114980 36964 114986
rect 36912 114922 36964 114928
rect 36820 114096 36872 114102
rect 36820 114038 36872 114044
rect 36820 112396 36872 112402
rect 36820 112338 36872 112344
rect 36636 101448 36688 101454
rect 36636 101390 36688 101396
rect 36544 101312 36596 101318
rect 36544 101254 36596 101260
rect 36556 84114 36584 101254
rect 36728 100768 36780 100774
rect 36728 100710 36780 100716
rect 36636 98592 36688 98598
rect 36636 98534 36688 98540
rect 36648 89486 36676 98534
rect 36636 89480 36688 89486
rect 36636 89422 36688 89428
rect 36636 89344 36688 89350
rect 36636 89286 36688 89292
rect 36648 85134 36676 89286
rect 36636 85128 36688 85134
rect 36636 85070 36688 85076
rect 36740 84590 36768 100710
rect 36832 98122 36860 112338
rect 36924 110022 36952 114922
rect 37016 113558 37044 118351
rect 37108 117230 37136 119200
rect 37096 117224 37148 117230
rect 37096 117166 37148 117172
rect 37094 117056 37150 117065
rect 37094 116991 37150 117000
rect 37108 115258 37136 116991
rect 37186 115832 37242 115841
rect 37186 115767 37242 115776
rect 37096 115252 37148 115258
rect 37096 115194 37148 115200
rect 37096 114572 37148 114578
rect 37096 114514 37148 114520
rect 37108 114481 37136 114514
rect 37094 114472 37150 114481
rect 37094 114407 37150 114416
rect 37200 114170 37228 115767
rect 37384 114442 37412 119200
rect 37568 115122 37596 119200
rect 37752 117230 37780 119200
rect 37936 117314 37964 119200
rect 37936 117286 38056 117314
rect 37740 117224 37792 117230
rect 37740 117166 37792 117172
rect 37924 117156 37976 117162
rect 37924 117098 37976 117104
rect 37646 116648 37702 116657
rect 37646 116583 37702 116592
rect 37660 116142 37688 116583
rect 37832 116204 37884 116210
rect 37832 116146 37884 116152
rect 37648 116136 37700 116142
rect 37844 116113 37872 116146
rect 37648 116078 37700 116084
rect 37830 116104 37886 116113
rect 37830 116039 37886 116048
rect 37646 115424 37702 115433
rect 37646 115359 37702 115368
rect 37556 115116 37608 115122
rect 37556 115058 37608 115064
rect 37660 115054 37688 115359
rect 37648 115048 37700 115054
rect 37648 114990 37700 114996
rect 37372 114436 37424 114442
rect 37372 114378 37424 114384
rect 37280 114368 37332 114374
rect 37280 114310 37332 114316
rect 37188 114164 37240 114170
rect 37188 114106 37240 114112
rect 37004 113552 37056 113558
rect 37004 113494 37056 113500
rect 37186 110256 37242 110265
rect 37186 110191 37188 110200
rect 37240 110191 37242 110200
rect 37188 110162 37240 110168
rect 36912 110016 36964 110022
rect 36912 109958 36964 109964
rect 37186 109712 37242 109721
rect 37186 109647 37242 109656
rect 37200 109614 37228 109647
rect 37188 109608 37240 109614
rect 37188 109550 37240 109556
rect 37188 109132 37240 109138
rect 37188 109074 37240 109080
rect 37200 108905 37228 109074
rect 37292 109034 37320 114310
rect 37370 114064 37426 114073
rect 37370 113999 37372 114008
rect 37424 113999 37426 114008
rect 37372 113970 37424 113976
rect 37464 113892 37516 113898
rect 37464 113834 37516 113840
rect 37372 113348 37424 113354
rect 37372 113290 37424 113296
rect 37384 113257 37412 113290
rect 37370 113248 37426 113257
rect 37370 113183 37426 113192
rect 37370 112840 37426 112849
rect 37370 112775 37372 112784
rect 37424 112775 37426 112784
rect 37372 112746 37424 112752
rect 37372 111172 37424 111178
rect 37372 111114 37424 111120
rect 37384 111081 37412 111114
rect 37476 111110 37504 113834
rect 37646 111888 37702 111897
rect 37646 111823 37702 111832
rect 37660 111790 37688 111823
rect 37648 111784 37700 111790
rect 37648 111726 37700 111732
rect 37464 111104 37516 111110
rect 37370 111072 37426 111081
rect 37464 111046 37516 111052
rect 37370 111007 37426 111016
rect 37464 110696 37516 110702
rect 37462 110664 37464 110673
rect 37516 110664 37518 110673
rect 37462 110599 37518 110608
rect 37832 110628 37884 110634
rect 37832 110570 37884 110576
rect 37844 109818 37872 110570
rect 37832 109812 37884 109818
rect 37832 109754 37884 109760
rect 37936 109698 37964 117098
rect 38028 115190 38056 117286
rect 38212 116278 38240 119200
rect 38200 116272 38252 116278
rect 38200 116214 38252 116220
rect 38016 115184 38068 115190
rect 38016 115126 38068 115132
rect 38292 114980 38344 114986
rect 38292 114922 38344 114928
rect 38108 112804 38160 112810
rect 38108 112746 38160 112752
rect 38120 112305 38148 112746
rect 38106 112296 38162 112305
rect 38106 112231 38162 112240
rect 38200 110084 38252 110090
rect 38200 110026 38252 110032
rect 37844 109670 37964 109698
rect 37292 109006 37412 109034
rect 37186 108896 37242 108905
rect 37186 108831 37242 108840
rect 37186 108080 37242 108089
rect 37186 108015 37188 108024
rect 37240 108015 37242 108024
rect 37188 107986 37240 107992
rect 37384 107642 37412 109006
rect 37372 107636 37424 107642
rect 37372 107578 37424 107584
rect 37186 107536 37242 107545
rect 37186 107471 37242 107480
rect 37200 107438 37228 107471
rect 37188 107432 37240 107438
rect 37188 107374 37240 107380
rect 37556 107364 37608 107370
rect 37556 107306 37608 107312
rect 36912 107296 36964 107302
rect 36912 107238 36964 107244
rect 36924 103562 36952 107238
rect 37188 106956 37240 106962
rect 37188 106898 37240 106904
rect 37200 106729 37228 106898
rect 37186 106720 37242 106729
rect 37186 106655 37242 106664
rect 37280 106344 37332 106350
rect 37278 106312 37280 106321
rect 37332 106312 37334 106321
rect 37278 106247 37334 106256
rect 37186 105904 37242 105913
rect 37186 105839 37188 105848
rect 37240 105839 37242 105848
rect 37188 105810 37240 105816
rect 37186 105496 37242 105505
rect 37186 105431 37242 105440
rect 37200 105262 37228 105431
rect 37188 105256 37240 105262
rect 37188 105198 37240 105204
rect 37188 104780 37240 104786
rect 37188 104722 37240 104728
rect 37004 104576 37056 104582
rect 37200 104553 37228 104722
rect 37004 104518 37056 104524
rect 37186 104544 37242 104553
rect 36912 103556 36964 103562
rect 36912 103498 36964 103504
rect 36912 102196 36964 102202
rect 36912 102138 36964 102144
rect 36820 98116 36872 98122
rect 36820 98058 36872 98064
rect 36820 96484 36872 96490
rect 36820 96426 36872 96432
rect 36728 84584 36780 84590
rect 36728 84526 36780 84532
rect 36544 84108 36596 84114
rect 36544 84050 36596 84056
rect 36728 80096 36780 80102
rect 36728 80038 36780 80044
rect 36452 63572 36504 63578
rect 36452 63514 36504 63520
rect 36740 60734 36768 80038
rect 36832 79762 36860 96426
rect 36924 86954 36952 102138
rect 37016 87514 37044 104518
rect 37186 104479 37242 104488
rect 37186 104136 37242 104145
rect 37186 104071 37188 104080
rect 37240 104071 37242 104080
rect 37372 104100 37424 104106
rect 37188 104042 37240 104048
rect 37372 104042 37424 104048
rect 37188 103692 37240 103698
rect 37188 103634 37240 103640
rect 37200 103329 37228 103634
rect 37186 103320 37242 103329
rect 37186 103255 37242 103264
rect 37280 103080 37332 103086
rect 37280 103022 37332 103028
rect 37292 102921 37320 103022
rect 37278 102912 37334 102921
rect 37278 102847 37334 102856
rect 37188 102604 37240 102610
rect 37188 102546 37240 102552
rect 37200 102377 37228 102546
rect 37280 102400 37332 102406
rect 37186 102368 37242 102377
rect 37280 102342 37332 102348
rect 37186 102303 37242 102312
rect 37186 101552 37242 101561
rect 37186 101487 37188 101496
rect 37240 101487 37242 101496
rect 37188 101458 37240 101464
rect 37188 100836 37240 100842
rect 37188 100778 37240 100784
rect 37200 100745 37228 100778
rect 37186 100736 37242 100745
rect 37186 100671 37242 100680
rect 37188 100428 37240 100434
rect 37188 100370 37240 100376
rect 37200 100337 37228 100370
rect 37186 100328 37242 100337
rect 37186 100263 37242 100272
rect 37292 99498 37320 102342
rect 37384 100978 37412 104042
rect 37372 100972 37424 100978
rect 37372 100914 37424 100920
rect 37108 99470 37320 99498
rect 37108 94738 37136 99470
rect 37186 99376 37242 99385
rect 37186 99311 37188 99320
rect 37240 99311 37242 99320
rect 37188 99282 37240 99288
rect 37186 98968 37242 98977
rect 37186 98903 37242 98912
rect 37200 98734 37228 98903
rect 37188 98728 37240 98734
rect 37188 98670 37240 98676
rect 37188 98252 37240 98258
rect 37188 98194 37240 98200
rect 37200 98161 37228 98194
rect 37186 98152 37242 98161
rect 37186 98087 37242 98096
rect 37186 97200 37242 97209
rect 37186 97135 37188 97144
rect 37240 97135 37242 97144
rect 37188 97106 37240 97112
rect 37188 96552 37240 96558
rect 37188 96494 37240 96500
rect 37200 96393 37228 96494
rect 37186 96384 37242 96393
rect 37186 96319 37242 96328
rect 37188 96076 37240 96082
rect 37188 96018 37240 96024
rect 37200 95985 37228 96018
rect 37186 95976 37242 95985
rect 37186 95911 37242 95920
rect 37278 95568 37334 95577
rect 37278 95503 37334 95512
rect 37292 95470 37320 95503
rect 37280 95464 37332 95470
rect 37280 95406 37332 95412
rect 37186 95024 37242 95033
rect 37186 94959 37188 94968
rect 37240 94959 37242 94968
rect 37188 94930 37240 94936
rect 37108 94710 37228 94738
rect 37200 93106 37228 94710
rect 37568 94450 37596 107306
rect 37844 107030 37872 109670
rect 37924 109540 37976 109546
rect 37924 109482 37976 109488
rect 37936 109313 37964 109482
rect 37922 109304 37978 109313
rect 37922 109239 37978 109248
rect 37922 108488 37978 108497
rect 37922 108423 37924 108432
rect 37976 108423 37978 108432
rect 37924 108394 37976 108400
rect 37924 107364 37976 107370
rect 37924 107306 37976 107312
rect 37936 107137 37964 107306
rect 37922 107128 37978 107137
rect 37922 107063 37978 107072
rect 37832 107024 37884 107030
rect 37832 106966 37884 106972
rect 37924 105188 37976 105194
rect 37924 105130 37976 105136
rect 37936 104961 37964 105130
rect 38016 105120 38068 105126
rect 38016 105062 38068 105068
rect 37922 104952 37978 104961
rect 37922 104887 37978 104896
rect 38028 104174 38056 105062
rect 38016 104168 38068 104174
rect 38016 104110 38068 104116
rect 37924 104100 37976 104106
rect 37924 104042 37976 104048
rect 37936 103737 37964 104042
rect 38016 104032 38068 104038
rect 38016 103974 38068 103980
rect 37922 103728 37978 103737
rect 37922 103663 37978 103672
rect 38028 102202 38056 103974
rect 38016 102196 38068 102202
rect 38016 102138 38068 102144
rect 37922 101960 37978 101969
rect 37922 101895 37924 101904
rect 37976 101895 37978 101904
rect 37924 101866 37976 101872
rect 37922 101144 37978 101153
rect 37922 101079 37978 101088
rect 37936 100910 37964 101079
rect 37924 100904 37976 100910
rect 37924 100846 37976 100852
rect 37648 100836 37700 100842
rect 37648 100778 37700 100784
rect 37660 94790 37688 100778
rect 37922 99784 37978 99793
rect 37922 99719 37924 99728
rect 37976 99719 37978 99728
rect 37924 99690 37976 99696
rect 37832 99680 37884 99686
rect 37832 99622 37884 99628
rect 37844 99374 37872 99622
rect 37844 99346 38148 99374
rect 37740 98660 37792 98666
rect 37740 98602 37792 98608
rect 37924 98660 37976 98666
rect 37924 98602 37976 98608
rect 37648 94784 37700 94790
rect 37648 94726 37700 94732
rect 37556 94444 37608 94450
rect 37556 94386 37608 94392
rect 37280 94376 37332 94382
rect 37280 94318 37332 94324
rect 37292 94217 37320 94318
rect 37464 94240 37516 94246
rect 37278 94208 37334 94217
rect 37464 94182 37516 94188
rect 37278 94143 37334 94152
rect 37278 93392 37334 93401
rect 37278 93327 37334 93336
rect 37292 93294 37320 93327
rect 37280 93288 37332 93294
rect 37280 93230 37332 93236
rect 37200 93078 37320 93106
rect 37186 92984 37242 92993
rect 37186 92919 37242 92928
rect 37200 92818 37228 92919
rect 37188 92812 37240 92818
rect 37188 92754 37240 92760
rect 37292 92698 37320 93078
rect 37200 92670 37320 92698
rect 37200 90930 37228 92670
rect 37372 92608 37424 92614
rect 37372 92550 37424 92556
rect 37280 92200 37332 92206
rect 37280 92142 37332 92148
rect 37292 92041 37320 92142
rect 37278 92032 37334 92041
rect 37278 91967 37334 91976
rect 37278 91216 37334 91225
rect 37278 91151 37334 91160
rect 37292 91118 37320 91151
rect 37280 91112 37332 91118
rect 37280 91054 37332 91060
rect 37200 90902 37320 90930
rect 37186 90808 37242 90817
rect 37186 90743 37242 90752
rect 37200 90642 37228 90743
rect 37188 90636 37240 90642
rect 37188 90578 37240 90584
rect 37292 90522 37320 90902
rect 37200 90494 37320 90522
rect 37200 89350 37228 90494
rect 37280 90024 37332 90030
rect 37280 89966 37332 89972
rect 37292 89865 37320 89966
rect 37278 89856 37334 89865
rect 37278 89791 37334 89800
rect 37188 89344 37240 89350
rect 37188 89286 37240 89292
rect 37278 89040 37334 89049
rect 37278 88975 37334 88984
rect 37292 88942 37320 88975
rect 37280 88936 37332 88942
rect 37280 88878 37332 88884
rect 37384 88874 37412 92550
rect 37476 91118 37504 94182
rect 37648 93152 37700 93158
rect 37648 93094 37700 93100
rect 37556 91248 37608 91254
rect 37556 91190 37608 91196
rect 37464 91112 37516 91118
rect 37464 91054 37516 91060
rect 37464 89888 37516 89894
rect 37464 89830 37516 89836
rect 37372 88868 37424 88874
rect 37372 88810 37424 88816
rect 37186 88632 37242 88641
rect 37186 88567 37242 88576
rect 37200 88466 37228 88567
rect 37188 88460 37240 88466
rect 37188 88402 37240 88408
rect 37280 87848 37332 87854
rect 37278 87816 37280 87825
rect 37332 87816 37334 87825
rect 37278 87751 37334 87760
rect 37004 87508 37056 87514
rect 37004 87450 37056 87456
rect 37476 86970 37504 89830
rect 37568 87446 37596 91190
rect 37660 89078 37688 93094
rect 37648 89072 37700 89078
rect 37648 89014 37700 89020
rect 37556 87440 37608 87446
rect 37556 87382 37608 87388
rect 37464 86964 37516 86970
rect 36924 86926 37136 86954
rect 37108 86222 37136 86926
rect 37464 86906 37516 86912
rect 37278 86864 37334 86873
rect 37278 86799 37334 86808
rect 37292 86766 37320 86799
rect 37280 86760 37332 86766
rect 37280 86702 37332 86708
rect 37556 86624 37608 86630
rect 37556 86566 37608 86572
rect 37648 86624 37700 86630
rect 37648 86566 37700 86572
rect 37186 86456 37242 86465
rect 37186 86391 37242 86400
rect 37200 86290 37228 86391
rect 37188 86284 37240 86290
rect 37188 86226 37240 86232
rect 37096 86216 37148 86222
rect 37096 86158 37148 86164
rect 37372 86080 37424 86086
rect 37372 86022 37424 86028
rect 36912 85808 36964 85814
rect 36912 85750 36964 85756
rect 36924 80170 36952 85750
rect 37280 85672 37332 85678
rect 37278 85640 37280 85649
rect 37332 85640 37334 85649
rect 37278 85575 37334 85584
rect 37278 84688 37334 84697
rect 37278 84623 37334 84632
rect 37292 84590 37320 84623
rect 37280 84584 37332 84590
rect 37280 84526 37332 84532
rect 37186 84280 37242 84289
rect 37186 84215 37242 84224
rect 37200 84114 37228 84215
rect 37188 84108 37240 84114
rect 37188 84050 37240 84056
rect 37280 83496 37332 83502
rect 37278 83464 37280 83473
rect 37332 83464 37334 83473
rect 37278 83399 37334 83408
rect 37384 82550 37412 86022
rect 37464 83360 37516 83366
rect 37464 83302 37516 83308
rect 37372 82544 37424 82550
rect 37278 82512 37334 82521
rect 37372 82486 37424 82492
rect 37278 82447 37334 82456
rect 37292 82414 37320 82447
rect 37280 82408 37332 82414
rect 37280 82350 37332 82356
rect 37280 82272 37332 82278
rect 37280 82214 37332 82220
rect 37186 82104 37242 82113
rect 37186 82039 37242 82048
rect 37200 81938 37228 82039
rect 37188 81932 37240 81938
rect 37188 81874 37240 81880
rect 37292 81410 37320 82214
rect 37016 81382 37320 81410
rect 36912 80164 36964 80170
rect 36912 80106 36964 80112
rect 36820 79756 36872 79762
rect 36820 79698 36872 79704
rect 36820 77376 36872 77382
rect 36820 77318 36872 77324
rect 36188 60706 36400 60734
rect 36648 60706 36768 60734
rect 36084 45892 36136 45898
rect 36084 45834 36136 45840
rect 36082 45656 36138 45665
rect 36082 45591 36084 45600
rect 36136 45591 36138 45600
rect 36084 45562 36136 45568
rect 36082 45112 36138 45121
rect 36082 45047 36138 45056
rect 36096 45014 36124 45047
rect 36084 45008 36136 45014
rect 36084 44950 36136 44956
rect 36084 44872 36136 44878
rect 36084 44814 36136 44820
rect 35992 44736 36044 44742
rect 35992 44678 36044 44684
rect 35898 44296 35954 44305
rect 35716 44260 35768 44266
rect 35898 44231 35954 44240
rect 35992 44260 36044 44266
rect 35716 44202 35768 44208
rect 35992 44202 36044 44208
rect 35728 43738 35756 44202
rect 35900 44192 35952 44198
rect 35806 44160 35862 44169
rect 35900 44134 35952 44140
rect 35806 44095 35862 44104
rect 35820 43858 35848 44095
rect 35912 43994 35940 44134
rect 35900 43988 35952 43994
rect 35900 43930 35952 43936
rect 35808 43852 35860 43858
rect 35808 43794 35860 43800
rect 35728 43710 35848 43738
rect 35714 42936 35770 42945
rect 35714 42871 35770 42880
rect 35728 42770 35756 42871
rect 35716 42764 35768 42770
rect 35716 42706 35768 42712
rect 35624 42628 35676 42634
rect 35624 42570 35676 42576
rect 35716 42628 35768 42634
rect 35716 42570 35768 42576
rect 35532 41608 35584 41614
rect 35532 41550 35584 41556
rect 35532 41472 35584 41478
rect 35532 41414 35584 41420
rect 35728 41414 35756 42570
rect 35820 41682 35848 43710
rect 35912 41818 35940 43930
rect 35900 41812 35952 41818
rect 35900 41754 35952 41760
rect 35808 41676 35860 41682
rect 35808 41618 35860 41624
rect 35900 41676 35952 41682
rect 35900 41618 35952 41624
rect 35808 41540 35860 41546
rect 35808 41482 35860 41488
rect 35440 40928 35492 40934
rect 35440 40870 35492 40876
rect 35440 40520 35492 40526
rect 35440 40462 35492 40468
rect 35268 38542 35388 38570
rect 34980 38276 35032 38282
rect 34980 38218 35032 38224
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 35164 37664 35216 37670
rect 35164 37606 35216 37612
rect 35176 37466 35204 37606
rect 35164 37460 35216 37466
rect 35164 37402 35216 37408
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34796 36372 34848 36378
rect 34796 36314 34848 36320
rect 34796 36236 34848 36242
rect 34796 36178 34848 36184
rect 34808 36145 34836 36178
rect 34794 36136 34850 36145
rect 34794 36071 34850 36080
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35268 35834 35296 38542
rect 35348 38412 35400 38418
rect 35348 38354 35400 38360
rect 35360 38185 35388 38354
rect 35346 38176 35402 38185
rect 35346 38111 35402 38120
rect 35348 37664 35400 37670
rect 35348 37606 35400 37612
rect 35360 36122 35388 37606
rect 35452 36530 35480 40462
rect 35544 39642 35572 41414
rect 35636 41386 35756 41414
rect 35532 39636 35584 39642
rect 35532 39578 35584 39584
rect 35532 39500 35584 39506
rect 35532 39442 35584 39448
rect 35544 39098 35572 39442
rect 35532 39092 35584 39098
rect 35532 39034 35584 39040
rect 35530 38992 35586 39001
rect 35530 38927 35586 38936
rect 35544 38826 35572 38927
rect 35532 38820 35584 38826
rect 35532 38762 35584 38768
rect 35636 38554 35664 41386
rect 35820 40712 35848 41482
rect 35728 40684 35848 40712
rect 35728 40050 35756 40684
rect 35808 40588 35860 40594
rect 35808 40530 35860 40536
rect 35820 40361 35848 40530
rect 35806 40352 35862 40361
rect 35806 40287 35862 40296
rect 35716 40044 35768 40050
rect 35716 39986 35768 39992
rect 35808 39908 35860 39914
rect 35808 39850 35860 39856
rect 35714 38992 35770 39001
rect 35714 38927 35770 38936
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 35728 38418 35756 38927
rect 35716 38412 35768 38418
rect 35716 38354 35768 38360
rect 35532 38344 35584 38350
rect 35532 38286 35584 38292
rect 35544 37670 35572 38286
rect 35716 37936 35768 37942
rect 35716 37878 35768 37884
rect 35532 37664 35584 37670
rect 35532 37606 35584 37612
rect 35532 37324 35584 37330
rect 35532 37266 35584 37272
rect 35544 37233 35572 37266
rect 35624 37256 35676 37262
rect 35530 37224 35586 37233
rect 35624 37198 35676 37204
rect 35530 37159 35586 37168
rect 35636 36650 35664 37198
rect 35624 36644 35676 36650
rect 35624 36586 35676 36592
rect 35728 36530 35756 37878
rect 35452 36502 35572 36530
rect 35438 36408 35494 36417
rect 35438 36343 35494 36352
rect 35452 36242 35480 36343
rect 35440 36236 35492 36242
rect 35440 36178 35492 36184
rect 35360 36094 35480 36122
rect 35256 35828 35308 35834
rect 35256 35770 35308 35776
rect 34796 35624 34848 35630
rect 34794 35592 34796 35601
rect 34848 35592 34850 35601
rect 34794 35527 34850 35536
rect 35348 35556 35400 35562
rect 35348 35498 35400 35504
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35256 32836 35308 32842
rect 35256 32778 35308 32784
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34796 31748 34848 31754
rect 34796 31690 34848 31696
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 34624 30110 34744 30138
rect 34612 29572 34664 29578
rect 34612 29514 34664 29520
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34624 28994 34652 29514
rect 34532 28966 34652 28994
rect 34532 22710 34560 28966
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34624 25226 34652 26930
rect 34612 25220 34664 25226
rect 34612 25162 34664 25168
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34428 18080 34480 18086
rect 34428 18022 34480 18028
rect 34336 17264 34388 17270
rect 34336 17206 34388 17212
rect 34520 14272 34572 14278
rect 34520 14214 34572 14220
rect 34532 4758 34560 14214
rect 34624 5234 34652 22442
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34612 5092 34664 5098
rect 34612 5034 34664 5040
rect 34520 4752 34572 4758
rect 34520 4694 34572 4700
rect 34336 4208 34388 4214
rect 34624 4162 34652 5034
rect 34336 4150 34388 4156
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 34348 3670 34376 4150
rect 34440 4134 34652 4162
rect 34336 3664 34388 3670
rect 34336 3606 34388 3612
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 34244 3596 34296 3602
rect 34244 3538 34296 3544
rect 33876 3188 33928 3194
rect 33876 3130 33928 3136
rect 33784 2644 33836 2650
rect 33784 2586 33836 2592
rect 33980 800 34008 3538
rect 34256 800 34284 3538
rect 34440 3398 34468 4134
rect 34520 4072 34572 4078
rect 34520 4014 34572 4020
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34428 2984 34480 2990
rect 34428 2926 34480 2932
rect 34440 2825 34468 2926
rect 34426 2816 34482 2825
rect 34426 2751 34482 2760
rect 34532 800 34560 4014
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34624 3670 34652 3878
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34716 2582 34744 30110
rect 34808 3738 34836 31690
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35268 30870 35296 32778
rect 35256 30864 35308 30870
rect 35256 30806 35308 30812
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34980 30116 35032 30122
rect 34980 30058 35032 30064
rect 34992 29578 35020 30058
rect 34980 29572 35032 29578
rect 34980 29514 35032 29520
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 35072 29232 35124 29238
rect 35072 29174 35124 29180
rect 35084 28694 35112 29174
rect 35164 29164 35216 29170
rect 35164 29106 35216 29112
rect 35072 28688 35124 28694
rect 35072 28630 35124 28636
rect 35176 28490 35204 29106
rect 35164 28484 35216 28490
rect 35164 28426 35216 28432
rect 35256 28416 35308 28422
rect 35256 28358 35308 28364
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35268 25294 35296 28358
rect 35360 26858 35388 35498
rect 35452 33538 35480 36094
rect 35544 35737 35572 36502
rect 35636 36502 35756 36530
rect 35530 35728 35586 35737
rect 35530 35663 35586 35672
rect 35532 35624 35584 35630
rect 35532 35566 35584 35572
rect 35544 34950 35572 35566
rect 35636 35154 35664 36502
rect 35820 36394 35848 39850
rect 35912 39506 35940 41618
rect 35900 39500 35952 39506
rect 35900 39442 35952 39448
rect 35912 36922 35940 39442
rect 36004 39370 36032 44202
rect 36096 40458 36124 44814
rect 36188 42158 36216 60706
rect 36544 59628 36596 59634
rect 36544 59570 36596 59576
rect 36268 59424 36320 59430
rect 36268 59366 36320 59372
rect 36280 56284 36308 59366
rect 36452 59084 36504 59090
rect 36452 59026 36504 59032
rect 36360 59016 36412 59022
rect 36360 58958 36412 58964
rect 36372 58562 36400 58958
rect 36464 58857 36492 59026
rect 36450 58848 36506 58857
rect 36450 58783 36506 58792
rect 36372 58534 36492 58562
rect 36464 58478 36492 58534
rect 36360 58472 36412 58478
rect 36360 58414 36412 58420
rect 36452 58472 36504 58478
rect 36452 58414 36504 58420
rect 36372 56794 36400 58414
rect 36450 58032 36506 58041
rect 36450 57967 36452 57976
rect 36504 57967 36506 57976
rect 36452 57938 36504 57944
rect 36556 57882 36584 59570
rect 36464 57854 36584 57882
rect 36464 57202 36492 57854
rect 36544 57792 36596 57798
rect 36544 57734 36596 57740
rect 36556 57594 36584 57734
rect 36544 57588 36596 57594
rect 36544 57530 36596 57536
rect 36464 57174 36584 57202
rect 36450 57080 36506 57089
rect 36450 57015 36506 57024
rect 36464 56982 36492 57015
rect 36452 56976 36504 56982
rect 36452 56918 36504 56924
rect 36372 56766 36492 56794
rect 36360 56296 36412 56302
rect 36280 56256 36360 56284
rect 36280 55962 36308 56256
rect 36360 56238 36412 56244
rect 36268 55956 36320 55962
rect 36320 55916 36400 55944
rect 36268 55898 36320 55904
rect 36268 55820 36320 55826
rect 36268 55762 36320 55768
rect 36280 54330 36308 55762
rect 36372 55350 36400 55916
rect 36464 55418 36492 56766
rect 36556 56438 36584 57174
rect 36544 56432 36596 56438
rect 36544 56374 36596 56380
rect 36544 56228 36596 56234
rect 36544 56170 36596 56176
rect 36556 55826 36584 56170
rect 36544 55820 36596 55826
rect 36544 55762 36596 55768
rect 36452 55412 36504 55418
rect 36452 55354 36504 55360
rect 36360 55344 36412 55350
rect 36360 55286 36412 55292
rect 36452 55276 36504 55282
rect 36452 55218 36504 55224
rect 36360 55208 36412 55214
rect 36360 55150 36412 55156
rect 36268 54324 36320 54330
rect 36268 54266 36320 54272
rect 36268 54052 36320 54058
rect 36268 53994 36320 54000
rect 36280 51338 36308 53994
rect 36372 52698 36400 55150
rect 36464 53786 36492 55218
rect 36556 55146 36584 55762
rect 36544 55140 36596 55146
rect 36544 55082 36596 55088
rect 36556 54738 36584 55082
rect 36544 54732 36596 54738
rect 36544 54674 36596 54680
rect 36452 53780 36504 53786
rect 36452 53722 36504 53728
rect 36360 52692 36412 52698
rect 36360 52634 36412 52640
rect 36556 52578 36584 54674
rect 36648 53038 36676 60706
rect 36728 59764 36780 59770
rect 36728 59706 36780 59712
rect 36740 59498 36768 59706
rect 36832 59634 36860 77318
rect 36820 59628 36872 59634
rect 36820 59570 36872 59576
rect 36912 59560 36964 59566
rect 36912 59502 36964 59508
rect 36728 59492 36780 59498
rect 36728 59434 36780 59440
rect 36740 58546 36768 59434
rect 36820 59424 36872 59430
rect 36820 59366 36872 59372
rect 36728 58540 36780 58546
rect 36728 58482 36780 58488
rect 36728 57996 36780 58002
rect 36728 57938 36780 57944
rect 36740 53786 36768 57938
rect 36832 55826 36860 59366
rect 36924 59265 36952 59502
rect 36910 59256 36966 59265
rect 36910 59191 36966 59200
rect 37016 59022 37044 81382
rect 37280 81320 37332 81326
rect 37278 81288 37280 81297
rect 37332 81288 37334 81297
rect 37278 81223 37334 81232
rect 37278 80472 37334 80481
rect 37278 80407 37334 80416
rect 37292 80238 37320 80407
rect 37280 80232 37332 80238
rect 37280 80174 37332 80180
rect 37186 79928 37242 79937
rect 37186 79863 37242 79872
rect 37200 79762 37228 79863
rect 37188 79756 37240 79762
rect 37188 79698 37240 79704
rect 37476 79150 37504 83302
rect 37568 82346 37596 86566
rect 37660 83434 37688 86566
rect 37752 84794 37780 98602
rect 37936 98569 37964 98602
rect 37922 98560 37978 98569
rect 37922 98495 37978 98504
rect 37922 97744 37978 97753
rect 37922 97679 37978 97688
rect 37936 97646 37964 97679
rect 37924 97640 37976 97646
rect 37924 97582 37976 97588
rect 37922 96792 37978 96801
rect 37922 96727 37978 96736
rect 37936 96558 37964 96727
rect 37924 96552 37976 96558
rect 37924 96494 37976 96500
rect 37924 95464 37976 95470
rect 37924 95406 37976 95412
rect 37936 94625 37964 95406
rect 37922 94616 37978 94625
rect 37922 94551 37978 94560
rect 37924 94376 37976 94382
rect 37924 94318 37976 94324
rect 37936 93809 37964 94318
rect 37922 93800 37978 93809
rect 37922 93735 37978 93744
rect 37924 92200 37976 92206
rect 37924 92142 37976 92148
rect 37936 91633 37964 92142
rect 37922 91624 37978 91633
rect 37922 91559 37978 91568
rect 37924 91112 37976 91118
rect 37924 91054 37976 91060
rect 37936 90409 37964 91054
rect 38016 90432 38068 90438
rect 37922 90400 37978 90409
rect 38016 90374 38068 90380
rect 37922 90335 37978 90344
rect 37924 90024 37976 90030
rect 37924 89966 37976 89972
rect 37936 89457 37964 89966
rect 37922 89448 37978 89457
rect 37922 89383 37978 89392
rect 37924 88936 37976 88942
rect 37924 88878 37976 88884
rect 37936 88233 37964 88878
rect 37922 88224 37978 88233
rect 37922 88159 37978 88168
rect 37924 87848 37976 87854
rect 37924 87790 37976 87796
rect 37936 87281 37964 87790
rect 37922 87272 37978 87281
rect 37922 87207 37978 87216
rect 37924 86760 37976 86766
rect 37924 86702 37976 86708
rect 37936 86057 37964 86702
rect 38028 86601 38056 90374
rect 38120 88942 38148 99346
rect 38108 88936 38160 88942
rect 38108 88878 38160 88884
rect 38108 88800 38160 88806
rect 38108 88742 38160 88748
rect 38120 88534 38148 88742
rect 38108 88528 38160 88534
rect 38108 88470 38160 88476
rect 38014 86592 38070 86601
rect 38014 86527 38070 86536
rect 37922 86048 37978 86057
rect 37922 85983 37978 85992
rect 37924 85672 37976 85678
rect 37924 85614 37976 85620
rect 37936 85241 37964 85614
rect 37922 85232 37978 85241
rect 37922 85167 37978 85176
rect 38212 84946 38240 110026
rect 38028 84918 38240 84946
rect 37740 84788 37792 84794
rect 37740 84730 37792 84736
rect 37924 84584 37976 84590
rect 37924 84526 37976 84532
rect 37740 84448 37792 84454
rect 37740 84390 37792 84396
rect 37648 83428 37700 83434
rect 37648 83370 37700 83376
rect 37556 82340 37608 82346
rect 37556 82282 37608 82288
rect 37556 81728 37608 81734
rect 37556 81670 37608 81676
rect 37464 79144 37516 79150
rect 37464 79086 37516 79092
rect 37188 78736 37240 78742
rect 37186 78704 37188 78713
rect 37240 78704 37242 78713
rect 37186 78639 37242 78648
rect 37186 78296 37242 78305
rect 37186 78231 37242 78240
rect 37200 78062 37228 78231
rect 37188 78056 37240 78062
rect 37188 77998 37240 78004
rect 37280 77920 37332 77926
rect 37280 77862 37332 77868
rect 37292 77722 37320 77862
rect 37280 77716 37332 77722
rect 37280 77658 37332 77664
rect 37188 77580 37240 77586
rect 37188 77522 37240 77528
rect 37200 77353 37228 77522
rect 37186 77344 37242 77353
rect 37186 77279 37242 77288
rect 37186 76528 37242 76537
rect 37186 76463 37188 76472
rect 37240 76463 37242 76472
rect 37188 76434 37240 76440
rect 37186 76120 37242 76129
rect 37186 76055 37242 76064
rect 37200 75886 37228 76055
rect 37188 75880 37240 75886
rect 37188 75822 37240 75828
rect 37280 75744 37332 75750
rect 37280 75686 37332 75692
rect 37292 75546 37320 75686
rect 37280 75540 37332 75546
rect 37280 75482 37332 75488
rect 37188 75404 37240 75410
rect 37188 75346 37240 75352
rect 37200 75313 37228 75346
rect 37186 75304 37242 75313
rect 37186 75239 37242 75248
rect 37186 74352 37242 74361
rect 37186 74287 37188 74296
rect 37240 74287 37242 74296
rect 37188 74258 37240 74264
rect 37186 73944 37242 73953
rect 37186 73879 37242 73888
rect 37200 73710 37228 73879
rect 37188 73704 37240 73710
rect 37188 73646 37240 73652
rect 37280 73568 37332 73574
rect 37280 73510 37332 73516
rect 37292 73370 37320 73510
rect 37280 73364 37332 73370
rect 37280 73306 37332 73312
rect 37188 73228 37240 73234
rect 37188 73170 37240 73176
rect 37200 73137 37228 73170
rect 37186 73128 37242 73137
rect 37186 73063 37242 73072
rect 37096 73024 37148 73030
rect 37096 72966 37148 72972
rect 37004 59016 37056 59022
rect 37004 58958 37056 58964
rect 37004 58608 37056 58614
rect 37004 58550 37056 58556
rect 36912 58472 36964 58478
rect 36912 58414 36964 58420
rect 36820 55820 36872 55826
rect 36820 55762 36872 55768
rect 36924 55434 36952 58414
rect 37016 58002 37044 58550
rect 37004 57996 37056 58002
rect 37004 57938 37056 57944
rect 37004 57384 37056 57390
rect 37004 57326 37056 57332
rect 37016 56273 37044 57326
rect 37002 56264 37058 56273
rect 37002 56199 37058 56208
rect 37108 56114 37136 72966
rect 37186 72176 37242 72185
rect 37186 72111 37188 72120
rect 37240 72111 37242 72120
rect 37188 72082 37240 72088
rect 37186 71768 37242 71777
rect 37186 71703 37242 71712
rect 37200 71534 37228 71703
rect 37188 71528 37240 71534
rect 37188 71470 37240 71476
rect 37188 71052 37240 71058
rect 37188 70994 37240 71000
rect 37200 70961 37228 70994
rect 37186 70952 37242 70961
rect 37186 70887 37242 70896
rect 37186 70000 37242 70009
rect 37186 69935 37188 69944
rect 37240 69935 37242 69944
rect 37188 69906 37240 69912
rect 37186 69592 37242 69601
rect 37186 69527 37242 69536
rect 37200 69290 37228 69527
rect 37188 69284 37240 69290
rect 37188 69226 37240 69232
rect 37188 68876 37240 68882
rect 37188 68818 37240 68824
rect 37200 68785 37228 68818
rect 37186 68776 37242 68785
rect 37186 68711 37242 68720
rect 37278 68368 37334 68377
rect 37278 68303 37334 68312
rect 37292 68270 37320 68303
rect 37280 68264 37332 68270
rect 37280 68206 37332 68212
rect 37186 67960 37242 67969
rect 37186 67895 37242 67904
rect 37200 67794 37228 67895
rect 37188 67788 37240 67794
rect 37188 67730 37240 67736
rect 37372 67652 37424 67658
rect 37372 67594 37424 67600
rect 37280 67176 37332 67182
rect 37280 67118 37332 67124
rect 37292 67017 37320 67118
rect 37278 67008 37334 67017
rect 37278 66943 37334 66952
rect 37278 66192 37334 66201
rect 37278 66127 37334 66136
rect 37292 66094 37320 66127
rect 37280 66088 37332 66094
rect 37280 66030 37332 66036
rect 37186 65784 37242 65793
rect 37186 65719 37242 65728
rect 37200 65618 37228 65719
rect 37188 65612 37240 65618
rect 37188 65554 37240 65560
rect 37188 65000 37240 65006
rect 37188 64942 37240 64948
rect 37200 64841 37228 64942
rect 37186 64832 37242 64841
rect 37186 64767 37242 64776
rect 37278 64016 37334 64025
rect 37278 63951 37334 63960
rect 37292 63918 37320 63951
rect 37280 63912 37332 63918
rect 37280 63854 37332 63860
rect 37186 63608 37242 63617
rect 37186 63543 37242 63552
rect 37200 63442 37228 63543
rect 37188 63436 37240 63442
rect 37188 63378 37240 63384
rect 37280 62824 37332 62830
rect 37278 62792 37280 62801
rect 37332 62792 37334 62801
rect 37278 62727 37334 62736
rect 37278 61840 37334 61849
rect 37278 61775 37334 61784
rect 37292 61742 37320 61775
rect 37280 61736 37332 61742
rect 37280 61678 37332 61684
rect 37186 61432 37242 61441
rect 37186 61367 37242 61376
rect 37200 61266 37228 61367
rect 37188 61260 37240 61266
rect 37188 61202 37240 61208
rect 37280 60648 37332 60654
rect 37278 60616 37280 60625
rect 37332 60616 37334 60625
rect 37278 60551 37334 60560
rect 37186 60208 37242 60217
rect 37186 60143 37188 60152
rect 37240 60143 37242 60152
rect 37188 60114 37240 60120
rect 37280 60036 37332 60042
rect 37280 59978 37332 59984
rect 37292 59566 37320 59978
rect 37280 59560 37332 59566
rect 37280 59502 37332 59508
rect 37188 59084 37240 59090
rect 37188 59026 37240 59032
rect 37200 58449 37228 59026
rect 37186 58440 37242 58449
rect 37186 58375 37242 58384
rect 37188 57996 37240 58002
rect 37188 57938 37240 57944
rect 37200 57497 37228 57938
rect 37186 57488 37242 57497
rect 37186 57423 37242 57432
rect 37280 57316 37332 57322
rect 37280 57258 37332 57264
rect 37188 56908 37240 56914
rect 37188 56850 37240 56856
rect 37200 56681 37228 56850
rect 37186 56672 37242 56681
rect 37186 56607 37242 56616
rect 37292 56506 37320 57258
rect 37280 56500 37332 56506
rect 37280 56442 37332 56448
rect 37188 56432 37240 56438
rect 37188 56374 37240 56380
rect 36832 55406 36952 55434
rect 37016 56086 37136 56114
rect 36728 53780 36780 53786
rect 36728 53722 36780 53728
rect 36726 53680 36782 53689
rect 36726 53615 36728 53624
rect 36780 53615 36782 53624
rect 36728 53586 36780 53592
rect 36636 53032 36688 53038
rect 36636 52974 36688 52980
rect 36726 53000 36782 53009
rect 36726 52935 36728 52944
rect 36780 52935 36782 52944
rect 36728 52906 36780 52912
rect 36636 52896 36688 52902
rect 36636 52838 36688 52844
rect 36372 52550 36584 52578
rect 36268 51332 36320 51338
rect 36268 51274 36320 51280
rect 36268 51060 36320 51066
rect 36268 51002 36320 51008
rect 36280 49858 36308 51002
rect 36372 50930 36400 52550
rect 36452 51808 36504 51814
rect 36452 51750 36504 51756
rect 36360 50924 36412 50930
rect 36360 50866 36412 50872
rect 36280 49830 36400 49858
rect 36268 49768 36320 49774
rect 36266 49736 36268 49745
rect 36320 49736 36322 49745
rect 36266 49671 36322 49680
rect 36372 49314 36400 49830
rect 36280 49286 36400 49314
rect 36280 48793 36308 49286
rect 36360 49224 36412 49230
rect 36360 49166 36412 49172
rect 36266 48784 36322 48793
rect 36266 48719 36322 48728
rect 36268 48680 36320 48686
rect 36268 48622 36320 48628
rect 36280 48521 36308 48622
rect 36266 48512 36322 48521
rect 36372 48498 36400 49166
rect 36464 48686 36492 51750
rect 36542 51504 36598 51513
rect 36542 51439 36544 51448
rect 36596 51439 36598 51448
rect 36544 51410 36596 51416
rect 36544 51332 36596 51338
rect 36544 51274 36596 51280
rect 36556 49178 36584 51274
rect 36648 49298 36676 52838
rect 36832 52698 36860 55406
rect 36912 55344 36964 55350
rect 36912 55286 36964 55292
rect 36924 54058 36952 55286
rect 36912 54052 36964 54058
rect 36912 53994 36964 54000
rect 36912 53032 36964 53038
rect 36912 52974 36964 52980
rect 36820 52692 36872 52698
rect 36820 52634 36872 52640
rect 36728 52556 36780 52562
rect 36728 52498 36780 52504
rect 36740 52329 36768 52498
rect 36820 52420 36872 52426
rect 36820 52362 36872 52368
rect 36726 52320 36782 52329
rect 36726 52255 36782 52264
rect 36832 51338 36860 52362
rect 36820 51332 36872 51338
rect 36820 51274 36872 51280
rect 36924 51074 36952 52974
rect 36740 51046 36952 51074
rect 37016 51066 37044 56086
rect 37200 55978 37228 56374
rect 37108 55950 37228 55978
rect 37108 54584 37136 55950
rect 37188 55276 37240 55282
rect 37188 55218 37240 55224
rect 37200 54806 37228 55218
rect 37188 54800 37240 54806
rect 37188 54742 37240 54748
rect 37108 54556 37228 54584
rect 37094 54496 37150 54505
rect 37094 54431 37150 54440
rect 37108 54126 37136 54431
rect 37096 54120 37148 54126
rect 37096 54062 37148 54068
rect 37200 53990 37228 54556
rect 37188 53984 37240 53990
rect 37188 53926 37240 53932
rect 37188 52896 37240 52902
rect 37108 52856 37188 52884
rect 37004 51060 37056 51066
rect 36636 49292 36688 49298
rect 36636 49234 36688 49240
rect 36556 49150 36676 49178
rect 36544 49088 36596 49094
rect 36544 49030 36596 49036
rect 36452 48680 36504 48686
rect 36452 48622 36504 48628
rect 36372 48470 36492 48498
rect 36266 48447 36322 48456
rect 36268 48272 36320 48278
rect 36268 48214 36320 48220
rect 36280 47530 36308 48214
rect 36360 48204 36412 48210
rect 36360 48146 36412 48152
rect 36372 48113 36400 48146
rect 36358 48104 36414 48113
rect 36358 48039 36414 48048
rect 36464 47954 36492 48470
rect 36372 47926 36492 47954
rect 36372 47734 36400 47926
rect 36360 47728 36412 47734
rect 36360 47670 36412 47676
rect 36268 47524 36320 47530
rect 36268 47466 36320 47472
rect 36280 45558 36308 47466
rect 36372 47462 36400 47670
rect 36360 47456 36412 47462
rect 36360 47398 36412 47404
rect 36452 47456 36504 47462
rect 36452 47398 36504 47404
rect 36358 46744 36414 46753
rect 36358 46679 36414 46688
rect 36372 46510 36400 46679
rect 36360 46504 36412 46510
rect 36360 46446 36412 46452
rect 36360 45892 36412 45898
rect 36360 45834 36412 45840
rect 36268 45552 36320 45558
rect 36268 45494 36320 45500
rect 36268 45348 36320 45354
rect 36268 45290 36320 45296
rect 36280 42362 36308 45290
rect 36372 42770 36400 45834
rect 36464 44470 36492 47398
rect 36556 46034 36584 49030
rect 36648 48210 36676 49150
rect 36636 48204 36688 48210
rect 36636 48146 36688 48152
rect 36636 47728 36688 47734
rect 36636 47670 36688 47676
rect 36648 47598 36676 47670
rect 36636 47592 36688 47598
rect 36636 47534 36688 47540
rect 36636 47116 36688 47122
rect 36636 47058 36688 47064
rect 36544 46028 36596 46034
rect 36544 45970 36596 45976
rect 36544 45892 36596 45898
rect 36544 45834 36596 45840
rect 36556 45558 36584 45834
rect 36544 45552 36596 45558
rect 36544 45494 36596 45500
rect 36556 44810 36584 45494
rect 36544 44804 36596 44810
rect 36544 44746 36596 44752
rect 36452 44464 36504 44470
rect 36452 44406 36504 44412
rect 36450 44296 36506 44305
rect 36450 44231 36506 44240
rect 36360 42764 36412 42770
rect 36360 42706 36412 42712
rect 36464 42650 36492 44231
rect 36556 44198 36584 44746
rect 36544 44192 36596 44198
rect 36544 44134 36596 44140
rect 36542 44024 36598 44033
rect 36542 43959 36544 43968
rect 36596 43959 36598 43968
rect 36544 43930 36596 43936
rect 36544 43852 36596 43858
rect 36544 43794 36596 43800
rect 36556 43382 36584 43794
rect 36544 43376 36596 43382
rect 36544 43318 36596 43324
rect 36372 42622 36492 42650
rect 36268 42356 36320 42362
rect 36268 42298 36320 42304
rect 36176 42152 36228 42158
rect 36176 42094 36228 42100
rect 36268 42016 36320 42022
rect 36268 41958 36320 41964
rect 36174 41032 36230 41041
rect 36174 40967 36230 40976
rect 36084 40452 36136 40458
rect 36084 40394 36136 40400
rect 36084 39976 36136 39982
rect 36082 39944 36084 39953
rect 36136 39944 36138 39953
rect 36082 39879 36138 39888
rect 36082 39672 36138 39681
rect 36082 39607 36138 39616
rect 36096 39574 36124 39607
rect 36084 39568 36136 39574
rect 36084 39510 36136 39516
rect 35992 39364 36044 39370
rect 35992 39306 36044 39312
rect 36084 39364 36136 39370
rect 36084 39306 36136 39312
rect 35992 39092 36044 39098
rect 35992 39034 36044 39040
rect 36004 38418 36032 39034
rect 36096 39030 36124 39306
rect 36084 39024 36136 39030
rect 36084 38966 36136 38972
rect 36188 38654 36216 40967
rect 36280 39506 36308 41958
rect 36372 41414 36400 42622
rect 36544 42560 36596 42566
rect 36544 42502 36596 42508
rect 36372 41386 36492 41414
rect 36360 40588 36412 40594
rect 36360 40530 36412 40536
rect 36268 39500 36320 39506
rect 36268 39442 36320 39448
rect 36268 39296 36320 39302
rect 36268 39238 36320 39244
rect 36096 38626 36216 38654
rect 35992 38412 36044 38418
rect 35992 38354 36044 38360
rect 36004 38282 36032 38354
rect 35992 38276 36044 38282
rect 35992 38218 36044 38224
rect 36004 37670 36032 38218
rect 35992 37664 36044 37670
rect 35992 37606 36044 37612
rect 35992 37188 36044 37194
rect 35992 37130 36044 37136
rect 35900 36916 35952 36922
rect 35900 36858 35952 36864
rect 36004 36802 36032 37130
rect 35728 36366 35848 36394
rect 35912 36774 36032 36802
rect 35912 36378 35940 36774
rect 36096 36718 36124 38626
rect 36176 37800 36228 37806
rect 36174 37768 36176 37777
rect 36228 37768 36230 37777
rect 36174 37703 36230 37712
rect 36176 37664 36228 37670
rect 36176 37606 36228 37612
rect 36188 37097 36216 37606
rect 36174 37088 36230 37097
rect 36174 37023 36230 37032
rect 36176 36916 36228 36922
rect 36176 36858 36228 36864
rect 36084 36712 36136 36718
rect 36084 36654 36136 36660
rect 35992 36576 36044 36582
rect 35992 36518 36044 36524
rect 36084 36576 36136 36582
rect 36084 36518 36136 36524
rect 35900 36372 35952 36378
rect 35624 35148 35676 35154
rect 35624 35090 35676 35096
rect 35532 34944 35584 34950
rect 35532 34886 35584 34892
rect 35624 34944 35676 34950
rect 35624 34886 35676 34892
rect 35530 34776 35586 34785
rect 35530 34711 35586 34720
rect 35544 34542 35572 34711
rect 35532 34536 35584 34542
rect 35532 34478 35584 34484
rect 35636 34474 35664 34886
rect 35624 34468 35676 34474
rect 35624 34410 35676 34416
rect 35622 34232 35678 34241
rect 35622 34167 35678 34176
rect 35532 34128 35584 34134
rect 35530 34096 35532 34105
rect 35584 34096 35586 34105
rect 35636 34066 35664 34167
rect 35530 34031 35586 34040
rect 35624 34060 35676 34066
rect 35624 34002 35676 34008
rect 35728 33862 35756 36366
rect 35900 36314 35952 36320
rect 35898 36272 35954 36281
rect 35898 36207 35900 36216
rect 35952 36207 35954 36216
rect 35900 36178 35952 36184
rect 35808 36168 35860 36174
rect 35808 36110 35860 36116
rect 35716 33856 35768 33862
rect 35716 33798 35768 33804
rect 35452 33510 35572 33538
rect 35438 33416 35494 33425
rect 35438 33351 35494 33360
rect 35452 32978 35480 33351
rect 35440 32972 35492 32978
rect 35440 32914 35492 32920
rect 35544 32858 35572 33510
rect 35624 33312 35676 33318
rect 35624 33254 35676 33260
rect 35452 32830 35572 32858
rect 35452 30598 35480 32830
rect 35530 32056 35586 32065
rect 35530 31991 35586 32000
rect 35544 31890 35572 31991
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 35636 31754 35664 33254
rect 35544 31726 35664 31754
rect 35440 30592 35492 30598
rect 35440 30534 35492 30540
rect 35440 29572 35492 29578
rect 35440 29514 35492 29520
rect 35348 26852 35400 26858
rect 35348 26794 35400 26800
rect 35452 25378 35480 29514
rect 35544 26994 35572 31726
rect 35820 31634 35848 36110
rect 35900 35828 35952 35834
rect 35900 35770 35952 35776
rect 35912 35630 35940 35770
rect 35900 35624 35952 35630
rect 35900 35566 35952 35572
rect 35900 35216 35952 35222
rect 35900 35158 35952 35164
rect 35912 34513 35940 35158
rect 35898 34504 35954 34513
rect 35898 34439 35954 34448
rect 35900 34128 35952 34134
rect 35900 34070 35952 34076
rect 35912 33697 35940 34070
rect 35898 33688 35954 33697
rect 35898 33623 35954 33632
rect 35900 33584 35952 33590
rect 35900 33526 35952 33532
rect 35912 32366 35940 33526
rect 35900 32360 35952 32366
rect 35900 32302 35952 32308
rect 35900 31748 35952 31754
rect 35900 31690 35952 31696
rect 35636 31606 35848 31634
rect 35532 26988 35584 26994
rect 35532 26930 35584 26936
rect 35532 26852 35584 26858
rect 35532 26794 35584 26800
rect 35360 25350 35480 25378
rect 35256 25288 35308 25294
rect 35256 25230 35308 25236
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35360 22094 35388 25350
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35268 22066 35388 22094
rect 35268 21962 35296 22066
rect 35256 21956 35308 21962
rect 35256 21898 35308 21904
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35452 20534 35480 25230
rect 35440 20528 35492 20534
rect 35440 20470 35492 20476
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35544 16250 35572 26794
rect 35532 16244 35584 16250
rect 35532 16186 35584 16192
rect 35256 16040 35308 16046
rect 35256 15982 35308 15988
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 35268 6866 35296 15982
rect 35636 15162 35664 31606
rect 35806 30832 35862 30841
rect 35806 30767 35808 30776
rect 35860 30767 35862 30776
rect 35808 30738 35860 30744
rect 35716 30592 35768 30598
rect 35716 30534 35768 30540
rect 35624 15156 35676 15162
rect 35624 15098 35676 15104
rect 35728 15094 35756 30534
rect 35808 29708 35860 29714
rect 35808 29650 35860 29656
rect 35820 29481 35848 29650
rect 35806 29472 35862 29481
rect 35806 29407 35862 29416
rect 35912 29017 35940 31690
rect 36004 30598 36032 36518
rect 36096 33454 36124 36518
rect 36188 34785 36216 36858
rect 36280 35306 36308 39238
rect 36372 37466 36400 40530
rect 36360 37460 36412 37466
rect 36360 37402 36412 37408
rect 36360 37324 36412 37330
rect 36360 37266 36412 37272
rect 36372 36825 36400 37266
rect 36358 36816 36414 36825
rect 36358 36751 36414 36760
rect 36464 36718 36492 41386
rect 36556 41002 36584 42502
rect 36648 41138 36676 47058
rect 36740 46170 36768 51046
rect 37004 51002 37056 51008
rect 36820 50856 36872 50862
rect 36820 50798 36872 50804
rect 36832 49978 36860 50798
rect 36912 50788 36964 50794
rect 36912 50730 36964 50736
rect 36924 50522 36952 50730
rect 37004 50720 37056 50726
rect 37004 50662 37056 50668
rect 37016 50522 37044 50662
rect 36912 50516 36964 50522
rect 36912 50458 36964 50464
rect 37004 50516 37056 50522
rect 37004 50458 37056 50464
rect 36912 50380 36964 50386
rect 36912 50322 36964 50328
rect 36820 49972 36872 49978
rect 36820 49914 36872 49920
rect 36820 49768 36872 49774
rect 36820 49710 36872 49716
rect 36832 47258 36860 49710
rect 36924 48890 36952 50322
rect 37016 49688 37044 50458
rect 37108 49910 37136 52856
rect 37188 52838 37240 52844
rect 37188 52556 37240 52562
rect 37188 52498 37240 52504
rect 37200 51921 37228 52498
rect 37186 51912 37242 51921
rect 37186 51847 37242 51856
rect 37292 50998 37320 56442
rect 37384 55214 37412 67594
rect 37464 62688 37516 62694
rect 37464 62630 37516 62636
rect 37476 62529 37504 62630
rect 37462 62520 37518 62529
rect 37462 62455 37518 62464
rect 37464 60512 37516 60518
rect 37464 60454 37516 60460
rect 37476 60246 37504 60454
rect 37464 60240 37516 60246
rect 37464 60182 37516 60188
rect 37568 58478 37596 81670
rect 37752 79898 37780 84390
rect 37936 83881 37964 84526
rect 37922 83872 37978 83881
rect 37922 83807 37978 83816
rect 37924 83496 37976 83502
rect 37924 83438 37976 83444
rect 37936 83065 37964 83438
rect 37922 83056 37978 83065
rect 37922 82991 37978 83000
rect 37924 82408 37976 82414
rect 37924 82350 37976 82356
rect 37936 81705 37964 82350
rect 37922 81696 37978 81705
rect 37922 81631 37978 81640
rect 37924 81320 37976 81326
rect 37924 81262 37976 81268
rect 37936 80889 37964 81262
rect 37922 80880 37978 80889
rect 37922 80815 37978 80824
rect 38028 80646 38056 84918
rect 38200 84788 38252 84794
rect 38200 84730 38252 84736
rect 38108 83360 38160 83366
rect 38108 83302 38160 83308
rect 38016 80640 38068 80646
rect 38016 80582 38068 80588
rect 37924 80232 37976 80238
rect 37924 80174 37976 80180
rect 37740 79892 37792 79898
rect 37740 79834 37792 79840
rect 37936 79529 37964 80174
rect 37922 79520 37978 79529
rect 37922 79455 37978 79464
rect 37924 79144 37976 79150
rect 37922 79112 37924 79121
rect 37976 79112 37978 79121
rect 37922 79047 37978 79056
rect 38120 78810 38148 83302
rect 38212 81394 38240 84730
rect 38200 81388 38252 81394
rect 38200 81330 38252 81336
rect 38108 78804 38160 78810
rect 38108 78746 38160 78752
rect 37924 77988 37976 77994
rect 37924 77930 37976 77936
rect 37936 77897 37964 77930
rect 37922 77888 37978 77897
rect 37922 77823 37978 77832
rect 37922 76936 37978 76945
rect 37922 76871 37924 76880
rect 37976 76871 37978 76880
rect 37924 76842 37976 76848
rect 38016 76832 38068 76838
rect 38016 76774 38068 76780
rect 38028 76634 38056 76774
rect 38016 76628 38068 76634
rect 38016 76570 38068 76576
rect 38304 75954 38332 114922
rect 38396 114102 38424 119200
rect 38384 114096 38436 114102
rect 38384 114038 38436 114044
rect 38580 113626 38608 119200
rect 38856 116618 38884 119200
rect 39040 117094 39068 119200
rect 39028 117088 39080 117094
rect 39028 117030 39080 117036
rect 38844 116612 38896 116618
rect 38844 116554 38896 116560
rect 39224 114646 39252 119200
rect 39500 115530 39528 119200
rect 39488 115524 39540 115530
rect 39488 115466 39540 115472
rect 39212 114640 39264 114646
rect 39212 114582 39264 114588
rect 39684 114510 39712 119200
rect 39672 114504 39724 114510
rect 39672 114446 39724 114452
rect 38568 113620 38620 113626
rect 38568 113562 38620 113568
rect 39868 112470 39896 119200
rect 39856 112464 39908 112470
rect 39856 112406 39908 112412
rect 38660 109540 38712 109546
rect 38660 109482 38712 109488
rect 38384 109472 38436 109478
rect 38384 109414 38436 109420
rect 38396 94586 38424 109414
rect 38476 106820 38528 106826
rect 38476 106762 38528 106768
rect 38384 94580 38436 94586
rect 38384 94522 38436 94528
rect 38384 93152 38436 93158
rect 38384 93094 38436 93100
rect 38396 89146 38424 93094
rect 38488 89622 38516 106762
rect 38672 99374 38700 109482
rect 38672 99346 38792 99374
rect 38660 94784 38712 94790
rect 38660 94726 38712 94732
rect 38568 94444 38620 94450
rect 38568 94386 38620 94392
rect 38476 89616 38528 89622
rect 38476 89558 38528 89564
rect 38384 89140 38436 89146
rect 38384 89082 38436 89088
rect 38580 89010 38608 94386
rect 38568 89004 38620 89010
rect 38568 88946 38620 88952
rect 38384 88936 38436 88942
rect 38384 88878 38436 88884
rect 38396 81870 38424 88878
rect 38672 84522 38700 94726
rect 38764 86737 38792 99346
rect 38844 94580 38896 94586
rect 38844 94522 38896 94528
rect 38750 86728 38806 86737
rect 38750 86663 38806 86672
rect 38660 84516 38712 84522
rect 38660 84458 38712 84464
rect 38384 81864 38436 81870
rect 38384 81806 38436 81812
rect 38856 80345 38884 94522
rect 38936 92540 38988 92546
rect 38936 92482 38988 92488
rect 38948 92449 38976 92482
rect 38934 92440 38990 92449
rect 38934 92375 38990 92384
rect 39212 82544 39264 82550
rect 39212 82486 39264 82492
rect 39028 80368 39080 80374
rect 38842 80336 38898 80345
rect 39028 80310 39080 80316
rect 38842 80271 38898 80280
rect 38292 75948 38344 75954
rect 38292 75890 38344 75896
rect 37924 75812 37976 75818
rect 37924 75754 37976 75760
rect 37936 75721 37964 75754
rect 37922 75712 37978 75721
rect 37922 75647 37978 75656
rect 37922 74760 37978 74769
rect 37922 74695 37924 74704
rect 37976 74695 37978 74704
rect 37924 74666 37976 74672
rect 37924 73636 37976 73642
rect 37924 73578 37976 73584
rect 37936 73545 37964 73578
rect 38016 73568 38068 73574
rect 37922 73536 37978 73545
rect 38016 73510 38068 73516
rect 37922 73471 37978 73480
rect 38028 73302 38056 73510
rect 38016 73296 38068 73302
rect 38016 73238 38068 73244
rect 37922 72720 37978 72729
rect 37922 72655 37978 72664
rect 37936 72622 37964 72655
rect 37924 72616 37976 72622
rect 37924 72558 37976 72564
rect 37648 72480 37700 72486
rect 37648 72422 37700 72428
rect 37556 58472 37608 58478
rect 37556 58414 37608 58420
rect 37556 57248 37608 57254
rect 37556 57190 37608 57196
rect 37372 55208 37424 55214
rect 37372 55150 37424 55156
rect 37464 55072 37516 55078
rect 37464 55014 37516 55020
rect 37372 53644 37424 53650
rect 37372 53586 37424 53592
rect 37384 53281 37412 53586
rect 37370 53272 37426 53281
rect 37370 53207 37426 53216
rect 37372 51468 37424 51474
rect 37372 51410 37424 51416
rect 37384 51105 37412 51410
rect 37370 51096 37426 51105
rect 37370 51031 37426 51040
rect 37280 50992 37332 50998
rect 37280 50934 37332 50940
rect 37476 50930 37504 55014
rect 37568 54670 37596 57190
rect 37556 54664 37608 54670
rect 37556 54606 37608 54612
rect 37556 53984 37608 53990
rect 37556 53926 37608 53932
rect 37464 50924 37516 50930
rect 37464 50866 37516 50872
rect 37372 50720 37424 50726
rect 37568 50674 37596 53926
rect 37372 50662 37424 50668
rect 37384 49978 37412 50662
rect 37476 50646 37596 50674
rect 37476 50250 37504 50646
rect 37556 50312 37608 50318
rect 37556 50254 37608 50260
rect 37464 50244 37516 50250
rect 37464 50186 37516 50192
rect 37372 49972 37424 49978
rect 37372 49914 37424 49920
rect 37096 49904 37148 49910
rect 37096 49846 37148 49852
rect 37372 49836 37424 49842
rect 37568 49824 37596 50254
rect 37424 49796 37596 49824
rect 37372 49778 37424 49784
rect 37096 49700 37148 49706
rect 37016 49660 37096 49688
rect 37016 49298 37044 49660
rect 37096 49642 37148 49648
rect 37384 49366 37412 49778
rect 37556 49428 37608 49434
rect 37556 49370 37608 49376
rect 37372 49360 37424 49366
rect 37372 49302 37424 49308
rect 37004 49292 37056 49298
rect 37004 49234 37056 49240
rect 36912 48884 36964 48890
rect 36912 48826 36964 48832
rect 37016 48618 37044 49234
rect 37280 49088 37332 49094
rect 37280 49030 37332 49036
rect 37292 48822 37320 49030
rect 37280 48816 37332 48822
rect 37280 48758 37332 48764
rect 37384 48754 37412 49302
rect 37372 48748 37424 48754
rect 37372 48690 37424 48696
rect 36912 48612 36964 48618
rect 36912 48554 36964 48560
rect 37004 48612 37056 48618
rect 37004 48554 37056 48560
rect 36820 47252 36872 47258
rect 36820 47194 36872 47200
rect 36924 47138 36952 48554
rect 36832 47110 36952 47138
rect 36728 46164 36780 46170
rect 36728 46106 36780 46112
rect 36728 46028 36780 46034
rect 36728 45970 36780 45976
rect 36740 43450 36768 45970
rect 36832 45490 36860 47110
rect 36912 46912 36964 46918
rect 36912 46854 36964 46860
rect 36924 46646 36952 46854
rect 36912 46640 36964 46646
rect 36912 46582 36964 46588
rect 36912 46028 36964 46034
rect 36912 45970 36964 45976
rect 36820 45484 36872 45490
rect 36820 45426 36872 45432
rect 36924 45370 36952 45970
rect 36832 45354 36952 45370
rect 36820 45348 36952 45354
rect 36872 45342 36952 45348
rect 36820 45290 36872 45296
rect 36832 44946 36860 45290
rect 36820 44940 36872 44946
rect 36820 44882 36872 44888
rect 36832 44266 36860 44882
rect 36912 44464 36964 44470
rect 36912 44406 36964 44412
rect 36820 44260 36872 44266
rect 36820 44202 36872 44208
rect 36832 43897 36860 44202
rect 36818 43888 36874 43897
rect 36818 43823 36874 43832
rect 36728 43444 36780 43450
rect 36728 43386 36780 43392
rect 36728 42628 36780 42634
rect 36728 42570 36780 42576
rect 36820 42628 36872 42634
rect 36820 42570 36872 42576
rect 36740 41682 36768 42570
rect 36832 42226 36860 42570
rect 36820 42220 36872 42226
rect 36820 42162 36872 42168
rect 36728 41676 36780 41682
rect 36728 41618 36780 41624
rect 36820 41608 36872 41614
rect 36820 41550 36872 41556
rect 36924 41562 36952 44406
rect 37016 43450 37044 48554
rect 37096 48544 37148 48550
rect 37096 48486 37148 48492
rect 37004 43444 37056 43450
rect 37004 43386 37056 43392
rect 37108 43330 37136 48486
rect 37280 48272 37332 48278
rect 37200 48220 37280 48226
rect 37200 48214 37332 48220
rect 37200 48198 37320 48214
rect 37200 47734 37228 48198
rect 37372 48000 37424 48006
rect 37372 47942 37424 47948
rect 37188 47728 37240 47734
rect 37188 47670 37240 47676
rect 37280 47592 37332 47598
rect 37280 47534 37332 47540
rect 37188 47524 37240 47530
rect 37188 47466 37240 47472
rect 37200 46442 37228 47466
rect 37292 47054 37320 47534
rect 37280 47048 37332 47054
rect 37280 46990 37332 46996
rect 37188 46436 37240 46442
rect 37188 46378 37240 46384
rect 37280 46368 37332 46374
rect 37280 46310 37332 46316
rect 37186 45792 37242 45801
rect 37186 45727 37242 45736
rect 37200 45626 37228 45727
rect 37188 45620 37240 45626
rect 37188 45562 37240 45568
rect 37188 45484 37240 45490
rect 37188 45426 37240 45432
rect 37200 44538 37228 45426
rect 37188 44532 37240 44538
rect 37188 44474 37240 44480
rect 37186 44432 37242 44441
rect 37186 44367 37188 44376
rect 37240 44367 37242 44376
rect 37188 44338 37240 44344
rect 37188 43988 37240 43994
rect 37188 43930 37240 43936
rect 37016 43302 37136 43330
rect 37016 41682 37044 43302
rect 37096 43172 37148 43178
rect 37096 43114 37148 43120
rect 37108 41750 37136 43114
rect 37200 43110 37228 43930
rect 37292 43722 37320 46310
rect 37384 45121 37412 47942
rect 37464 47456 37516 47462
rect 37464 47398 37516 47404
rect 37370 45112 37426 45121
rect 37370 45047 37426 45056
rect 37372 44192 37424 44198
rect 37372 44134 37424 44140
rect 37280 43716 37332 43722
rect 37280 43658 37332 43664
rect 37188 43104 37240 43110
rect 37188 43046 37240 43052
rect 37280 42764 37332 42770
rect 37200 42724 37280 42752
rect 37096 41744 37148 41750
rect 37096 41686 37148 41692
rect 37004 41676 37056 41682
rect 37004 41618 37056 41624
rect 36728 41200 36780 41206
rect 36728 41142 36780 41148
rect 36636 41132 36688 41138
rect 36636 41074 36688 41080
rect 36544 40996 36596 41002
rect 36544 40938 36596 40944
rect 36636 40996 36688 41002
rect 36636 40938 36688 40944
rect 36556 40662 36584 40938
rect 36544 40656 36596 40662
rect 36544 40598 36596 40604
rect 36556 39982 36584 40598
rect 36648 40594 36676 40938
rect 36740 40594 36768 41142
rect 36636 40588 36688 40594
rect 36636 40530 36688 40536
rect 36728 40588 36780 40594
rect 36728 40530 36780 40536
rect 36544 39976 36596 39982
rect 36544 39918 36596 39924
rect 36556 39574 36584 39918
rect 36648 39914 36676 40530
rect 36636 39908 36688 39914
rect 36636 39850 36688 39856
rect 36544 39568 36596 39574
rect 36544 39510 36596 39516
rect 36556 39137 36584 39510
rect 36648 39506 36676 39850
rect 36728 39636 36780 39642
rect 36728 39578 36780 39584
rect 36636 39500 36688 39506
rect 36636 39442 36688 39448
rect 36542 39128 36598 39137
rect 36542 39063 36598 39072
rect 36544 38956 36596 38962
rect 36544 38898 36596 38904
rect 36556 38536 36584 38898
rect 36648 38826 36676 39442
rect 36740 38978 36768 39578
rect 36740 38950 36773 38978
rect 36745 38876 36773 38950
rect 36740 38848 36773 38876
rect 36636 38820 36688 38826
rect 36636 38762 36688 38768
rect 36556 38508 36676 38536
rect 36544 38412 36596 38418
rect 36544 38354 36596 38360
rect 36360 36712 36412 36718
rect 36360 36654 36412 36660
rect 36452 36712 36504 36718
rect 36452 36654 36504 36660
rect 36372 36242 36400 36654
rect 36360 36236 36412 36242
rect 36360 36178 36412 36184
rect 36372 35816 36400 36178
rect 36450 35864 36506 35873
rect 36372 35808 36450 35816
rect 36372 35799 36506 35808
rect 36372 35788 36492 35799
rect 36358 35728 36414 35737
rect 36464 35698 36492 35788
rect 36358 35663 36414 35672
rect 36452 35692 36504 35698
rect 36372 35630 36400 35663
rect 36452 35634 36504 35640
rect 36360 35624 36412 35630
rect 36360 35566 36412 35572
rect 36280 35278 36405 35306
rect 36377 35222 36405 35278
rect 36365 35216 36417 35222
rect 36365 35158 36417 35164
rect 36268 35148 36320 35154
rect 36268 35090 36320 35096
rect 36372 35142 36405 35158
rect 36452 35148 36504 35154
rect 36174 34776 36230 34785
rect 36174 34711 36230 34720
rect 36174 34504 36230 34513
rect 36174 34439 36230 34448
rect 36188 33590 36216 34439
rect 36176 33584 36228 33590
rect 36176 33526 36228 33532
rect 36084 33448 36136 33454
rect 36084 33390 36136 33396
rect 36176 33448 36228 33454
rect 36176 33390 36228 33396
rect 36082 33144 36138 33153
rect 36082 33079 36138 33088
rect 36096 32978 36124 33079
rect 36084 32972 36136 32978
rect 36084 32914 36136 32920
rect 36188 32008 36216 33390
rect 36096 31980 36216 32008
rect 35992 30592 36044 30598
rect 35992 30534 36044 30540
rect 35990 30288 36046 30297
rect 35990 30223 36046 30232
rect 36004 30190 36032 30223
rect 35992 30184 36044 30190
rect 35992 30126 36044 30132
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 36004 29238 36032 29446
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 35992 29096 36044 29102
rect 36096 29073 36124 31980
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 36188 31249 36216 31826
rect 36174 31240 36230 31249
rect 36174 31175 36230 31184
rect 36280 30938 36308 35090
rect 36372 34542 36400 35142
rect 36452 35090 36504 35096
rect 36360 34536 36412 34542
rect 36360 34478 36412 34484
rect 36464 34538 36492 35090
rect 36372 34134 36400 34478
rect 36464 34474 36493 34538
rect 36453 34468 36505 34474
rect 36453 34410 36505 34416
rect 36360 34128 36412 34134
rect 36360 34070 36412 34076
rect 36372 33386 36400 34070
rect 36464 34066 36492 34410
rect 36452 34060 36504 34066
rect 36452 34002 36504 34008
rect 36464 33386 36492 34002
rect 36360 33380 36412 33386
rect 36360 33322 36412 33328
rect 36452 33380 36504 33386
rect 36452 33322 36504 33328
rect 36372 33046 36400 33322
rect 36360 33040 36412 33046
rect 36360 32982 36412 32988
rect 36464 32978 36492 33322
rect 36556 33114 36584 38354
rect 36648 38298 36676 38508
rect 36740 38418 36768 38848
rect 36728 38412 36780 38418
rect 36728 38354 36780 38360
rect 36648 38270 36768 38298
rect 36636 38208 36688 38214
rect 36636 38150 36688 38156
rect 36648 36281 36676 38150
rect 36634 36272 36690 36281
rect 36634 36207 36690 36216
rect 36636 34944 36688 34950
rect 36636 34886 36688 34892
rect 36648 34678 36676 34886
rect 36636 34672 36688 34678
rect 36636 34614 36688 34620
rect 36740 34490 36768 38270
rect 36832 36378 36860 41550
rect 36924 41534 37044 41562
rect 36912 40928 36964 40934
rect 36912 40870 36964 40876
rect 36924 40089 36952 40870
rect 37016 40730 37044 41534
rect 37108 41041 37136 41686
rect 37094 41032 37150 41041
rect 37094 40967 37150 40976
rect 37096 40928 37148 40934
rect 37096 40870 37148 40876
rect 37004 40724 37056 40730
rect 37004 40666 37056 40672
rect 36910 40080 36966 40089
rect 36910 40015 36966 40024
rect 36912 39840 36964 39846
rect 36912 39782 36964 39788
rect 36924 39681 36952 39782
rect 36910 39672 36966 39681
rect 36910 39607 36966 39616
rect 36910 39536 36966 39545
rect 36910 39471 36966 39480
rect 36924 38944 36952 39471
rect 37108 39098 37136 40870
rect 37096 39092 37148 39098
rect 37096 39034 37148 39040
rect 36924 38916 37136 38944
rect 37108 38758 37136 38916
rect 37096 38752 37148 38758
rect 37096 38694 37148 38700
rect 36910 38448 36966 38457
rect 36910 38383 36912 38392
rect 36964 38383 36966 38392
rect 36912 38354 36964 38360
rect 36910 38040 36966 38049
rect 36910 37975 36912 37984
rect 36964 37975 36966 37984
rect 36912 37946 36964 37952
rect 37096 37732 37148 37738
rect 37096 37674 37148 37680
rect 36912 37120 36964 37126
rect 36912 37062 36964 37068
rect 36820 36372 36872 36378
rect 36820 36314 36872 36320
rect 36832 35698 36860 36314
rect 36820 35692 36872 35698
rect 36820 35634 36872 35640
rect 36820 35556 36872 35562
rect 36820 35498 36872 35504
rect 36648 34462 36768 34490
rect 36648 33946 36676 34462
rect 36728 34400 36780 34406
rect 36728 34342 36780 34348
rect 36740 34202 36768 34342
rect 36728 34196 36780 34202
rect 36728 34138 36780 34144
rect 36726 34096 36782 34105
rect 36726 34031 36728 34040
rect 36780 34031 36782 34040
rect 36728 34002 36780 34008
rect 36648 33918 36768 33946
rect 36634 33688 36690 33697
rect 36634 33623 36690 33632
rect 36544 33108 36596 33114
rect 36544 33050 36596 33056
rect 36452 32972 36504 32978
rect 36452 32914 36504 32920
rect 36544 32972 36596 32978
rect 36544 32914 36596 32920
rect 36360 32768 36412 32774
rect 36360 32710 36412 32716
rect 36268 30932 36320 30938
rect 36268 30874 36320 30880
rect 36372 30666 36400 32710
rect 36464 32570 36492 32914
rect 36556 32570 36584 32914
rect 36452 32564 36504 32570
rect 36452 32506 36504 32512
rect 36544 32564 36596 32570
rect 36544 32506 36596 32512
rect 36544 32428 36596 32434
rect 36544 32370 36596 32376
rect 36452 31952 36504 31958
rect 36452 31894 36504 31900
rect 36464 31482 36492 31894
rect 36556 31890 36584 32370
rect 36544 31884 36596 31890
rect 36544 31826 36596 31832
rect 36544 31680 36596 31686
rect 36544 31622 36596 31628
rect 36452 31476 36504 31482
rect 36452 31418 36504 31424
rect 36360 30660 36412 30666
rect 36360 30602 36412 30608
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 36188 30190 36216 30534
rect 36176 30184 36228 30190
rect 36360 30184 36412 30190
rect 36228 30144 36308 30172
rect 36176 30126 36228 30132
rect 36176 29844 36228 29850
rect 36176 29786 36228 29792
rect 36188 29170 36216 29786
rect 36280 29714 36308 30144
rect 36360 30126 36412 30132
rect 36372 29782 36400 30126
rect 36452 30048 36504 30054
rect 36452 29990 36504 29996
rect 36360 29776 36412 29782
rect 36360 29718 36412 29724
rect 36268 29708 36320 29714
rect 36268 29650 36320 29656
rect 36176 29164 36228 29170
rect 36176 29106 36228 29112
rect 35992 29038 36044 29044
rect 36082 29064 36138 29073
rect 35898 29008 35954 29017
rect 35808 28960 35860 28966
rect 36004 28994 36032 29038
rect 36082 28999 36138 29008
rect 36176 29028 36228 29034
rect 36004 28966 36033 28994
rect 36280 29016 36308 29650
rect 36228 28988 36308 29016
rect 36372 29016 36400 29718
rect 36464 29714 36492 29990
rect 36452 29708 36504 29714
rect 36452 29650 36504 29656
rect 36452 29028 36504 29034
rect 36372 28988 36452 29016
rect 36176 28970 36228 28976
rect 35898 28943 35954 28952
rect 36005 28948 36033 28966
rect 36005 28920 36124 28948
rect 35808 28902 35860 28908
rect 35820 20806 35848 28902
rect 36096 28778 36124 28920
rect 35900 28756 35952 28762
rect 35900 28698 35952 28704
rect 36004 28750 36124 28778
rect 35912 28014 35940 28698
rect 35900 28008 35952 28014
rect 35900 27950 35952 27956
rect 35900 27532 35952 27538
rect 35900 27474 35952 27480
rect 35808 20800 35860 20806
rect 35808 20742 35860 20748
rect 35716 15088 35768 15094
rect 35716 15030 35768 15036
rect 35256 6860 35308 6866
rect 35256 6802 35308 6808
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35624 5568 35676 5574
rect 35624 5510 35676 5516
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35532 5228 35584 5234
rect 35532 5170 35584 5176
rect 35440 4480 35492 4486
rect 35440 4422 35492 4428
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 34704 2576 34756 2582
rect 34704 2518 34756 2524
rect 34796 2508 34848 2514
rect 34796 2450 34848 2456
rect 34808 800 34836 2450
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35268 1578 35296 2926
rect 35360 2922 35388 3878
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 35176 1550 35296 1578
rect 35176 800 35204 1550
rect 35452 800 35480 4422
rect 35544 2650 35572 5170
rect 35636 3126 35664 5510
rect 35808 4684 35860 4690
rect 35808 4626 35860 4632
rect 35820 3641 35848 4626
rect 35912 3738 35940 27474
rect 36004 21690 36032 28750
rect 36084 28688 36136 28694
rect 36084 28630 36136 28636
rect 36096 27130 36124 28630
rect 36188 28626 36216 28970
rect 36372 28914 36400 28988
rect 36452 28970 36504 28976
rect 36280 28886 36400 28914
rect 36280 28694 36308 28886
rect 36358 28792 36414 28801
rect 36358 28727 36414 28736
rect 36268 28688 36320 28694
rect 36268 28630 36320 28636
rect 36176 28620 36228 28626
rect 36176 28562 36228 28568
rect 36280 28614 36316 28630
rect 36188 27946 36216 28562
rect 36280 28014 36308 28614
rect 36377 28608 36405 28727
rect 36372 28580 36405 28608
rect 36268 28008 36320 28014
rect 36268 27950 36320 27956
rect 36176 27940 36228 27946
rect 36176 27882 36228 27888
rect 36280 27674 36308 27950
rect 36268 27668 36320 27674
rect 36268 27610 36320 27616
rect 36372 27538 36400 28580
rect 36452 28144 36504 28150
rect 36452 28086 36504 28092
rect 36360 27532 36412 27538
rect 36360 27474 36412 27480
rect 36084 27124 36136 27130
rect 36084 27066 36136 27072
rect 35992 21684 36044 21690
rect 35992 21626 36044 21632
rect 36464 20942 36492 28086
rect 36556 26042 36584 31622
rect 36648 28642 36676 33623
rect 36740 32570 36768 33918
rect 36728 32564 36780 32570
rect 36728 32506 36780 32512
rect 36728 32360 36780 32366
rect 36728 32302 36780 32308
rect 36740 31754 36768 32302
rect 36728 31748 36780 31754
rect 36728 31690 36780 31696
rect 36728 30796 36780 30802
rect 36728 30738 36780 30744
rect 36740 30433 36768 30738
rect 36726 30424 36782 30433
rect 36726 30359 36782 30368
rect 36728 30048 36780 30054
rect 36728 29990 36780 29996
rect 36740 28762 36768 29990
rect 36728 28756 36780 28762
rect 36728 28698 36780 28704
rect 36648 28614 36768 28642
rect 36636 28552 36688 28558
rect 36636 28494 36688 28500
rect 36544 26036 36596 26042
rect 36544 25978 36596 25984
rect 36648 25242 36676 28494
rect 36740 28218 36768 28614
rect 36728 28212 36780 28218
rect 36728 28154 36780 28160
rect 36832 25362 36860 35498
rect 36924 33930 36952 37062
rect 37004 36712 37056 36718
rect 37004 36654 37056 36660
rect 36912 33924 36964 33930
rect 36912 33866 36964 33872
rect 36912 32360 36964 32366
rect 36912 32302 36964 32308
rect 36924 31657 36952 32302
rect 37016 31686 37044 36654
rect 37108 32008 37136 37674
rect 37200 34202 37228 42724
rect 37280 42706 37332 42712
rect 37280 42560 37332 42566
rect 37280 42502 37332 42508
rect 37292 40050 37320 42502
rect 37384 42362 37412 44134
rect 37476 43246 37504 47398
rect 37568 43994 37596 49370
rect 37556 43988 37608 43994
rect 37556 43930 37608 43936
rect 37554 43888 37610 43897
rect 37554 43823 37610 43832
rect 37568 43790 37596 43823
rect 37556 43784 37608 43790
rect 37556 43726 37608 43732
rect 37464 43240 37516 43246
rect 37464 43182 37516 43188
rect 37372 42356 37424 42362
rect 37372 42298 37424 42304
rect 37464 42288 37516 42294
rect 37464 42230 37516 42236
rect 37372 42152 37424 42158
rect 37372 42094 37424 42100
rect 37384 41478 37412 42094
rect 37372 41472 37424 41478
rect 37372 41414 37424 41420
rect 37384 41206 37412 41414
rect 37372 41200 37424 41206
rect 37372 41142 37424 41148
rect 37372 41064 37424 41070
rect 37372 41006 37424 41012
rect 37280 40044 37332 40050
rect 37280 39986 37332 39992
rect 37280 38956 37332 38962
rect 37280 38898 37332 38904
rect 37292 38865 37320 38898
rect 37278 38856 37334 38865
rect 37278 38791 37334 38800
rect 37280 38752 37332 38758
rect 37280 38694 37332 38700
rect 37292 35698 37320 38694
rect 37384 38350 37412 41006
rect 37476 41002 37504 42230
rect 37568 41818 37596 43726
rect 37556 41812 37608 41818
rect 37556 41754 37608 41760
rect 37556 41064 37608 41070
rect 37556 41006 37608 41012
rect 37464 40996 37516 41002
rect 37464 40938 37516 40944
rect 37568 40186 37596 41006
rect 37556 40180 37608 40186
rect 37556 40122 37608 40128
rect 37556 39840 37608 39846
rect 37556 39782 37608 39788
rect 37464 38888 37516 38894
rect 37464 38830 37516 38836
rect 37372 38344 37424 38350
rect 37372 38286 37424 38292
rect 37372 37664 37424 37670
rect 37372 37606 37424 37612
rect 37384 37398 37412 37606
rect 37372 37392 37424 37398
rect 37372 37334 37424 37340
rect 37384 36650 37412 37334
rect 37372 36644 37424 36650
rect 37372 36586 37424 36592
rect 37370 36544 37426 36553
rect 37370 36479 37426 36488
rect 37280 35692 37332 35698
rect 37280 35634 37332 35640
rect 37384 35306 37412 36479
rect 37476 36310 37504 38830
rect 37464 36304 37516 36310
rect 37464 36246 37516 36252
rect 37462 35864 37518 35873
rect 37568 35834 37596 39782
rect 37462 35799 37518 35808
rect 37556 35828 37608 35834
rect 37476 35562 37504 35799
rect 37556 35770 37608 35776
rect 37464 35556 37516 35562
rect 37464 35498 37516 35504
rect 37292 35278 37412 35306
rect 37292 35154 37320 35278
rect 37280 35148 37332 35154
rect 37280 35090 37332 35096
rect 37188 34196 37240 34202
rect 37188 34138 37240 34144
rect 37292 34082 37320 35090
rect 37462 35048 37518 35057
rect 37462 34983 37518 34992
rect 37200 34054 37320 34082
rect 37372 34060 37424 34066
rect 37200 32774 37228 34054
rect 37372 34002 37424 34008
rect 37384 33833 37412 34002
rect 37370 33824 37426 33833
rect 37370 33759 37426 33768
rect 37476 33454 37504 34983
rect 37556 34672 37608 34678
rect 37556 34614 37608 34620
rect 37464 33448 37516 33454
rect 37464 33390 37516 33396
rect 37370 33008 37426 33017
rect 37370 32943 37372 32952
rect 37424 32943 37426 32952
rect 37372 32914 37424 32920
rect 37188 32768 37240 32774
rect 37188 32710 37240 32716
rect 37464 32224 37516 32230
rect 37464 32166 37516 32172
rect 37188 32020 37240 32026
rect 37108 31980 37188 32008
rect 37188 31962 37240 31968
rect 37188 31884 37240 31890
rect 37108 31844 37188 31872
rect 37004 31680 37056 31686
rect 36910 31648 36966 31657
rect 37004 31622 37056 31628
rect 36910 31583 36966 31592
rect 36912 31272 36964 31278
rect 36912 31214 36964 31220
rect 36820 25356 36872 25362
rect 36820 25298 36872 25304
rect 36648 25214 36860 25242
rect 36728 25152 36780 25158
rect 36728 25094 36780 25100
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36544 19984 36596 19990
rect 36544 19926 36596 19932
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 36096 6914 36124 18022
rect 36176 15972 36228 15978
rect 36176 15914 36228 15920
rect 36004 6886 36124 6914
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 35806 3632 35862 3641
rect 35716 3596 35768 3602
rect 35806 3567 35862 3576
rect 35716 3538 35768 3544
rect 35624 3120 35676 3126
rect 35624 3062 35676 3068
rect 35532 2644 35584 2650
rect 35532 2586 35584 2592
rect 35728 800 35756 3538
rect 36004 3058 36032 6886
rect 36084 5568 36136 5574
rect 36084 5510 36136 5516
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36096 2802 36124 5510
rect 36188 4758 36216 15914
rect 36556 15706 36584 19926
rect 36544 15700 36596 15706
rect 36544 15642 36596 15648
rect 36648 12442 36676 24074
rect 36740 17338 36768 25094
rect 36832 20602 36860 25214
rect 36820 20596 36872 20602
rect 36820 20538 36872 20544
rect 36924 19242 36952 31214
rect 37004 31136 37056 31142
rect 37004 31078 37056 31084
rect 37016 28490 37044 31078
rect 37004 28484 37056 28490
rect 37004 28426 37056 28432
rect 37004 27872 37056 27878
rect 37004 27814 37056 27820
rect 36912 19236 36964 19242
rect 36912 19178 36964 19184
rect 37016 18970 37044 27814
rect 37108 21622 37136 31844
rect 37188 31826 37240 31832
rect 37372 31680 37424 31686
rect 37372 31622 37424 31628
rect 37280 31204 37332 31210
rect 37280 31146 37332 31152
rect 37188 31136 37240 31142
rect 37188 31078 37240 31084
rect 37200 29646 37228 31078
rect 37292 30938 37320 31146
rect 37280 30932 37332 30938
rect 37280 30874 37332 30880
rect 37280 30116 37332 30122
rect 37280 30058 37332 30064
rect 37188 29640 37240 29646
rect 37188 29582 37240 29588
rect 37186 29200 37242 29209
rect 37186 29135 37242 29144
rect 37200 28762 37228 29135
rect 37188 28756 37240 28762
rect 37188 28698 37240 28704
rect 37188 28620 37240 28626
rect 37188 28562 37240 28568
rect 37200 28257 37228 28562
rect 37186 28248 37242 28257
rect 37186 28183 37242 28192
rect 37292 27010 37320 30058
rect 37384 30002 37412 31622
rect 37476 30297 37504 32166
rect 37462 30288 37518 30297
rect 37462 30223 37518 30232
rect 37384 29974 37504 30002
rect 37370 29880 37426 29889
rect 37370 29815 37426 29824
rect 37384 29714 37412 29815
rect 37372 29708 37424 29714
rect 37372 29650 37424 29656
rect 37476 29238 37504 29974
rect 37568 29306 37596 34614
rect 37660 34542 37688 72422
rect 38384 72004 38436 72010
rect 38384 71946 38436 71952
rect 37924 71460 37976 71466
rect 37924 71402 37976 71408
rect 37936 71369 37964 71402
rect 37922 71360 37978 71369
rect 37922 71295 37978 71304
rect 38292 70916 38344 70922
rect 38292 70858 38344 70864
rect 37922 70544 37978 70553
rect 37922 70479 37978 70488
rect 37936 70446 37964 70479
rect 37924 70440 37976 70446
rect 37924 70382 37976 70388
rect 37924 69284 37976 69290
rect 37924 69226 37976 69232
rect 37936 69193 37964 69226
rect 37922 69184 37978 69193
rect 37922 69119 37978 69128
rect 37832 68128 37884 68134
rect 37832 68070 37884 68076
rect 38200 68128 38252 68134
rect 38200 68070 38252 68076
rect 37740 59560 37792 59566
rect 37740 59502 37792 59508
rect 37752 58410 37780 59502
rect 37740 58404 37792 58410
rect 37740 58346 37792 58352
rect 37752 57322 37780 58346
rect 37740 57316 37792 57322
rect 37740 57258 37792 57264
rect 37844 56302 37872 68070
rect 37924 67176 37976 67182
rect 37924 67118 37976 67124
rect 37936 66609 37964 67118
rect 37922 66600 37978 66609
rect 37922 66535 37978 66544
rect 37924 66088 37976 66094
rect 37924 66030 37976 66036
rect 37936 65385 37964 66030
rect 37922 65376 37978 65385
rect 37922 65311 37978 65320
rect 37924 65000 37976 65006
rect 37924 64942 37976 64948
rect 37936 64433 37964 64942
rect 37922 64424 37978 64433
rect 37922 64359 37978 64368
rect 37924 63912 37976 63918
rect 37924 63854 37976 63860
rect 37936 63209 37964 63854
rect 37922 63200 37978 63209
rect 37922 63135 37978 63144
rect 37924 62824 37976 62830
rect 37924 62766 37976 62772
rect 37936 62257 37964 62766
rect 38108 62688 38160 62694
rect 38108 62630 38160 62636
rect 37922 62248 37978 62257
rect 38120 62218 38148 62630
rect 37922 62183 37978 62192
rect 38108 62212 38160 62218
rect 38108 62154 38160 62160
rect 37924 61736 37976 61742
rect 37924 61678 37976 61684
rect 37936 61033 37964 61678
rect 38108 61600 38160 61606
rect 38108 61542 38160 61548
rect 38120 61334 38148 61542
rect 38108 61328 38160 61334
rect 38108 61270 38160 61276
rect 37922 61024 37978 61033
rect 37922 60959 37978 60968
rect 37924 60648 37976 60654
rect 37924 60590 37976 60596
rect 37936 59673 37964 60590
rect 38108 60512 38160 60518
rect 38108 60454 38160 60460
rect 38120 60314 38148 60454
rect 38108 60308 38160 60314
rect 38108 60250 38160 60256
rect 37922 59664 37978 59673
rect 37922 59599 37978 59608
rect 38016 59560 38068 59566
rect 38016 59502 38068 59508
rect 38028 58682 38056 59502
rect 38016 58676 38068 58682
rect 38016 58618 38068 58624
rect 38108 58336 38160 58342
rect 38108 58278 38160 58284
rect 38016 57384 38068 57390
rect 38016 57326 38068 57332
rect 37832 56296 37884 56302
rect 37832 56238 37884 56244
rect 37924 55208 37976 55214
rect 37924 55150 37976 55156
rect 37740 55140 37792 55146
rect 37740 55082 37792 55088
rect 37832 55140 37884 55146
rect 37832 55082 37884 55088
rect 37752 54058 37780 55082
rect 37844 54058 37872 55082
rect 37740 54052 37792 54058
rect 37740 53994 37792 54000
rect 37832 54052 37884 54058
rect 37832 53994 37884 54000
rect 37752 53038 37780 53994
rect 37740 53032 37792 53038
rect 37738 53000 37740 53009
rect 37792 53000 37794 53009
rect 37844 52970 37872 53994
rect 37738 52935 37794 52944
rect 37832 52964 37884 52970
rect 37752 51882 37780 52935
rect 37832 52906 37884 52912
rect 37844 51882 37872 52906
rect 37740 51876 37792 51882
rect 37740 51818 37792 51824
rect 37832 51876 37884 51882
rect 37832 51818 37884 51824
rect 37752 48890 37780 51818
rect 37740 48884 37792 48890
rect 37740 48826 37792 48832
rect 37740 48612 37792 48618
rect 37740 48554 37792 48560
rect 37752 45626 37780 48554
rect 37844 46646 37872 51818
rect 37936 49978 37964 55150
rect 38028 51066 38056 57326
rect 38120 57050 38148 58278
rect 38108 57044 38160 57050
rect 38108 56986 38160 56992
rect 38212 54738 38240 68070
rect 38200 54732 38252 54738
rect 38200 54674 38252 54680
rect 38200 54120 38252 54126
rect 38200 54062 38252 54068
rect 38108 53032 38160 53038
rect 38108 52974 38160 52980
rect 38016 51060 38068 51066
rect 38016 51002 38068 51008
rect 38120 50946 38148 52974
rect 38028 50918 38148 50946
rect 37924 49972 37976 49978
rect 37924 49914 37976 49920
rect 37924 48136 37976 48142
rect 37924 48078 37976 48084
rect 37832 46640 37884 46646
rect 37832 46582 37884 46588
rect 37936 46594 37964 48078
rect 38028 46918 38056 50918
rect 38108 50856 38160 50862
rect 38108 50798 38160 50804
rect 38120 50697 38148 50798
rect 38106 50688 38162 50697
rect 38106 50623 38162 50632
rect 38108 49768 38160 49774
rect 38108 49710 38160 49716
rect 38120 49337 38148 49710
rect 38106 49328 38162 49337
rect 38106 49263 38162 49272
rect 38212 48074 38240 54062
rect 38200 48068 38252 48074
rect 38200 48010 38252 48016
rect 38108 47456 38160 47462
rect 38108 47398 38160 47404
rect 38016 46912 38068 46918
rect 38016 46854 38068 46860
rect 37936 46566 38056 46594
rect 37924 46504 37976 46510
rect 37924 46446 37976 46452
rect 37740 45620 37792 45626
rect 37740 45562 37792 45568
rect 37752 45393 37780 45562
rect 37738 45384 37794 45393
rect 37738 45319 37794 45328
rect 37740 45280 37792 45286
rect 37738 45248 37740 45257
rect 37792 45248 37794 45257
rect 37738 45183 37794 45192
rect 37740 45076 37792 45082
rect 37740 45018 37792 45024
rect 37752 44334 37780 45018
rect 37740 44328 37792 44334
rect 37740 44270 37792 44276
rect 37752 43246 37780 44270
rect 37832 44260 37884 44266
rect 37832 44202 37884 44208
rect 37740 43240 37792 43246
rect 37740 43182 37792 43188
rect 37752 42906 37780 43182
rect 37844 43178 37872 44202
rect 37832 43172 37884 43178
rect 37832 43114 37884 43120
rect 37740 42900 37792 42906
rect 37740 42842 37792 42848
rect 37752 42294 37780 42842
rect 37844 42838 37872 43114
rect 37832 42832 37884 42838
rect 37832 42774 37884 42780
rect 37740 42288 37792 42294
rect 37740 42230 37792 42236
rect 37740 42152 37792 42158
rect 37740 42094 37792 42100
rect 37752 40066 37780 42094
rect 37832 41676 37884 41682
rect 37832 41618 37884 41624
rect 37844 40186 37872 41618
rect 37832 40180 37884 40186
rect 37832 40122 37884 40128
rect 37752 40038 37872 40066
rect 37740 39976 37792 39982
rect 37740 39918 37792 39924
rect 37752 38826 37780 39918
rect 37740 38820 37792 38826
rect 37740 38762 37792 38768
rect 37752 38457 37780 38762
rect 37738 38448 37794 38457
rect 37738 38383 37794 38392
rect 37740 37800 37792 37806
rect 37844 37788 37872 40038
rect 37936 38049 37964 46446
rect 38028 44946 38056 46566
rect 38120 45665 38148 47398
rect 38304 46170 38332 70858
rect 38292 46164 38344 46170
rect 38292 46106 38344 46112
rect 38106 45656 38162 45665
rect 38106 45591 38162 45600
rect 38292 45620 38344 45626
rect 38292 45562 38344 45568
rect 38200 45416 38252 45422
rect 38200 45358 38252 45364
rect 38016 44940 38068 44946
rect 38016 44882 38068 44888
rect 38014 44704 38070 44713
rect 38014 44639 38070 44648
rect 38028 39914 38056 44639
rect 38108 43920 38160 43926
rect 38108 43862 38160 43868
rect 38120 43217 38148 43862
rect 38106 43208 38162 43217
rect 38106 43143 38162 43152
rect 38108 43104 38160 43110
rect 38108 43046 38160 43052
rect 38120 41274 38148 43046
rect 38212 42226 38240 45358
rect 38200 42220 38252 42226
rect 38200 42162 38252 42168
rect 38200 42084 38252 42090
rect 38200 42026 38252 42032
rect 38108 41268 38160 41274
rect 38108 41210 38160 41216
rect 38108 39976 38160 39982
rect 38106 39944 38108 39953
rect 38160 39944 38162 39953
rect 38016 39908 38068 39914
rect 38106 39879 38162 39888
rect 38016 39850 38068 39856
rect 38028 39030 38056 39850
rect 38108 39092 38160 39098
rect 38108 39034 38160 39040
rect 38016 39024 38068 39030
rect 38016 38966 38068 38972
rect 38028 38554 38056 38966
rect 38120 38729 38148 39034
rect 38106 38720 38162 38729
rect 38106 38655 38162 38664
rect 38016 38548 38068 38554
rect 38016 38490 38068 38496
rect 37922 38040 37978 38049
rect 37922 37975 37978 37984
rect 37792 37760 37872 37788
rect 37740 37742 37792 37748
rect 37752 37262 37780 37742
rect 37740 37256 37792 37262
rect 37740 37198 37792 37204
rect 37752 36650 37780 37198
rect 37924 36712 37976 36718
rect 37924 36654 37976 36660
rect 37740 36644 37792 36650
rect 37740 36586 37792 36592
rect 37832 36644 37884 36650
rect 37832 36586 37884 36592
rect 37648 34536 37700 34542
rect 37648 34478 37700 34484
rect 37752 34474 37780 36586
rect 37844 34950 37872 36586
rect 37832 34944 37884 34950
rect 37832 34886 37884 34892
rect 37844 34542 37872 34886
rect 37832 34536 37884 34542
rect 37832 34478 37884 34484
rect 37740 34468 37792 34474
rect 37740 34410 37792 34416
rect 37648 32904 37700 32910
rect 37648 32846 37700 32852
rect 37556 29300 37608 29306
rect 37556 29242 37608 29248
rect 37464 29232 37516 29238
rect 37464 29174 37516 29180
rect 37464 29096 37516 29102
rect 37462 29064 37464 29073
rect 37516 29064 37518 29073
rect 37462 28999 37518 29008
rect 37370 28656 37426 28665
rect 37370 28591 37426 28600
rect 37384 28558 37412 28591
rect 37372 28552 37424 28558
rect 37372 28494 37424 28500
rect 37464 28008 37516 28014
rect 37464 27950 37516 27956
rect 37476 27849 37504 27950
rect 37462 27840 37518 27849
rect 37462 27775 37518 27784
rect 37292 26982 37412 27010
rect 37280 26920 37332 26926
rect 37278 26888 37280 26897
rect 37332 26888 37334 26897
rect 37278 26823 37334 26832
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 37292 25673 37320 25774
rect 37278 25664 37334 25673
rect 37278 25599 37334 25608
rect 37188 25356 37240 25362
rect 37188 25298 37240 25304
rect 37200 25265 37228 25298
rect 37186 25256 37242 25265
rect 37186 25191 37242 25200
rect 37186 24304 37242 24313
rect 37186 24239 37188 24248
rect 37240 24239 37242 24248
rect 37188 24210 37240 24216
rect 37384 23866 37412 26982
rect 37660 25498 37688 32846
rect 37740 32292 37792 32298
rect 37740 32234 37792 32240
rect 37832 32292 37884 32298
rect 37832 32234 37884 32240
rect 37752 31482 37780 32234
rect 37844 31958 37872 32234
rect 37832 31952 37884 31958
rect 37832 31894 37884 31900
rect 37740 31476 37792 31482
rect 37740 31418 37792 31424
rect 37752 31210 37780 31418
rect 37844 31278 37872 31894
rect 37832 31272 37884 31278
rect 37832 31214 37884 31220
rect 37740 31204 37792 31210
rect 37740 31146 37792 31152
rect 37752 30122 37780 31146
rect 37844 30190 37872 31214
rect 37832 30184 37884 30190
rect 37832 30126 37884 30132
rect 37740 30116 37792 30122
rect 37740 30058 37792 30064
rect 37740 29776 37792 29782
rect 37740 29718 37792 29724
rect 37648 25492 37700 25498
rect 37648 25434 37700 25440
rect 37556 24200 37608 24206
rect 37556 24142 37608 24148
rect 37462 23896 37518 23905
rect 37372 23860 37424 23866
rect 37462 23831 37518 23840
rect 37372 23802 37424 23808
rect 37476 23662 37504 23831
rect 37464 23656 37516 23662
rect 37464 23598 37516 23604
rect 37188 23180 37240 23186
rect 37188 23122 37240 23128
rect 37200 23089 37228 23122
rect 37186 23080 37242 23089
rect 37186 23015 37242 23024
rect 37280 22568 37332 22574
rect 37278 22536 37280 22545
rect 37332 22536 37334 22545
rect 37278 22471 37334 22480
rect 37188 22092 37240 22098
rect 37188 22034 37240 22040
rect 37200 21729 37228 22034
rect 37186 21720 37242 21729
rect 37186 21655 37242 21664
rect 37096 21616 37148 21622
rect 37096 21558 37148 21564
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 37292 21321 37320 21422
rect 37278 21312 37334 21321
rect 37278 21247 37334 21256
rect 37278 20496 37334 20505
rect 37278 20431 37334 20440
rect 37292 20398 37320 20431
rect 37280 20392 37332 20398
rect 37280 20334 37332 20340
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37292 19145 37320 19246
rect 37278 19136 37334 19145
rect 37278 19071 37334 19080
rect 37004 18964 37056 18970
rect 37004 18906 37056 18912
rect 37188 18828 37240 18834
rect 37188 18770 37240 18776
rect 37004 18760 37056 18766
rect 37200 18737 37228 18770
rect 37004 18702 37056 18708
rect 37186 18728 37242 18737
rect 36728 17332 36780 17338
rect 36728 17274 36780 17280
rect 37016 16794 37044 18702
rect 37186 18663 37242 18672
rect 37186 17912 37242 17921
rect 37186 17847 37242 17856
rect 37200 17746 37228 17847
rect 37464 17808 37516 17814
rect 37464 17750 37516 17756
rect 37188 17740 37240 17746
rect 37188 17682 37240 17688
rect 37278 17368 37334 17377
rect 37278 17303 37334 17312
rect 37096 17196 37148 17202
rect 37096 17138 37148 17144
rect 37004 16788 37056 16794
rect 37004 16730 37056 16736
rect 36912 13252 36964 13258
rect 36912 13194 36964 13200
rect 36636 12436 36688 12442
rect 36636 12378 36688 12384
rect 36268 11824 36320 11830
rect 36268 11766 36320 11772
rect 36280 4826 36308 11766
rect 36728 11756 36780 11762
rect 36728 11698 36780 11704
rect 36452 7812 36504 7818
rect 36452 7754 36504 7760
rect 36360 6180 36412 6186
rect 36360 6122 36412 6128
rect 36268 4820 36320 4826
rect 36268 4762 36320 4768
rect 36176 4752 36228 4758
rect 36176 4694 36228 4700
rect 36268 4616 36320 4622
rect 36268 4558 36320 4564
rect 36176 4480 36228 4486
rect 36176 4422 36228 4428
rect 36188 3398 36216 4422
rect 36280 4078 36308 4558
rect 36372 4146 36400 6122
rect 36464 4146 36492 7754
rect 36544 6860 36596 6866
rect 36544 6802 36596 6808
rect 36556 5370 36584 6802
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36636 5092 36688 5098
rect 36636 5034 36688 5040
rect 36544 4684 36596 4690
rect 36544 4626 36596 4632
rect 36360 4140 36412 4146
rect 36360 4082 36412 4088
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 36268 4072 36320 4078
rect 36268 4014 36320 4020
rect 36452 4004 36504 4010
rect 36452 3946 36504 3952
rect 36268 3460 36320 3466
rect 36268 3402 36320 3408
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36004 2774 36124 2802
rect 36004 800 36032 2774
rect 36280 800 36308 3402
rect 36464 2281 36492 3946
rect 36556 2825 36584 4626
rect 36648 3233 36676 5034
rect 36740 3738 36768 11698
rect 36924 6390 36952 13194
rect 37108 6458 37136 17138
rect 37292 17134 37320 17303
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37372 17060 37424 17066
rect 37372 17002 37424 17008
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 37200 16561 37228 16594
rect 37186 16552 37242 16561
rect 37186 16487 37242 16496
rect 37278 16144 37334 16153
rect 37278 16079 37334 16088
rect 37292 16046 37320 16079
rect 37280 16040 37332 16046
rect 37280 15982 37332 15988
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37200 15337 37228 15506
rect 37186 15328 37242 15337
rect 37186 15263 37242 15272
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 37292 14793 37320 14894
rect 37278 14784 37334 14793
rect 37278 14719 37334 14728
rect 37280 14612 37332 14618
rect 37280 14554 37332 14560
rect 37186 13968 37242 13977
rect 37186 13903 37242 13912
rect 37200 13870 37228 13903
rect 37188 13864 37240 13870
rect 37188 13806 37240 13812
rect 37188 13388 37240 13394
rect 37188 13330 37240 13336
rect 37200 13161 37228 13330
rect 37186 13152 37242 13161
rect 37186 13087 37242 13096
rect 37188 12300 37240 12306
rect 37188 12242 37240 12248
rect 37200 12209 37228 12242
rect 37186 12200 37242 12209
rect 37186 12135 37242 12144
rect 37186 11792 37242 11801
rect 37186 11727 37242 11736
rect 37200 11694 37228 11727
rect 37188 11688 37240 11694
rect 37188 11630 37240 11636
rect 37188 11212 37240 11218
rect 37188 11154 37240 11160
rect 37200 10985 37228 11154
rect 37186 10976 37242 10985
rect 37186 10911 37242 10920
rect 37188 10124 37240 10130
rect 37188 10066 37240 10072
rect 37200 10033 37228 10066
rect 37186 10024 37242 10033
rect 37186 9959 37242 9968
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 37200 9518 37228 9551
rect 37188 9512 37240 9518
rect 37188 9454 37240 9460
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37200 8809 37228 8978
rect 37186 8800 37242 8809
rect 37186 8735 37242 8744
rect 37186 7984 37242 7993
rect 37186 7919 37188 7928
rect 37240 7919 37242 7928
rect 37188 7890 37240 7896
rect 37186 7440 37242 7449
rect 37186 7375 37242 7384
rect 37200 7342 37228 7375
rect 37188 7336 37240 7342
rect 37188 7278 37240 7284
rect 37292 6866 37320 14554
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37280 6860 37332 6866
rect 37280 6802 37332 6808
rect 37200 6633 37228 6802
rect 37186 6624 37242 6633
rect 37186 6559 37242 6568
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 36912 6384 36964 6390
rect 36912 6326 36964 6332
rect 37004 6180 37056 6186
rect 37004 6122 37056 6128
rect 37096 6180 37148 6186
rect 37096 6122 37148 6128
rect 36912 5160 36964 5166
rect 36912 5102 36964 5108
rect 36820 4004 36872 4010
rect 36820 3946 36872 3952
rect 36728 3732 36780 3738
rect 36728 3674 36780 3680
rect 36634 3224 36690 3233
rect 36634 3159 36690 3168
rect 36728 2916 36780 2922
rect 36728 2858 36780 2864
rect 36542 2816 36598 2825
rect 36542 2751 36598 2760
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36450 2272 36506 2281
rect 36450 2207 36506 2216
rect 36556 800 36584 2450
rect 2778 504 2834 513
rect 2778 439 2834 448
rect 2962 -800 3018 800
rect 3238 -800 3294 800
rect 3606 -800 3662 800
rect 3882 -800 3938 800
rect 4158 -800 4214 800
rect 4434 -800 4490 800
rect 4710 -800 4766 800
rect 4986 -800 5042 800
rect 5354 -800 5410 800
rect 5630 -800 5686 800
rect 5906 -800 5962 800
rect 6182 -800 6238 800
rect 6458 -800 6514 800
rect 6826 -800 6882 800
rect 7102 -800 7158 800
rect 7378 -800 7434 800
rect 7654 -800 7710 800
rect 7930 -800 7986 800
rect 8206 -800 8262 800
rect 8574 -800 8630 800
rect 8850 -800 8906 800
rect 9126 -800 9182 800
rect 9402 -800 9458 800
rect 9678 -800 9734 800
rect 9954 -800 10010 800
rect 10322 -800 10378 800
rect 10598 -800 10654 800
rect 10874 -800 10930 800
rect 11150 -800 11206 800
rect 11426 -800 11482 800
rect 11794 -800 11850 800
rect 12070 -800 12126 800
rect 12346 -800 12402 800
rect 12622 -800 12678 800
rect 12898 -800 12954 800
rect 13174 -800 13230 800
rect 13542 -800 13598 800
rect 13818 -800 13874 800
rect 14094 -800 14150 800
rect 14370 -800 14426 800
rect 14646 -800 14702 800
rect 14922 -800 14978 800
rect 15290 -800 15346 800
rect 15566 -800 15622 800
rect 15842 -800 15898 800
rect 16118 -800 16174 800
rect 16394 -800 16450 800
rect 16670 -800 16726 800
rect 17038 -800 17094 800
rect 17314 -800 17370 800
rect 17590 -800 17646 800
rect 17866 -800 17922 800
rect 18142 -800 18198 800
rect 18510 -800 18566 800
rect 18786 -800 18842 800
rect 19062 -800 19118 800
rect 19338 -800 19394 800
rect 19614 -800 19670 800
rect 19890 -800 19946 800
rect 20258 -800 20314 800
rect 20534 -800 20590 800
rect 20810 -800 20866 800
rect 21086 -800 21142 800
rect 21362 -800 21418 800
rect 21638 -800 21694 800
rect 22006 -800 22062 800
rect 22282 -800 22338 800
rect 22558 -800 22614 800
rect 22834 -800 22890 800
rect 23110 -800 23166 800
rect 23478 -800 23534 800
rect 23754 -800 23810 800
rect 24030 -800 24086 800
rect 24306 -800 24362 800
rect 24582 -800 24638 800
rect 24858 -800 24914 800
rect 25226 -800 25282 800
rect 25502 -800 25558 800
rect 25778 -800 25834 800
rect 26054 -800 26110 800
rect 26330 -800 26386 800
rect 26606 -800 26662 800
rect 26974 -800 27030 800
rect 27250 -800 27306 800
rect 27526 -800 27582 800
rect 27802 -800 27858 800
rect 28078 -800 28134 800
rect 28354 -800 28410 800
rect 28722 -800 28778 800
rect 28998 -800 29054 800
rect 29274 -800 29330 800
rect 29550 -800 29606 800
rect 29826 -800 29882 800
rect 30194 -800 30250 800
rect 30470 -800 30526 800
rect 30746 -800 30802 800
rect 31022 -800 31078 800
rect 31298 -800 31354 800
rect 31574 -800 31630 800
rect 31942 -800 31998 800
rect 32218 -800 32274 800
rect 32494 -800 32550 800
rect 32770 -800 32826 800
rect 33046 -800 33102 800
rect 33322 -800 33378 800
rect 33690 -800 33746 800
rect 33966 -800 34022 800
rect 34242 -800 34298 800
rect 34518 -800 34574 800
rect 34794 -800 34850 800
rect 35162 -800 35218 800
rect 35438 -800 35494 800
rect 35714 -800 35770 800
rect 35990 -800 36046 800
rect 36266 -800 36322 800
rect 36542 -800 36598 800
rect 36740 649 36768 2858
rect 36832 1873 36860 3946
rect 36924 3942 36952 5102
rect 36912 3936 36964 3942
rect 36912 3878 36964 3884
rect 36912 3664 36964 3670
rect 36912 3606 36964 3612
rect 36818 1864 36874 1873
rect 36818 1799 36874 1808
rect 36924 800 36952 3606
rect 37016 898 37044 6122
rect 37108 4049 37136 6122
rect 37280 6112 37332 6118
rect 37280 6054 37332 6060
rect 37186 5808 37242 5817
rect 37186 5743 37188 5752
rect 37240 5743 37242 5752
rect 37188 5714 37240 5720
rect 37186 5400 37242 5409
rect 37186 5335 37242 5344
rect 37200 5166 37228 5335
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 37188 4684 37240 4690
rect 37188 4626 37240 4632
rect 37200 4457 37228 4626
rect 37186 4448 37242 4457
rect 37186 4383 37242 4392
rect 37094 4040 37150 4049
rect 37094 3975 37150 3984
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 37200 1057 37228 3538
rect 37292 3058 37320 6054
rect 37384 5302 37412 17002
rect 37372 5296 37424 5302
rect 37372 5238 37424 5244
rect 37476 4758 37504 17750
rect 37568 9654 37596 24142
rect 37752 22778 37780 29718
rect 37936 29306 37964 36654
rect 38108 34400 38160 34406
rect 38108 34342 38160 34348
rect 38016 33448 38068 33454
rect 38016 33390 38068 33396
rect 38028 32473 38056 33390
rect 38120 33153 38148 34342
rect 38212 33658 38240 42026
rect 38304 40050 38332 45562
rect 38292 40044 38344 40050
rect 38292 39986 38344 39992
rect 38292 37800 38344 37806
rect 38292 37742 38344 37748
rect 38200 33652 38252 33658
rect 38200 33594 38252 33600
rect 38106 33144 38162 33153
rect 38106 33079 38162 33088
rect 38014 32464 38070 32473
rect 38014 32399 38070 32408
rect 38016 31272 38068 31278
rect 38016 31214 38068 31220
rect 37924 29300 37976 29306
rect 37924 29242 37976 29248
rect 37830 28928 37886 28937
rect 37830 28863 37886 28872
rect 37844 27130 37872 28863
rect 37924 28008 37976 28014
rect 37924 27950 37976 27956
rect 37936 27305 37964 27950
rect 37922 27296 37978 27305
rect 37922 27231 37978 27240
rect 37832 27124 37884 27130
rect 37832 27066 37884 27072
rect 37924 26920 37976 26926
rect 37924 26862 37976 26868
rect 37936 26489 37964 26862
rect 37922 26480 37978 26489
rect 37922 26415 37978 26424
rect 37922 26072 37978 26081
rect 37922 26007 37978 26016
rect 37936 25838 37964 26007
rect 37924 25832 37976 25838
rect 37924 25774 37976 25780
rect 37924 24744 37976 24750
rect 37922 24712 37924 24721
rect 37976 24712 37978 24721
rect 37922 24647 37978 24656
rect 38028 22778 38056 31214
rect 38200 30184 38252 30190
rect 38200 30126 38252 30132
rect 38108 29096 38160 29102
rect 38108 29038 38160 29044
rect 38120 28665 38148 29038
rect 38106 28656 38162 28665
rect 38106 28591 38162 28600
rect 38108 23656 38160 23662
rect 38108 23598 38160 23604
rect 38120 23497 38148 23598
rect 38106 23488 38162 23497
rect 38106 23423 38162 23432
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 38016 22772 38068 22778
rect 38016 22714 38068 22720
rect 37924 22568 37976 22574
rect 37924 22510 37976 22516
rect 37936 22137 37964 22510
rect 37922 22128 37978 22137
rect 37922 22063 37978 22072
rect 37924 21480 37976 21486
rect 37924 21422 37976 21428
rect 37936 20913 37964 21422
rect 37922 20904 37978 20913
rect 37922 20839 37978 20848
rect 37924 20392 37976 20398
rect 37924 20334 37976 20340
rect 37936 19961 37964 20334
rect 37922 19952 37978 19961
rect 37922 19887 37978 19896
rect 37922 19544 37978 19553
rect 37922 19479 37978 19488
rect 37936 19310 37964 19479
rect 37924 19304 37976 19310
rect 37924 19246 37976 19252
rect 37648 18692 37700 18698
rect 37648 18634 37700 18640
rect 37556 9648 37608 9654
rect 37556 9590 37608 9596
rect 37556 9104 37608 9110
rect 37556 9046 37608 9052
rect 37464 4752 37516 4758
rect 37464 4694 37516 4700
rect 37568 4146 37596 9046
rect 37660 7546 37688 18634
rect 38212 18426 38240 30126
rect 38304 29850 38332 37742
rect 38396 32434 38424 71946
rect 38844 68672 38896 68678
rect 38844 68614 38896 68620
rect 38752 67312 38804 67318
rect 38752 67254 38804 67260
rect 38660 67040 38712 67046
rect 38660 66982 38712 66988
rect 38568 66224 38620 66230
rect 38568 66166 38620 66172
rect 38476 63232 38528 63238
rect 38476 63174 38528 63180
rect 38488 44198 38516 63174
rect 38580 49842 38608 66166
rect 38672 50386 38700 66982
rect 38764 50930 38792 67254
rect 38856 66042 38884 68614
rect 38936 67652 38988 67658
rect 38936 67594 38988 67600
rect 38948 67425 38976 67594
rect 38934 67416 38990 67425
rect 38934 67351 38990 67360
rect 38856 66014 38976 66042
rect 38844 65952 38896 65958
rect 38844 65894 38896 65900
rect 38752 50924 38804 50930
rect 38752 50866 38804 50872
rect 38660 50380 38712 50386
rect 38660 50322 38712 50328
rect 38568 49836 38620 49842
rect 38568 49778 38620 49784
rect 38856 48686 38884 65894
rect 38948 55962 38976 66014
rect 38936 55956 38988 55962
rect 38936 55898 38988 55904
rect 38936 54596 38988 54602
rect 38936 54538 38988 54544
rect 38844 48680 38896 48686
rect 38844 48622 38896 48628
rect 38568 48204 38620 48210
rect 38568 48146 38620 48152
rect 38476 44192 38528 44198
rect 38476 44134 38528 44140
rect 38476 42220 38528 42226
rect 38476 42162 38528 42168
rect 38488 37874 38516 42162
rect 38580 40526 38608 48146
rect 38660 46164 38712 46170
rect 38660 46106 38712 46112
rect 38568 40520 38620 40526
rect 38568 40462 38620 40468
rect 38568 40180 38620 40186
rect 38568 40122 38620 40128
rect 38580 38321 38608 40122
rect 38566 38312 38622 38321
rect 38566 38247 38622 38256
rect 38476 37868 38528 37874
rect 38476 37810 38528 37816
rect 38476 37324 38528 37330
rect 38476 37266 38528 37272
rect 38384 32428 38436 32434
rect 38384 32370 38436 32376
rect 38292 29844 38344 29850
rect 38292 29786 38344 29792
rect 38488 28218 38516 37266
rect 38568 34536 38620 34542
rect 38568 34478 38620 34484
rect 38476 28212 38528 28218
rect 38476 28154 38528 28160
rect 38580 24614 38608 34478
rect 38672 31414 38700 46106
rect 38752 44328 38804 44334
rect 38752 44270 38804 44276
rect 38764 37194 38792 44270
rect 38844 41064 38896 41070
rect 38844 41006 38896 41012
rect 38752 37188 38804 37194
rect 38752 37130 38804 37136
rect 38752 35488 38804 35494
rect 38752 35430 38804 35436
rect 38660 31408 38712 31414
rect 38660 31350 38712 31356
rect 38764 29510 38792 35430
rect 38856 31822 38884 41006
rect 38948 36378 38976 54538
rect 39040 54194 39068 80310
rect 39120 71528 39172 71534
rect 39120 71470 39172 71476
rect 39028 54188 39080 54194
rect 39028 54130 39080 54136
rect 39028 51944 39080 51950
rect 39028 51886 39080 51892
rect 39040 43654 39068 51886
rect 39028 43648 39080 43654
rect 39028 43590 39080 43596
rect 39028 43240 39080 43246
rect 39028 43182 39080 43188
rect 38936 36372 38988 36378
rect 38936 36314 38988 36320
rect 39040 33590 39068 43182
rect 39028 33584 39080 33590
rect 39028 33526 39080 33532
rect 38936 32360 38988 32366
rect 38936 32302 38988 32308
rect 38844 31816 38896 31822
rect 38844 31758 38896 31764
rect 38752 29504 38804 29510
rect 38752 29446 38804 29452
rect 38568 24608 38620 24614
rect 38568 24550 38620 24556
rect 38948 23866 38976 32302
rect 39132 31346 39160 71470
rect 39224 60042 39252 82486
rect 39396 81252 39448 81258
rect 39396 81194 39448 81200
rect 39304 81184 39356 81190
rect 39304 81126 39356 81132
rect 39212 60036 39264 60042
rect 39212 59978 39264 59984
rect 39212 57316 39264 57322
rect 39212 57258 39264 57264
rect 39224 46986 39252 57258
rect 39316 55214 39344 81126
rect 39408 57458 39436 81194
rect 39488 71460 39540 71466
rect 39488 71402 39540 71408
rect 39396 57452 39448 57458
rect 39396 57394 39448 57400
rect 39396 56160 39448 56166
rect 39396 56102 39448 56108
rect 39304 55208 39356 55214
rect 39304 55150 39356 55156
rect 39212 46980 39264 46986
rect 39212 46922 39264 46928
rect 39408 45422 39436 56102
rect 39396 45416 39448 45422
rect 39396 45358 39448 45364
rect 39500 32502 39528 71402
rect 39580 65408 39632 65414
rect 39580 65350 39632 65356
rect 39592 49298 39620 65350
rect 39580 49292 39632 49298
rect 39580 49234 39632 49240
rect 39488 32496 39540 32502
rect 39488 32438 39540 32444
rect 39120 31340 39172 31346
rect 39120 31282 39172 31288
rect 38936 23860 38988 23866
rect 38936 23802 38988 23808
rect 38200 18420 38252 18426
rect 38200 18362 38252 18368
rect 37922 18320 37978 18329
rect 37922 18255 37978 18264
rect 37936 18222 37964 18255
rect 37924 18216 37976 18222
rect 37924 18158 37976 18164
rect 37924 17128 37976 17134
rect 37924 17070 37976 17076
rect 37936 16969 37964 17070
rect 37922 16960 37978 16969
rect 37922 16895 37978 16904
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 37740 10532 37792 10538
rect 37740 10474 37792 10480
rect 37648 7540 37700 7546
rect 37648 7482 37700 7488
rect 37752 5370 37780 10474
rect 37844 9654 37872 16050
rect 37924 16040 37976 16046
rect 37924 15982 37976 15988
rect 37936 15745 37964 15982
rect 37922 15736 37978 15745
rect 37922 15671 37978 15680
rect 37924 14952 37976 14958
rect 37924 14894 37976 14900
rect 37936 14385 37964 14894
rect 38016 14544 38068 14550
rect 38016 14486 38068 14492
rect 37922 14376 37978 14385
rect 37922 14311 37978 14320
rect 37924 13864 37976 13870
rect 37924 13806 37976 13812
rect 37936 13569 37964 13806
rect 37922 13560 37978 13569
rect 37922 13495 37978 13504
rect 37922 12744 37978 12753
rect 37922 12679 37924 12688
rect 37976 12679 37978 12688
rect 37924 12650 37976 12656
rect 37924 11620 37976 11626
rect 37924 11562 37976 11568
rect 37936 11393 37964 11562
rect 37922 11384 37978 11393
rect 37922 11319 37978 11328
rect 37922 10568 37978 10577
rect 37922 10503 37924 10512
rect 37976 10503 37978 10512
rect 37924 10474 37976 10480
rect 37832 9648 37884 9654
rect 37832 9590 37884 9596
rect 37924 9444 37976 9450
rect 37924 9386 37976 9392
rect 37936 9217 37964 9386
rect 37922 9208 37978 9217
rect 37922 9143 37978 9152
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37740 5364 37792 5370
rect 37740 5306 37792 5312
rect 37844 4146 37872 8910
rect 37922 8392 37978 8401
rect 37922 8327 37924 8336
rect 37976 8327 37978 8336
rect 37924 8298 37976 8304
rect 37924 7268 37976 7274
rect 37924 7210 37976 7216
rect 37936 7041 37964 7210
rect 37922 7032 37978 7041
rect 37922 6967 37978 6976
rect 37922 6216 37978 6225
rect 37922 6151 37924 6160
rect 37976 6151 37978 6160
rect 37924 6122 37976 6128
rect 37924 5092 37976 5098
rect 37924 5034 37976 5040
rect 37936 4865 37964 5034
rect 37922 4856 37978 4865
rect 37922 4791 37978 4800
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37186 1048 37242 1057
rect 37186 983 37242 992
rect 37016 870 37228 898
rect 37200 800 37228 870
rect 37476 800 37504 3878
rect 38028 3194 38056 14486
rect 38936 5024 38988 5030
rect 38936 4966 38988 4972
rect 38108 4004 38160 4010
rect 38108 3946 38160 3952
rect 37832 3188 37884 3194
rect 37832 3130 37884 3136
rect 38016 3188 38068 3194
rect 38016 3130 38068 3136
rect 37740 2984 37792 2990
rect 37740 2926 37792 2932
rect 37752 800 37780 2926
rect 37844 2854 37872 3130
rect 38016 3052 38068 3058
rect 38016 2994 38068 3000
rect 37924 2916 37976 2922
rect 37924 2858 37976 2864
rect 37832 2848 37884 2854
rect 37832 2790 37884 2796
rect 36726 640 36782 649
rect 36726 575 36782 584
rect 36910 -800 36966 800
rect 37186 -800 37242 800
rect 37462 -800 37518 800
rect 37738 -800 37794 800
rect 37936 241 37964 2858
rect 38028 800 38056 2994
rect 38120 1465 38148 3946
rect 38660 3392 38712 3398
rect 38660 3334 38712 3340
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 38106 1456 38162 1465
rect 38106 1391 38162 1400
rect 38304 800 38332 2450
rect 38672 800 38700 3334
rect 38948 800 38976 4966
rect 39488 4072 39540 4078
rect 39488 4014 39540 4020
rect 39212 3528 39264 3534
rect 39212 3470 39264 3476
rect 39224 800 39252 3470
rect 39500 800 39528 4014
rect 39764 2848 39816 2854
rect 39764 2790 39816 2796
rect 39776 800 39804 2790
rect 37922 232 37978 241
rect 37922 167 37978 176
rect 38014 -800 38070 800
rect 38290 -800 38346 800
rect 38658 -800 38714 800
rect 38934 -800 38990 800
rect 39210 -800 39266 800
rect 39486 -800 39542 800
rect 39762 -800 39818 800
<< via2 >>
rect 3330 119448 3386 119504
rect 1398 116184 1454 116240
rect 1950 115404 1952 115424
rect 1952 115404 2004 115424
rect 2004 115404 2006 115424
rect 1950 115368 2006 115404
rect 2042 114552 2098 114608
rect 1950 113772 1952 113792
rect 1952 113772 2004 113792
rect 2004 113772 2006 113792
rect 1950 113736 2006 113772
rect 1398 111308 1454 111344
rect 1398 111288 1400 111308
rect 1400 111288 1452 111308
rect 1452 111288 1454 111308
rect 1858 112920 1914 112976
rect 1950 112140 1952 112160
rect 1952 112140 2004 112160
rect 2004 112140 2006 112160
rect 1950 112104 2006 112140
rect 1950 110508 1952 110528
rect 1952 110508 2004 110528
rect 2004 110508 2006 110528
rect 1950 110472 2006 110508
rect 2042 109556 2044 109576
rect 2044 109556 2096 109576
rect 2096 109556 2098 109576
rect 2042 109520 2098 109556
rect 1950 108724 2006 108760
rect 1950 108704 1952 108724
rect 1952 108704 2004 108724
rect 2004 108704 2006 108724
rect 2042 107908 2098 107944
rect 2042 107888 2044 107908
rect 2044 107888 2096 107908
rect 2096 107888 2098 107908
rect 1950 107092 2006 107128
rect 1950 107072 1952 107092
rect 1952 107072 2004 107092
rect 2004 107072 2006 107092
rect 1766 106292 1768 106312
rect 1768 106292 1820 106312
rect 1820 106292 1822 106312
rect 1766 106256 1822 106292
rect 1398 105440 1454 105496
rect 1858 104624 1914 104680
rect 1858 103808 1914 103864
rect 1858 103012 1914 103048
rect 1858 102992 1860 103012
rect 1860 102992 1912 103012
rect 1912 102992 1914 103012
rect 1858 102176 1914 102232
rect 1858 101360 1914 101416
rect 1858 100544 1914 100600
rect 1858 99592 1914 99648
rect 1858 98776 1914 98832
rect 1858 97960 1914 98016
rect 1858 97164 1914 97200
rect 1858 97144 1860 97164
rect 1860 97144 1912 97164
rect 1912 97144 1914 97164
rect 1858 96328 1914 96384
rect 1858 95512 1914 95568
rect 1858 94696 1914 94752
rect 1858 93900 1914 93936
rect 1858 93880 1860 93900
rect 1860 93880 1912 93900
rect 1912 93880 1914 93900
rect 2962 117816 3018 117872
rect 2870 117000 2926 117056
rect 3146 118632 3202 118688
rect 36358 119584 36414 119640
rect 4220 117530 4276 117532
rect 4300 117530 4356 117532
rect 4380 117530 4436 117532
rect 4460 117530 4516 117532
rect 4220 117478 4246 117530
rect 4246 117478 4276 117530
rect 4300 117478 4310 117530
rect 4310 117478 4356 117530
rect 4380 117478 4426 117530
rect 4426 117478 4436 117530
rect 4460 117478 4490 117530
rect 4490 117478 4516 117530
rect 4220 117476 4276 117478
rect 4300 117476 4356 117478
rect 4380 117476 4436 117478
rect 4460 117476 4516 117478
rect 4220 116442 4276 116444
rect 4300 116442 4356 116444
rect 4380 116442 4436 116444
rect 4460 116442 4516 116444
rect 4220 116390 4246 116442
rect 4246 116390 4276 116442
rect 4300 116390 4310 116442
rect 4310 116390 4356 116442
rect 4380 116390 4426 116442
rect 4426 116390 4436 116442
rect 4460 116390 4490 116442
rect 4490 116390 4516 116442
rect 4220 116388 4276 116390
rect 4300 116388 4356 116390
rect 4380 116388 4436 116390
rect 4460 116388 4516 116390
rect 4220 115354 4276 115356
rect 4300 115354 4356 115356
rect 4380 115354 4436 115356
rect 4460 115354 4516 115356
rect 4220 115302 4246 115354
rect 4246 115302 4276 115354
rect 4300 115302 4310 115354
rect 4310 115302 4356 115354
rect 4380 115302 4426 115354
rect 4426 115302 4436 115354
rect 4460 115302 4490 115354
rect 4490 115302 4516 115354
rect 4220 115300 4276 115302
rect 4300 115300 4356 115302
rect 4380 115300 4436 115302
rect 4460 115300 4516 115302
rect 1858 93064 1914 93120
rect 1858 92248 1914 92304
rect 1858 91432 1914 91488
rect 1858 90636 1914 90672
rect 1858 90616 1860 90636
rect 1860 90616 1912 90636
rect 1912 90616 1914 90636
rect 1858 89664 1914 89720
rect 1858 88868 1914 88904
rect 1858 88848 1860 88868
rect 1860 88848 1912 88868
rect 1912 88848 1914 88868
rect 1858 88032 1914 88088
rect 1858 87216 1914 87272
rect 1858 86400 1914 86456
rect 1858 85620 1860 85640
rect 1860 85620 1912 85640
rect 1912 85620 1914 85640
rect 1858 85584 1914 85620
rect 1858 84768 1914 84824
rect 1858 83952 1914 84008
rect 1398 83136 1454 83192
rect 1858 82340 1914 82376
rect 1858 82320 1860 82340
rect 1860 82320 1912 82340
rect 1912 82320 1914 82340
rect 1858 81504 1914 81560
rect 1398 80688 1454 80744
rect 1398 79756 1454 79792
rect 1398 79736 1400 79756
rect 1400 79736 1452 79756
rect 1452 79736 1454 79756
rect 1858 78920 1914 78976
rect 1858 78104 1914 78160
rect 1398 77288 1454 77344
rect 1398 76492 1454 76528
rect 1398 76472 1400 76492
rect 1400 76472 1452 76492
rect 1452 76472 1454 76492
rect 1858 75656 1914 75712
rect 1858 74840 1914 74896
rect 1858 74024 1914 74080
rect 1858 73228 1914 73264
rect 1858 73208 1860 73228
rect 1860 73208 1912 73228
rect 1912 73208 1914 73228
rect 1858 72392 1914 72448
rect 1858 71576 1914 71632
rect 1858 70760 1914 70816
rect 1858 69808 1914 69864
rect 1858 68992 1914 69048
rect 1858 68212 1860 68232
rect 1860 68212 1912 68232
rect 1912 68212 1914 68232
rect 1858 68176 1914 68212
rect 1398 67360 1454 67416
rect 1398 66544 1454 66600
rect 1398 65728 1454 65784
rect 1398 64948 1400 64968
rect 1400 64948 1452 64968
rect 1452 64948 1454 64968
rect 1398 64912 1454 64948
rect 1398 64096 1454 64152
rect 1398 63280 1454 63336
rect 1398 62464 1454 62520
rect 1398 61684 1400 61704
rect 1400 61684 1452 61704
rect 1452 61684 1454 61704
rect 1398 61648 1454 61684
rect 1398 60832 1454 60888
rect 1398 59880 1454 59936
rect 1398 59084 1454 59120
rect 1398 59064 1400 59084
rect 1400 59064 1452 59084
rect 1452 59064 1454 59084
rect 1398 58248 1454 58304
rect 1398 57432 1454 57488
rect 1398 56616 1454 56672
rect 1398 55820 1454 55856
rect 1398 55800 1400 55820
rect 1400 55800 1452 55820
rect 1452 55800 1454 55820
rect 1398 54984 1454 55040
rect 1398 54168 1454 54224
rect 1398 53352 1454 53408
rect 1398 47540 1400 47560
rect 1400 47540 1452 47560
rect 1452 47540 1454 47560
rect 1398 47504 1454 47540
rect 1398 46688 1454 46744
rect 1858 52556 1914 52592
rect 1858 52536 1860 52556
rect 1860 52536 1912 52556
rect 1912 52536 1914 52556
rect 1858 51720 1914 51776
rect 1858 50904 1914 50960
rect 1858 49952 1914 50008
rect 1858 49136 1914 49192
rect 1858 48320 1914 48376
rect 1858 45872 1914 45928
rect 1858 45056 1914 45112
rect 1858 44276 1860 44296
rect 1860 44276 1912 44296
rect 1912 44276 1914 44296
rect 1858 44240 1914 44276
rect 1858 43424 1914 43480
rect 1858 42608 1914 42664
rect 1858 41792 1914 41848
rect 1858 41012 1860 41032
rect 1860 41012 1912 41032
rect 1912 41012 1914 41032
rect 1858 40976 1914 41012
rect 1858 40024 1914 40080
rect 1858 39208 1914 39264
rect 1858 38428 1860 38448
rect 1860 38428 1912 38448
rect 1912 38428 1914 38448
rect 1858 38392 1914 38428
rect 1398 36760 1454 36816
rect 1858 37576 1914 37632
rect 1398 35944 1454 36000
rect 1398 35148 1454 35184
rect 1398 35128 1400 35148
rect 1400 35128 1452 35148
rect 1452 35128 1454 35148
rect 1398 34312 1454 34368
rect 1858 33496 1914 33552
rect 1398 32680 1454 32736
rect 1398 31884 1454 31920
rect 1398 31864 1400 31884
rect 1400 31864 1452 31884
rect 1452 31864 1454 31884
rect 1398 31048 1454 31104
rect 1398 30132 1400 30152
rect 1400 30132 1452 30152
rect 1452 30132 1454 30152
rect 1398 30096 1454 30132
rect 1398 29280 1454 29336
rect 1398 28500 1400 28520
rect 1400 28500 1452 28520
rect 1452 28500 1454 28520
rect 1398 28464 1454 28500
rect 1858 27648 1914 27704
rect 1858 26852 1914 26888
rect 1858 26832 1860 26852
rect 1860 26832 1912 26852
rect 1912 26832 1914 26852
rect 1858 26016 1914 26072
rect 1858 25200 1914 25256
rect 1398 22752 1454 22808
rect 1858 24384 1914 24440
rect 1398 21936 1454 21992
rect 1858 23604 1860 23624
rect 1860 23604 1912 23624
rect 1912 23604 1914 23624
rect 1858 23568 1914 23604
rect 1398 21120 1454 21176
rect 1398 20168 1454 20224
rect 1398 19352 1454 19408
rect 1398 18536 1454 18592
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 16904 1454 16960
rect 1398 16088 1454 16144
rect 1398 15272 1454 15328
rect 1398 14476 1454 14512
rect 1398 14456 1400 14476
rect 1400 14456 1452 14476
rect 1452 14456 1454 14476
rect 1398 13640 1454 13696
rect 1398 12824 1454 12880
rect 1398 12008 1454 12064
rect 1398 11212 1454 11248
rect 1398 11192 1400 11212
rect 1400 11192 1452 11212
rect 1452 11192 1454 11212
rect 1398 10240 1454 10296
rect 1398 9460 1400 9480
rect 1400 9460 1452 9480
rect 1452 9460 1454 9480
rect 1398 9424 1454 9460
rect 1398 8608 1454 8664
rect 1398 7792 1454 7848
rect 1398 6976 1454 7032
rect 1398 6196 1400 6216
rect 1400 6196 1452 6216
rect 1452 6196 1454 6216
rect 1398 6160 1454 6196
rect 2042 5344 2098 5400
rect 1398 4528 1454 4584
rect 1306 2896 1362 2952
rect 2778 3712 2834 3768
rect 4220 114266 4276 114268
rect 4300 114266 4356 114268
rect 4380 114266 4436 114268
rect 4460 114266 4516 114268
rect 4220 114214 4246 114266
rect 4246 114214 4276 114266
rect 4300 114214 4310 114266
rect 4310 114214 4356 114266
rect 4380 114214 4426 114266
rect 4426 114214 4436 114266
rect 4460 114214 4490 114266
rect 4490 114214 4516 114266
rect 4220 114212 4276 114214
rect 4300 114212 4356 114214
rect 4380 114212 4436 114214
rect 4460 114212 4516 114214
rect 4220 113178 4276 113180
rect 4300 113178 4356 113180
rect 4380 113178 4436 113180
rect 4460 113178 4516 113180
rect 4220 113126 4246 113178
rect 4246 113126 4276 113178
rect 4300 113126 4310 113178
rect 4310 113126 4356 113178
rect 4380 113126 4426 113178
rect 4426 113126 4436 113178
rect 4460 113126 4490 113178
rect 4490 113126 4516 113178
rect 4220 113124 4276 113126
rect 4300 113124 4356 113126
rect 4380 113124 4436 113126
rect 4460 113124 4516 113126
rect 4220 112090 4276 112092
rect 4300 112090 4356 112092
rect 4380 112090 4436 112092
rect 4460 112090 4516 112092
rect 4220 112038 4246 112090
rect 4246 112038 4276 112090
rect 4300 112038 4310 112090
rect 4310 112038 4356 112090
rect 4380 112038 4426 112090
rect 4426 112038 4436 112090
rect 4460 112038 4490 112090
rect 4490 112038 4516 112090
rect 4220 112036 4276 112038
rect 4300 112036 4356 112038
rect 4380 112036 4436 112038
rect 4460 112036 4516 112038
rect 4220 111002 4276 111004
rect 4300 111002 4356 111004
rect 4380 111002 4436 111004
rect 4460 111002 4516 111004
rect 4220 110950 4246 111002
rect 4246 110950 4276 111002
rect 4300 110950 4310 111002
rect 4310 110950 4356 111002
rect 4380 110950 4426 111002
rect 4426 110950 4436 111002
rect 4460 110950 4490 111002
rect 4490 110950 4516 111002
rect 4220 110948 4276 110950
rect 4300 110948 4356 110950
rect 4380 110948 4436 110950
rect 4460 110948 4516 110950
rect 4220 109914 4276 109916
rect 4300 109914 4356 109916
rect 4380 109914 4436 109916
rect 4460 109914 4516 109916
rect 4220 109862 4246 109914
rect 4246 109862 4276 109914
rect 4300 109862 4310 109914
rect 4310 109862 4356 109914
rect 4380 109862 4426 109914
rect 4426 109862 4436 109914
rect 4460 109862 4490 109914
rect 4490 109862 4516 109914
rect 4220 109860 4276 109862
rect 4300 109860 4356 109862
rect 4380 109860 4436 109862
rect 4460 109860 4516 109862
rect 4220 108826 4276 108828
rect 4300 108826 4356 108828
rect 4380 108826 4436 108828
rect 4460 108826 4516 108828
rect 4220 108774 4246 108826
rect 4246 108774 4276 108826
rect 4300 108774 4310 108826
rect 4310 108774 4356 108826
rect 4380 108774 4426 108826
rect 4426 108774 4436 108826
rect 4460 108774 4490 108826
rect 4490 108774 4516 108826
rect 4220 108772 4276 108774
rect 4300 108772 4356 108774
rect 4380 108772 4436 108774
rect 4460 108772 4516 108774
rect 4220 107738 4276 107740
rect 4300 107738 4356 107740
rect 4380 107738 4436 107740
rect 4460 107738 4516 107740
rect 4220 107686 4246 107738
rect 4246 107686 4276 107738
rect 4300 107686 4310 107738
rect 4310 107686 4356 107738
rect 4380 107686 4426 107738
rect 4426 107686 4436 107738
rect 4460 107686 4490 107738
rect 4490 107686 4516 107738
rect 4220 107684 4276 107686
rect 4300 107684 4356 107686
rect 4380 107684 4436 107686
rect 4460 107684 4516 107686
rect 4220 106650 4276 106652
rect 4300 106650 4356 106652
rect 4380 106650 4436 106652
rect 4460 106650 4516 106652
rect 4220 106598 4246 106650
rect 4246 106598 4276 106650
rect 4300 106598 4310 106650
rect 4310 106598 4356 106650
rect 4380 106598 4426 106650
rect 4426 106598 4436 106650
rect 4460 106598 4490 106650
rect 4490 106598 4516 106650
rect 4220 106596 4276 106598
rect 4300 106596 4356 106598
rect 4380 106596 4436 106598
rect 4460 106596 4516 106598
rect 4220 105562 4276 105564
rect 4300 105562 4356 105564
rect 4380 105562 4436 105564
rect 4460 105562 4516 105564
rect 4220 105510 4246 105562
rect 4246 105510 4276 105562
rect 4300 105510 4310 105562
rect 4310 105510 4356 105562
rect 4380 105510 4426 105562
rect 4426 105510 4436 105562
rect 4460 105510 4490 105562
rect 4490 105510 4516 105562
rect 4220 105508 4276 105510
rect 4300 105508 4356 105510
rect 4380 105508 4436 105510
rect 4460 105508 4516 105510
rect 4220 104474 4276 104476
rect 4300 104474 4356 104476
rect 4380 104474 4436 104476
rect 4460 104474 4516 104476
rect 4220 104422 4246 104474
rect 4246 104422 4276 104474
rect 4300 104422 4310 104474
rect 4310 104422 4356 104474
rect 4380 104422 4426 104474
rect 4426 104422 4436 104474
rect 4460 104422 4490 104474
rect 4490 104422 4516 104474
rect 4220 104420 4276 104422
rect 4300 104420 4356 104422
rect 4380 104420 4436 104422
rect 4460 104420 4516 104422
rect 4220 103386 4276 103388
rect 4300 103386 4356 103388
rect 4380 103386 4436 103388
rect 4460 103386 4516 103388
rect 4220 103334 4246 103386
rect 4246 103334 4276 103386
rect 4300 103334 4310 103386
rect 4310 103334 4356 103386
rect 4380 103334 4426 103386
rect 4426 103334 4436 103386
rect 4460 103334 4490 103386
rect 4490 103334 4516 103386
rect 4220 103332 4276 103334
rect 4300 103332 4356 103334
rect 4380 103332 4436 103334
rect 4460 103332 4516 103334
rect 4220 102298 4276 102300
rect 4300 102298 4356 102300
rect 4380 102298 4436 102300
rect 4460 102298 4516 102300
rect 4220 102246 4246 102298
rect 4246 102246 4276 102298
rect 4300 102246 4310 102298
rect 4310 102246 4356 102298
rect 4380 102246 4426 102298
rect 4426 102246 4436 102298
rect 4460 102246 4490 102298
rect 4490 102246 4516 102298
rect 4220 102244 4276 102246
rect 4300 102244 4356 102246
rect 4380 102244 4436 102246
rect 4460 102244 4516 102246
rect 4220 101210 4276 101212
rect 4300 101210 4356 101212
rect 4380 101210 4436 101212
rect 4460 101210 4516 101212
rect 4220 101158 4246 101210
rect 4246 101158 4276 101210
rect 4300 101158 4310 101210
rect 4310 101158 4356 101210
rect 4380 101158 4426 101210
rect 4426 101158 4436 101210
rect 4460 101158 4490 101210
rect 4490 101158 4516 101210
rect 4220 101156 4276 101158
rect 4300 101156 4356 101158
rect 4380 101156 4436 101158
rect 4460 101156 4516 101158
rect 4220 100122 4276 100124
rect 4300 100122 4356 100124
rect 4380 100122 4436 100124
rect 4460 100122 4516 100124
rect 4220 100070 4246 100122
rect 4246 100070 4276 100122
rect 4300 100070 4310 100122
rect 4310 100070 4356 100122
rect 4380 100070 4426 100122
rect 4426 100070 4436 100122
rect 4460 100070 4490 100122
rect 4490 100070 4516 100122
rect 4220 100068 4276 100070
rect 4300 100068 4356 100070
rect 4380 100068 4436 100070
rect 4460 100068 4516 100070
rect 4220 99034 4276 99036
rect 4300 99034 4356 99036
rect 4380 99034 4436 99036
rect 4460 99034 4516 99036
rect 4220 98982 4246 99034
rect 4246 98982 4276 99034
rect 4300 98982 4310 99034
rect 4310 98982 4356 99034
rect 4380 98982 4426 99034
rect 4426 98982 4436 99034
rect 4460 98982 4490 99034
rect 4490 98982 4516 99034
rect 4220 98980 4276 98982
rect 4300 98980 4356 98982
rect 4380 98980 4436 98982
rect 4460 98980 4516 98982
rect 4220 97946 4276 97948
rect 4300 97946 4356 97948
rect 4380 97946 4436 97948
rect 4460 97946 4516 97948
rect 4220 97894 4246 97946
rect 4246 97894 4276 97946
rect 4300 97894 4310 97946
rect 4310 97894 4356 97946
rect 4380 97894 4426 97946
rect 4426 97894 4436 97946
rect 4460 97894 4490 97946
rect 4490 97894 4516 97946
rect 4220 97892 4276 97894
rect 4300 97892 4356 97894
rect 4380 97892 4436 97894
rect 4460 97892 4516 97894
rect 4220 96858 4276 96860
rect 4300 96858 4356 96860
rect 4380 96858 4436 96860
rect 4460 96858 4516 96860
rect 4220 96806 4246 96858
rect 4246 96806 4276 96858
rect 4300 96806 4310 96858
rect 4310 96806 4356 96858
rect 4380 96806 4426 96858
rect 4426 96806 4436 96858
rect 4460 96806 4490 96858
rect 4490 96806 4516 96858
rect 4220 96804 4276 96806
rect 4300 96804 4356 96806
rect 4380 96804 4436 96806
rect 4460 96804 4516 96806
rect 4220 95770 4276 95772
rect 4300 95770 4356 95772
rect 4380 95770 4436 95772
rect 4460 95770 4516 95772
rect 4220 95718 4246 95770
rect 4246 95718 4276 95770
rect 4300 95718 4310 95770
rect 4310 95718 4356 95770
rect 4380 95718 4426 95770
rect 4426 95718 4436 95770
rect 4460 95718 4490 95770
rect 4490 95718 4516 95770
rect 4220 95716 4276 95718
rect 4300 95716 4356 95718
rect 4380 95716 4436 95718
rect 4460 95716 4516 95718
rect 4220 94682 4276 94684
rect 4300 94682 4356 94684
rect 4380 94682 4436 94684
rect 4460 94682 4516 94684
rect 4220 94630 4246 94682
rect 4246 94630 4276 94682
rect 4300 94630 4310 94682
rect 4310 94630 4356 94682
rect 4380 94630 4426 94682
rect 4426 94630 4436 94682
rect 4460 94630 4490 94682
rect 4490 94630 4516 94682
rect 4220 94628 4276 94630
rect 4300 94628 4356 94630
rect 4380 94628 4436 94630
rect 4460 94628 4516 94630
rect 4220 93594 4276 93596
rect 4300 93594 4356 93596
rect 4380 93594 4436 93596
rect 4460 93594 4516 93596
rect 4220 93542 4246 93594
rect 4246 93542 4276 93594
rect 4300 93542 4310 93594
rect 4310 93542 4356 93594
rect 4380 93542 4426 93594
rect 4426 93542 4436 93594
rect 4460 93542 4490 93594
rect 4490 93542 4516 93594
rect 4220 93540 4276 93542
rect 4300 93540 4356 93542
rect 4380 93540 4436 93542
rect 4460 93540 4516 93542
rect 4220 92506 4276 92508
rect 4300 92506 4356 92508
rect 4380 92506 4436 92508
rect 4460 92506 4516 92508
rect 4220 92454 4246 92506
rect 4246 92454 4276 92506
rect 4300 92454 4310 92506
rect 4310 92454 4356 92506
rect 4380 92454 4426 92506
rect 4426 92454 4436 92506
rect 4460 92454 4490 92506
rect 4490 92454 4516 92506
rect 4220 92452 4276 92454
rect 4300 92452 4356 92454
rect 4380 92452 4436 92454
rect 4460 92452 4516 92454
rect 4220 91418 4276 91420
rect 4300 91418 4356 91420
rect 4380 91418 4436 91420
rect 4460 91418 4516 91420
rect 4220 91366 4246 91418
rect 4246 91366 4276 91418
rect 4300 91366 4310 91418
rect 4310 91366 4356 91418
rect 4380 91366 4426 91418
rect 4426 91366 4436 91418
rect 4460 91366 4490 91418
rect 4490 91366 4516 91418
rect 4220 91364 4276 91366
rect 4300 91364 4356 91366
rect 4380 91364 4436 91366
rect 4460 91364 4516 91366
rect 4220 90330 4276 90332
rect 4300 90330 4356 90332
rect 4380 90330 4436 90332
rect 4460 90330 4516 90332
rect 4220 90278 4246 90330
rect 4246 90278 4276 90330
rect 4300 90278 4310 90330
rect 4310 90278 4356 90330
rect 4380 90278 4426 90330
rect 4426 90278 4436 90330
rect 4460 90278 4490 90330
rect 4490 90278 4516 90330
rect 4220 90276 4276 90278
rect 4300 90276 4356 90278
rect 4380 90276 4436 90278
rect 4460 90276 4516 90278
rect 4220 89242 4276 89244
rect 4300 89242 4356 89244
rect 4380 89242 4436 89244
rect 4460 89242 4516 89244
rect 4220 89190 4246 89242
rect 4246 89190 4276 89242
rect 4300 89190 4310 89242
rect 4310 89190 4356 89242
rect 4380 89190 4426 89242
rect 4426 89190 4436 89242
rect 4460 89190 4490 89242
rect 4490 89190 4516 89242
rect 4220 89188 4276 89190
rect 4300 89188 4356 89190
rect 4380 89188 4436 89190
rect 4460 89188 4516 89190
rect 4220 88154 4276 88156
rect 4300 88154 4356 88156
rect 4380 88154 4436 88156
rect 4460 88154 4516 88156
rect 4220 88102 4246 88154
rect 4246 88102 4276 88154
rect 4300 88102 4310 88154
rect 4310 88102 4356 88154
rect 4380 88102 4426 88154
rect 4426 88102 4436 88154
rect 4460 88102 4490 88154
rect 4490 88102 4516 88154
rect 4220 88100 4276 88102
rect 4300 88100 4356 88102
rect 4380 88100 4436 88102
rect 4460 88100 4516 88102
rect 4220 87066 4276 87068
rect 4300 87066 4356 87068
rect 4380 87066 4436 87068
rect 4460 87066 4516 87068
rect 4220 87014 4246 87066
rect 4246 87014 4276 87066
rect 4300 87014 4310 87066
rect 4310 87014 4356 87066
rect 4380 87014 4426 87066
rect 4426 87014 4436 87066
rect 4460 87014 4490 87066
rect 4490 87014 4516 87066
rect 4220 87012 4276 87014
rect 4300 87012 4356 87014
rect 4380 87012 4436 87014
rect 4460 87012 4516 87014
rect 4220 85978 4276 85980
rect 4300 85978 4356 85980
rect 4380 85978 4436 85980
rect 4460 85978 4516 85980
rect 4220 85926 4246 85978
rect 4246 85926 4276 85978
rect 4300 85926 4310 85978
rect 4310 85926 4356 85978
rect 4380 85926 4426 85978
rect 4426 85926 4436 85978
rect 4460 85926 4490 85978
rect 4490 85926 4516 85978
rect 4220 85924 4276 85926
rect 4300 85924 4356 85926
rect 4380 85924 4436 85926
rect 4460 85924 4516 85926
rect 4220 84890 4276 84892
rect 4300 84890 4356 84892
rect 4380 84890 4436 84892
rect 4460 84890 4516 84892
rect 4220 84838 4246 84890
rect 4246 84838 4276 84890
rect 4300 84838 4310 84890
rect 4310 84838 4356 84890
rect 4380 84838 4426 84890
rect 4426 84838 4436 84890
rect 4460 84838 4490 84890
rect 4490 84838 4516 84890
rect 4220 84836 4276 84838
rect 4300 84836 4356 84838
rect 4380 84836 4436 84838
rect 4460 84836 4516 84838
rect 4220 83802 4276 83804
rect 4300 83802 4356 83804
rect 4380 83802 4436 83804
rect 4460 83802 4516 83804
rect 4220 83750 4246 83802
rect 4246 83750 4276 83802
rect 4300 83750 4310 83802
rect 4310 83750 4356 83802
rect 4380 83750 4426 83802
rect 4426 83750 4436 83802
rect 4460 83750 4490 83802
rect 4490 83750 4516 83802
rect 4220 83748 4276 83750
rect 4300 83748 4356 83750
rect 4380 83748 4436 83750
rect 4460 83748 4516 83750
rect 4220 82714 4276 82716
rect 4300 82714 4356 82716
rect 4380 82714 4436 82716
rect 4460 82714 4516 82716
rect 4220 82662 4246 82714
rect 4246 82662 4276 82714
rect 4300 82662 4310 82714
rect 4310 82662 4356 82714
rect 4380 82662 4426 82714
rect 4426 82662 4436 82714
rect 4460 82662 4490 82714
rect 4490 82662 4516 82714
rect 4220 82660 4276 82662
rect 4300 82660 4356 82662
rect 4380 82660 4436 82662
rect 4460 82660 4516 82662
rect 4220 81626 4276 81628
rect 4300 81626 4356 81628
rect 4380 81626 4436 81628
rect 4460 81626 4516 81628
rect 4220 81574 4246 81626
rect 4246 81574 4276 81626
rect 4300 81574 4310 81626
rect 4310 81574 4356 81626
rect 4380 81574 4426 81626
rect 4426 81574 4436 81626
rect 4460 81574 4490 81626
rect 4490 81574 4516 81626
rect 4220 81572 4276 81574
rect 4300 81572 4356 81574
rect 4380 81572 4436 81574
rect 4460 81572 4516 81574
rect 4220 80538 4276 80540
rect 4300 80538 4356 80540
rect 4380 80538 4436 80540
rect 4460 80538 4516 80540
rect 4220 80486 4246 80538
rect 4246 80486 4276 80538
rect 4300 80486 4310 80538
rect 4310 80486 4356 80538
rect 4380 80486 4426 80538
rect 4426 80486 4436 80538
rect 4460 80486 4490 80538
rect 4490 80486 4516 80538
rect 4220 80484 4276 80486
rect 4300 80484 4356 80486
rect 4380 80484 4436 80486
rect 4460 80484 4516 80486
rect 4220 79450 4276 79452
rect 4300 79450 4356 79452
rect 4380 79450 4436 79452
rect 4460 79450 4516 79452
rect 4220 79398 4246 79450
rect 4246 79398 4276 79450
rect 4300 79398 4310 79450
rect 4310 79398 4356 79450
rect 4380 79398 4426 79450
rect 4426 79398 4436 79450
rect 4460 79398 4490 79450
rect 4490 79398 4516 79450
rect 4220 79396 4276 79398
rect 4300 79396 4356 79398
rect 4380 79396 4436 79398
rect 4460 79396 4516 79398
rect 4220 78362 4276 78364
rect 4300 78362 4356 78364
rect 4380 78362 4436 78364
rect 4460 78362 4516 78364
rect 4220 78310 4246 78362
rect 4246 78310 4276 78362
rect 4300 78310 4310 78362
rect 4310 78310 4356 78362
rect 4380 78310 4426 78362
rect 4426 78310 4436 78362
rect 4460 78310 4490 78362
rect 4490 78310 4516 78362
rect 4220 78308 4276 78310
rect 4300 78308 4356 78310
rect 4380 78308 4436 78310
rect 4460 78308 4516 78310
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4246 77274
rect 4246 77222 4276 77274
rect 4300 77222 4310 77274
rect 4310 77222 4356 77274
rect 4380 77222 4426 77274
rect 4426 77222 4436 77274
rect 4460 77222 4490 77274
rect 4490 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4246 76186
rect 4246 76134 4276 76186
rect 4300 76134 4310 76186
rect 4310 76134 4356 76186
rect 4380 76134 4426 76186
rect 4426 76134 4436 76186
rect 4460 76134 4490 76186
rect 4490 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4246 75098
rect 4246 75046 4276 75098
rect 4300 75046 4310 75098
rect 4310 75046 4356 75098
rect 4380 75046 4426 75098
rect 4426 75046 4436 75098
rect 4460 75046 4490 75098
rect 4490 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4246 74010
rect 4246 73958 4276 74010
rect 4300 73958 4310 74010
rect 4310 73958 4356 74010
rect 4380 73958 4426 74010
rect 4426 73958 4436 74010
rect 4460 73958 4490 74010
rect 4490 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4246 72922
rect 4246 72870 4276 72922
rect 4300 72870 4310 72922
rect 4310 72870 4356 72922
rect 4380 72870 4426 72922
rect 4426 72870 4436 72922
rect 4460 72870 4490 72922
rect 4490 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4246 71834
rect 4246 71782 4276 71834
rect 4300 71782 4310 71834
rect 4310 71782 4356 71834
rect 4380 71782 4426 71834
rect 4426 71782 4436 71834
rect 4460 71782 4490 71834
rect 4490 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4246 70746
rect 4246 70694 4276 70746
rect 4300 70694 4310 70746
rect 4310 70694 4356 70746
rect 4380 70694 4426 70746
rect 4426 70694 4436 70746
rect 4460 70694 4490 70746
rect 4490 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4246 69658
rect 4246 69606 4276 69658
rect 4300 69606 4310 69658
rect 4310 69606 4356 69658
rect 4380 69606 4426 69658
rect 4426 69606 4436 69658
rect 4460 69606 4490 69658
rect 4490 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4246 68570
rect 4246 68518 4276 68570
rect 4300 68518 4310 68570
rect 4310 68518 4356 68570
rect 4380 68518 4426 68570
rect 4426 68518 4436 68570
rect 4460 68518 4490 68570
rect 4490 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3054 1264 3110 1320
rect 3330 2080 3386 2136
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19890 117308 19892 117328
rect 19892 117308 19944 117328
rect 19944 117308 19946 117328
rect 19890 117272 19946 117308
rect 19580 116986 19636 116988
rect 19660 116986 19716 116988
rect 19740 116986 19796 116988
rect 19820 116986 19876 116988
rect 19580 116934 19606 116986
rect 19606 116934 19636 116986
rect 19660 116934 19670 116986
rect 19670 116934 19716 116986
rect 19740 116934 19786 116986
rect 19786 116934 19796 116986
rect 19820 116934 19850 116986
rect 19850 116934 19876 116986
rect 19580 116932 19636 116934
rect 19660 116932 19716 116934
rect 19740 116932 19796 116934
rect 19820 116932 19876 116934
rect 19580 115898 19636 115900
rect 19660 115898 19716 115900
rect 19740 115898 19796 115900
rect 19820 115898 19876 115900
rect 19580 115846 19606 115898
rect 19606 115846 19636 115898
rect 19660 115846 19670 115898
rect 19670 115846 19716 115898
rect 19740 115846 19786 115898
rect 19786 115846 19796 115898
rect 19820 115846 19850 115898
rect 19850 115846 19876 115898
rect 19580 115844 19636 115846
rect 19660 115844 19716 115846
rect 19740 115844 19796 115846
rect 19820 115844 19876 115846
rect 19580 114810 19636 114812
rect 19660 114810 19716 114812
rect 19740 114810 19796 114812
rect 19820 114810 19876 114812
rect 19580 114758 19606 114810
rect 19606 114758 19636 114810
rect 19660 114758 19670 114810
rect 19670 114758 19716 114810
rect 19740 114758 19786 114810
rect 19786 114758 19796 114810
rect 19820 114758 19850 114810
rect 19850 114758 19876 114810
rect 19580 114756 19636 114758
rect 19660 114756 19716 114758
rect 19740 114756 19796 114758
rect 19820 114756 19876 114758
rect 20258 115776 20314 115832
rect 20718 114552 20774 114608
rect 21454 116592 21510 116648
rect 20902 115232 20958 115288
rect 22098 116628 22100 116648
rect 22100 116628 22152 116648
rect 22152 116628 22154 116648
rect 22098 116592 22154 116628
rect 21914 116184 21970 116240
rect 19580 113722 19636 113724
rect 19660 113722 19716 113724
rect 19740 113722 19796 113724
rect 19820 113722 19876 113724
rect 19580 113670 19606 113722
rect 19606 113670 19636 113722
rect 19660 113670 19670 113722
rect 19670 113670 19716 113722
rect 19740 113670 19786 113722
rect 19786 113670 19796 113722
rect 19820 113670 19850 113722
rect 19850 113670 19876 113722
rect 19580 113668 19636 113670
rect 19660 113668 19716 113670
rect 19740 113668 19796 113670
rect 19820 113668 19876 113670
rect 10322 18808 10378 18864
rect 13450 19116 13452 19136
rect 13452 19116 13504 19136
rect 13504 19116 13506 19136
rect 13450 19080 13506 19116
rect 14462 28736 14518 28792
rect 19580 112634 19636 112636
rect 19660 112634 19716 112636
rect 19740 112634 19796 112636
rect 19820 112634 19876 112636
rect 19580 112582 19606 112634
rect 19606 112582 19636 112634
rect 19660 112582 19670 112634
rect 19670 112582 19716 112634
rect 19740 112582 19786 112634
rect 19786 112582 19796 112634
rect 19820 112582 19850 112634
rect 19850 112582 19876 112634
rect 19580 112580 19636 112582
rect 19660 112580 19716 112582
rect 19740 112580 19796 112582
rect 19820 112580 19876 112582
rect 19580 111546 19636 111548
rect 19660 111546 19716 111548
rect 19740 111546 19796 111548
rect 19820 111546 19876 111548
rect 19580 111494 19606 111546
rect 19606 111494 19636 111546
rect 19660 111494 19670 111546
rect 19670 111494 19716 111546
rect 19740 111494 19786 111546
rect 19786 111494 19796 111546
rect 19820 111494 19850 111546
rect 19850 111494 19876 111546
rect 19580 111492 19636 111494
rect 19660 111492 19716 111494
rect 19740 111492 19796 111494
rect 19820 111492 19876 111494
rect 19580 110458 19636 110460
rect 19660 110458 19716 110460
rect 19740 110458 19796 110460
rect 19820 110458 19876 110460
rect 19580 110406 19606 110458
rect 19606 110406 19636 110458
rect 19660 110406 19670 110458
rect 19670 110406 19716 110458
rect 19740 110406 19786 110458
rect 19786 110406 19796 110458
rect 19820 110406 19850 110458
rect 19850 110406 19876 110458
rect 19580 110404 19636 110406
rect 19660 110404 19716 110406
rect 19740 110404 19796 110406
rect 19820 110404 19876 110406
rect 19580 109370 19636 109372
rect 19660 109370 19716 109372
rect 19740 109370 19796 109372
rect 19820 109370 19876 109372
rect 19580 109318 19606 109370
rect 19606 109318 19636 109370
rect 19660 109318 19670 109370
rect 19670 109318 19716 109370
rect 19740 109318 19786 109370
rect 19786 109318 19796 109370
rect 19820 109318 19850 109370
rect 19850 109318 19876 109370
rect 19580 109316 19636 109318
rect 19660 109316 19716 109318
rect 19740 109316 19796 109318
rect 19820 109316 19876 109318
rect 19580 108282 19636 108284
rect 19660 108282 19716 108284
rect 19740 108282 19796 108284
rect 19820 108282 19876 108284
rect 19580 108230 19606 108282
rect 19606 108230 19636 108282
rect 19660 108230 19670 108282
rect 19670 108230 19716 108282
rect 19740 108230 19786 108282
rect 19786 108230 19796 108282
rect 19820 108230 19850 108282
rect 19850 108230 19876 108282
rect 19580 108228 19636 108230
rect 19660 108228 19716 108230
rect 19740 108228 19796 108230
rect 19820 108228 19876 108230
rect 19580 107194 19636 107196
rect 19660 107194 19716 107196
rect 19740 107194 19796 107196
rect 19820 107194 19876 107196
rect 19580 107142 19606 107194
rect 19606 107142 19636 107194
rect 19660 107142 19670 107194
rect 19670 107142 19716 107194
rect 19740 107142 19786 107194
rect 19786 107142 19796 107194
rect 19820 107142 19850 107194
rect 19850 107142 19876 107194
rect 19580 107140 19636 107142
rect 19660 107140 19716 107142
rect 19740 107140 19796 107142
rect 19820 107140 19876 107142
rect 19580 106106 19636 106108
rect 19660 106106 19716 106108
rect 19740 106106 19796 106108
rect 19820 106106 19876 106108
rect 19580 106054 19606 106106
rect 19606 106054 19636 106106
rect 19660 106054 19670 106106
rect 19670 106054 19716 106106
rect 19740 106054 19786 106106
rect 19786 106054 19796 106106
rect 19820 106054 19850 106106
rect 19850 106054 19876 106106
rect 19580 106052 19636 106054
rect 19660 106052 19716 106054
rect 19740 106052 19796 106054
rect 19820 106052 19876 106054
rect 19580 105018 19636 105020
rect 19660 105018 19716 105020
rect 19740 105018 19796 105020
rect 19820 105018 19876 105020
rect 19580 104966 19606 105018
rect 19606 104966 19636 105018
rect 19660 104966 19670 105018
rect 19670 104966 19716 105018
rect 19740 104966 19786 105018
rect 19786 104966 19796 105018
rect 19820 104966 19850 105018
rect 19850 104966 19876 105018
rect 19580 104964 19636 104966
rect 19660 104964 19716 104966
rect 19740 104964 19796 104966
rect 19820 104964 19876 104966
rect 19580 103930 19636 103932
rect 19660 103930 19716 103932
rect 19740 103930 19796 103932
rect 19820 103930 19876 103932
rect 19580 103878 19606 103930
rect 19606 103878 19636 103930
rect 19660 103878 19670 103930
rect 19670 103878 19716 103930
rect 19740 103878 19786 103930
rect 19786 103878 19796 103930
rect 19820 103878 19850 103930
rect 19850 103878 19876 103930
rect 19580 103876 19636 103878
rect 19660 103876 19716 103878
rect 19740 103876 19796 103878
rect 19820 103876 19876 103878
rect 17130 21972 17132 21992
rect 17132 21972 17184 21992
rect 17184 21972 17186 21992
rect 17130 21936 17186 21972
rect 17130 21428 17132 21448
rect 17132 21428 17184 21448
rect 17184 21428 17186 21448
rect 17130 21392 17186 21428
rect 17314 23704 17370 23760
rect 17682 21528 17738 21584
rect 17222 19250 17278 19306
rect 17222 19116 17224 19136
rect 17224 19116 17276 19136
rect 17276 19116 17278 19136
rect 17222 19080 17278 19116
rect 17314 18944 17370 19000
rect 19580 102842 19636 102844
rect 19660 102842 19716 102844
rect 19740 102842 19796 102844
rect 19820 102842 19876 102844
rect 19580 102790 19606 102842
rect 19606 102790 19636 102842
rect 19660 102790 19670 102842
rect 19670 102790 19716 102842
rect 19740 102790 19786 102842
rect 19786 102790 19796 102842
rect 19820 102790 19850 102842
rect 19850 102790 19876 102842
rect 19580 102788 19636 102790
rect 19660 102788 19716 102790
rect 19740 102788 19796 102790
rect 19820 102788 19876 102790
rect 19580 101754 19636 101756
rect 19660 101754 19716 101756
rect 19740 101754 19796 101756
rect 19820 101754 19876 101756
rect 19580 101702 19606 101754
rect 19606 101702 19636 101754
rect 19660 101702 19670 101754
rect 19670 101702 19716 101754
rect 19740 101702 19786 101754
rect 19786 101702 19796 101754
rect 19820 101702 19850 101754
rect 19850 101702 19876 101754
rect 19580 101700 19636 101702
rect 19660 101700 19716 101702
rect 19740 101700 19796 101702
rect 19820 101700 19876 101702
rect 19580 100666 19636 100668
rect 19660 100666 19716 100668
rect 19740 100666 19796 100668
rect 19820 100666 19876 100668
rect 19580 100614 19606 100666
rect 19606 100614 19636 100666
rect 19660 100614 19670 100666
rect 19670 100614 19716 100666
rect 19740 100614 19786 100666
rect 19786 100614 19796 100666
rect 19820 100614 19850 100666
rect 19850 100614 19876 100666
rect 19580 100612 19636 100614
rect 19660 100612 19716 100614
rect 19740 100612 19796 100614
rect 19820 100612 19876 100614
rect 19580 99578 19636 99580
rect 19660 99578 19716 99580
rect 19740 99578 19796 99580
rect 19820 99578 19876 99580
rect 19580 99526 19606 99578
rect 19606 99526 19636 99578
rect 19660 99526 19670 99578
rect 19670 99526 19716 99578
rect 19740 99526 19786 99578
rect 19786 99526 19796 99578
rect 19820 99526 19850 99578
rect 19850 99526 19876 99578
rect 19580 99524 19636 99526
rect 19660 99524 19716 99526
rect 19740 99524 19796 99526
rect 19820 99524 19876 99526
rect 19580 98490 19636 98492
rect 19660 98490 19716 98492
rect 19740 98490 19796 98492
rect 19820 98490 19876 98492
rect 19580 98438 19606 98490
rect 19606 98438 19636 98490
rect 19660 98438 19670 98490
rect 19670 98438 19716 98490
rect 19740 98438 19786 98490
rect 19786 98438 19796 98490
rect 19820 98438 19850 98490
rect 19850 98438 19876 98490
rect 19580 98436 19636 98438
rect 19660 98436 19716 98438
rect 19740 98436 19796 98438
rect 19820 98436 19876 98438
rect 19580 97402 19636 97404
rect 19660 97402 19716 97404
rect 19740 97402 19796 97404
rect 19820 97402 19876 97404
rect 19580 97350 19606 97402
rect 19606 97350 19636 97402
rect 19660 97350 19670 97402
rect 19670 97350 19716 97402
rect 19740 97350 19786 97402
rect 19786 97350 19796 97402
rect 19820 97350 19850 97402
rect 19850 97350 19876 97402
rect 19580 97348 19636 97350
rect 19660 97348 19716 97350
rect 19740 97348 19796 97350
rect 19820 97348 19876 97350
rect 19580 96314 19636 96316
rect 19660 96314 19716 96316
rect 19740 96314 19796 96316
rect 19820 96314 19876 96316
rect 19580 96262 19606 96314
rect 19606 96262 19636 96314
rect 19660 96262 19670 96314
rect 19670 96262 19716 96314
rect 19740 96262 19786 96314
rect 19786 96262 19796 96314
rect 19820 96262 19850 96314
rect 19850 96262 19876 96314
rect 19580 96260 19636 96262
rect 19660 96260 19716 96262
rect 19740 96260 19796 96262
rect 19820 96260 19876 96262
rect 19580 95226 19636 95228
rect 19660 95226 19716 95228
rect 19740 95226 19796 95228
rect 19820 95226 19876 95228
rect 19580 95174 19606 95226
rect 19606 95174 19636 95226
rect 19660 95174 19670 95226
rect 19670 95174 19716 95226
rect 19740 95174 19786 95226
rect 19786 95174 19796 95226
rect 19820 95174 19850 95226
rect 19850 95174 19876 95226
rect 19580 95172 19636 95174
rect 19660 95172 19716 95174
rect 19740 95172 19796 95174
rect 19820 95172 19876 95174
rect 19580 94138 19636 94140
rect 19660 94138 19716 94140
rect 19740 94138 19796 94140
rect 19820 94138 19876 94140
rect 19580 94086 19606 94138
rect 19606 94086 19636 94138
rect 19660 94086 19670 94138
rect 19670 94086 19716 94138
rect 19740 94086 19786 94138
rect 19786 94086 19796 94138
rect 19820 94086 19850 94138
rect 19850 94086 19876 94138
rect 19580 94084 19636 94086
rect 19660 94084 19716 94086
rect 19740 94084 19796 94086
rect 19820 94084 19876 94086
rect 18234 28192 18290 28248
rect 18050 23976 18106 24032
rect 18602 21528 18658 21584
rect 18510 21412 18566 21448
rect 18510 21392 18512 21412
rect 18512 21392 18564 21412
rect 18564 21392 18566 21412
rect 18418 18828 18474 18864
rect 18418 18808 18420 18828
rect 18420 18808 18472 18828
rect 18472 18808 18474 18828
rect 18878 23840 18934 23896
rect 18878 21972 18880 21992
rect 18880 21972 18932 21992
rect 18932 21972 18934 21992
rect 18878 21936 18934 21972
rect 18786 21528 18842 21584
rect 19580 93050 19636 93052
rect 19660 93050 19716 93052
rect 19740 93050 19796 93052
rect 19820 93050 19876 93052
rect 19580 92998 19606 93050
rect 19606 92998 19636 93050
rect 19660 92998 19670 93050
rect 19670 92998 19716 93050
rect 19740 92998 19786 93050
rect 19786 92998 19796 93050
rect 19820 92998 19850 93050
rect 19850 92998 19876 93050
rect 19580 92996 19636 92998
rect 19660 92996 19716 92998
rect 19740 92996 19796 92998
rect 19820 92996 19876 92998
rect 19580 91962 19636 91964
rect 19660 91962 19716 91964
rect 19740 91962 19796 91964
rect 19820 91962 19876 91964
rect 19580 91910 19606 91962
rect 19606 91910 19636 91962
rect 19660 91910 19670 91962
rect 19670 91910 19716 91962
rect 19740 91910 19786 91962
rect 19786 91910 19796 91962
rect 19820 91910 19850 91962
rect 19850 91910 19876 91962
rect 19580 91908 19636 91910
rect 19660 91908 19716 91910
rect 19740 91908 19796 91910
rect 19820 91908 19876 91910
rect 19580 90874 19636 90876
rect 19660 90874 19716 90876
rect 19740 90874 19796 90876
rect 19820 90874 19876 90876
rect 19580 90822 19606 90874
rect 19606 90822 19636 90874
rect 19660 90822 19670 90874
rect 19670 90822 19716 90874
rect 19740 90822 19786 90874
rect 19786 90822 19796 90874
rect 19820 90822 19850 90874
rect 19850 90822 19876 90874
rect 19580 90820 19636 90822
rect 19660 90820 19716 90822
rect 19740 90820 19796 90822
rect 19820 90820 19876 90822
rect 19580 89786 19636 89788
rect 19660 89786 19716 89788
rect 19740 89786 19796 89788
rect 19820 89786 19876 89788
rect 19580 89734 19606 89786
rect 19606 89734 19636 89786
rect 19660 89734 19670 89786
rect 19670 89734 19716 89786
rect 19740 89734 19786 89786
rect 19786 89734 19796 89786
rect 19820 89734 19850 89786
rect 19850 89734 19876 89786
rect 19580 89732 19636 89734
rect 19660 89732 19716 89734
rect 19740 89732 19796 89734
rect 19820 89732 19876 89734
rect 19580 88698 19636 88700
rect 19660 88698 19716 88700
rect 19740 88698 19796 88700
rect 19820 88698 19876 88700
rect 19580 88646 19606 88698
rect 19606 88646 19636 88698
rect 19660 88646 19670 88698
rect 19670 88646 19716 88698
rect 19740 88646 19786 88698
rect 19786 88646 19796 88698
rect 19820 88646 19850 88698
rect 19850 88646 19876 88698
rect 19580 88644 19636 88646
rect 19660 88644 19716 88646
rect 19740 88644 19796 88646
rect 19820 88644 19876 88646
rect 19580 87610 19636 87612
rect 19660 87610 19716 87612
rect 19740 87610 19796 87612
rect 19820 87610 19876 87612
rect 19580 87558 19606 87610
rect 19606 87558 19636 87610
rect 19660 87558 19670 87610
rect 19670 87558 19716 87610
rect 19740 87558 19786 87610
rect 19786 87558 19796 87610
rect 19820 87558 19850 87610
rect 19850 87558 19876 87610
rect 19580 87556 19636 87558
rect 19660 87556 19716 87558
rect 19740 87556 19796 87558
rect 19820 87556 19876 87558
rect 19246 23840 19302 23896
rect 19246 21528 19302 21584
rect 19580 86522 19636 86524
rect 19660 86522 19716 86524
rect 19740 86522 19796 86524
rect 19820 86522 19876 86524
rect 19580 86470 19606 86522
rect 19606 86470 19636 86522
rect 19660 86470 19670 86522
rect 19670 86470 19716 86522
rect 19740 86470 19786 86522
rect 19786 86470 19796 86522
rect 19820 86470 19850 86522
rect 19850 86470 19876 86522
rect 19580 86468 19636 86470
rect 19660 86468 19716 86470
rect 19740 86468 19796 86470
rect 19820 86468 19876 86470
rect 19580 85434 19636 85436
rect 19660 85434 19716 85436
rect 19740 85434 19796 85436
rect 19820 85434 19876 85436
rect 19580 85382 19606 85434
rect 19606 85382 19636 85434
rect 19660 85382 19670 85434
rect 19670 85382 19716 85434
rect 19740 85382 19786 85434
rect 19786 85382 19796 85434
rect 19820 85382 19850 85434
rect 19850 85382 19876 85434
rect 19580 85380 19636 85382
rect 19660 85380 19716 85382
rect 19740 85380 19796 85382
rect 19820 85380 19876 85382
rect 19580 84346 19636 84348
rect 19660 84346 19716 84348
rect 19740 84346 19796 84348
rect 19820 84346 19876 84348
rect 19580 84294 19606 84346
rect 19606 84294 19636 84346
rect 19660 84294 19670 84346
rect 19670 84294 19716 84346
rect 19740 84294 19786 84346
rect 19786 84294 19796 84346
rect 19820 84294 19850 84346
rect 19850 84294 19876 84346
rect 19580 84292 19636 84294
rect 19660 84292 19716 84294
rect 19740 84292 19796 84294
rect 19820 84292 19876 84294
rect 19580 83258 19636 83260
rect 19660 83258 19716 83260
rect 19740 83258 19796 83260
rect 19820 83258 19876 83260
rect 19580 83206 19606 83258
rect 19606 83206 19636 83258
rect 19660 83206 19670 83258
rect 19670 83206 19716 83258
rect 19740 83206 19786 83258
rect 19786 83206 19796 83258
rect 19820 83206 19850 83258
rect 19850 83206 19876 83258
rect 19580 83204 19636 83206
rect 19660 83204 19716 83206
rect 19740 83204 19796 83206
rect 19820 83204 19876 83206
rect 19580 82170 19636 82172
rect 19660 82170 19716 82172
rect 19740 82170 19796 82172
rect 19820 82170 19876 82172
rect 19580 82118 19606 82170
rect 19606 82118 19636 82170
rect 19660 82118 19670 82170
rect 19670 82118 19716 82170
rect 19740 82118 19786 82170
rect 19786 82118 19796 82170
rect 19820 82118 19850 82170
rect 19850 82118 19876 82170
rect 19580 82116 19636 82118
rect 19660 82116 19716 82118
rect 19740 82116 19796 82118
rect 19820 82116 19876 82118
rect 19580 81082 19636 81084
rect 19660 81082 19716 81084
rect 19740 81082 19796 81084
rect 19820 81082 19876 81084
rect 19580 81030 19606 81082
rect 19606 81030 19636 81082
rect 19660 81030 19670 81082
rect 19670 81030 19716 81082
rect 19740 81030 19786 81082
rect 19786 81030 19796 81082
rect 19820 81030 19850 81082
rect 19850 81030 19876 81082
rect 19580 81028 19636 81030
rect 19660 81028 19716 81030
rect 19740 81028 19796 81030
rect 19820 81028 19876 81030
rect 19580 79994 19636 79996
rect 19660 79994 19716 79996
rect 19740 79994 19796 79996
rect 19820 79994 19876 79996
rect 19580 79942 19606 79994
rect 19606 79942 19636 79994
rect 19660 79942 19670 79994
rect 19670 79942 19716 79994
rect 19740 79942 19786 79994
rect 19786 79942 19796 79994
rect 19820 79942 19850 79994
rect 19850 79942 19876 79994
rect 19580 79940 19636 79942
rect 19660 79940 19716 79942
rect 19740 79940 19796 79942
rect 19820 79940 19876 79942
rect 19580 78906 19636 78908
rect 19660 78906 19716 78908
rect 19740 78906 19796 78908
rect 19820 78906 19876 78908
rect 19580 78854 19606 78906
rect 19606 78854 19636 78906
rect 19660 78854 19670 78906
rect 19670 78854 19716 78906
rect 19740 78854 19786 78906
rect 19786 78854 19796 78906
rect 19820 78854 19850 78906
rect 19850 78854 19876 78906
rect 19580 78852 19636 78854
rect 19660 78852 19716 78854
rect 19740 78852 19796 78854
rect 19820 78852 19876 78854
rect 19580 77818 19636 77820
rect 19660 77818 19716 77820
rect 19740 77818 19796 77820
rect 19820 77818 19876 77820
rect 19580 77766 19606 77818
rect 19606 77766 19636 77818
rect 19660 77766 19670 77818
rect 19670 77766 19716 77818
rect 19740 77766 19786 77818
rect 19786 77766 19796 77818
rect 19820 77766 19850 77818
rect 19850 77766 19876 77818
rect 19580 77764 19636 77766
rect 19660 77764 19716 77766
rect 19740 77764 19796 77766
rect 19820 77764 19876 77766
rect 19580 76730 19636 76732
rect 19660 76730 19716 76732
rect 19740 76730 19796 76732
rect 19820 76730 19876 76732
rect 19580 76678 19606 76730
rect 19606 76678 19636 76730
rect 19660 76678 19670 76730
rect 19670 76678 19716 76730
rect 19740 76678 19786 76730
rect 19786 76678 19796 76730
rect 19820 76678 19850 76730
rect 19850 76678 19876 76730
rect 19580 76676 19636 76678
rect 19660 76676 19716 76678
rect 19740 76676 19796 76678
rect 19820 76676 19876 76678
rect 19580 75642 19636 75644
rect 19660 75642 19716 75644
rect 19740 75642 19796 75644
rect 19820 75642 19876 75644
rect 19580 75590 19606 75642
rect 19606 75590 19636 75642
rect 19660 75590 19670 75642
rect 19670 75590 19716 75642
rect 19740 75590 19786 75642
rect 19786 75590 19796 75642
rect 19820 75590 19850 75642
rect 19850 75590 19876 75642
rect 19580 75588 19636 75590
rect 19660 75588 19716 75590
rect 19740 75588 19796 75590
rect 19820 75588 19876 75590
rect 19580 74554 19636 74556
rect 19660 74554 19716 74556
rect 19740 74554 19796 74556
rect 19820 74554 19876 74556
rect 19580 74502 19606 74554
rect 19606 74502 19636 74554
rect 19660 74502 19670 74554
rect 19670 74502 19716 74554
rect 19740 74502 19786 74554
rect 19786 74502 19796 74554
rect 19820 74502 19850 74554
rect 19850 74502 19876 74554
rect 19580 74500 19636 74502
rect 19660 74500 19716 74502
rect 19740 74500 19796 74502
rect 19820 74500 19876 74502
rect 19580 73466 19636 73468
rect 19660 73466 19716 73468
rect 19740 73466 19796 73468
rect 19820 73466 19876 73468
rect 19580 73414 19606 73466
rect 19606 73414 19636 73466
rect 19660 73414 19670 73466
rect 19670 73414 19716 73466
rect 19740 73414 19786 73466
rect 19786 73414 19796 73466
rect 19820 73414 19850 73466
rect 19850 73414 19876 73466
rect 19580 73412 19636 73414
rect 19660 73412 19716 73414
rect 19740 73412 19796 73414
rect 19820 73412 19876 73414
rect 19580 72378 19636 72380
rect 19660 72378 19716 72380
rect 19740 72378 19796 72380
rect 19820 72378 19876 72380
rect 19580 72326 19606 72378
rect 19606 72326 19636 72378
rect 19660 72326 19670 72378
rect 19670 72326 19716 72378
rect 19740 72326 19786 72378
rect 19786 72326 19796 72378
rect 19820 72326 19850 72378
rect 19850 72326 19876 72378
rect 19580 72324 19636 72326
rect 19660 72324 19716 72326
rect 19740 72324 19796 72326
rect 19820 72324 19876 72326
rect 19580 71290 19636 71292
rect 19660 71290 19716 71292
rect 19740 71290 19796 71292
rect 19820 71290 19876 71292
rect 19580 71238 19606 71290
rect 19606 71238 19636 71290
rect 19660 71238 19670 71290
rect 19670 71238 19716 71290
rect 19740 71238 19786 71290
rect 19786 71238 19796 71290
rect 19820 71238 19850 71290
rect 19850 71238 19876 71290
rect 19580 71236 19636 71238
rect 19660 71236 19716 71238
rect 19740 71236 19796 71238
rect 19820 71236 19876 71238
rect 19580 70202 19636 70204
rect 19660 70202 19716 70204
rect 19740 70202 19796 70204
rect 19820 70202 19876 70204
rect 19580 70150 19606 70202
rect 19606 70150 19636 70202
rect 19660 70150 19670 70202
rect 19670 70150 19716 70202
rect 19740 70150 19786 70202
rect 19786 70150 19796 70202
rect 19820 70150 19850 70202
rect 19850 70150 19876 70202
rect 19580 70148 19636 70150
rect 19660 70148 19716 70150
rect 19740 70148 19796 70150
rect 19820 70148 19876 70150
rect 19580 69114 19636 69116
rect 19660 69114 19716 69116
rect 19740 69114 19796 69116
rect 19820 69114 19876 69116
rect 19580 69062 19606 69114
rect 19606 69062 19636 69114
rect 19660 69062 19670 69114
rect 19670 69062 19716 69114
rect 19740 69062 19786 69114
rect 19786 69062 19796 69114
rect 19820 69062 19850 69114
rect 19850 69062 19876 69114
rect 19580 69060 19636 69062
rect 19660 69060 19716 69062
rect 19740 69060 19796 69062
rect 19820 69060 19876 69062
rect 19580 68026 19636 68028
rect 19660 68026 19716 68028
rect 19740 68026 19796 68028
rect 19820 68026 19876 68028
rect 19580 67974 19606 68026
rect 19606 67974 19636 68026
rect 19660 67974 19670 68026
rect 19670 67974 19716 68026
rect 19740 67974 19786 68026
rect 19786 67974 19796 68026
rect 19820 67974 19850 68026
rect 19850 67974 19876 68026
rect 19580 67972 19636 67974
rect 19660 67972 19716 67974
rect 19740 67972 19796 67974
rect 19820 67972 19876 67974
rect 19580 66938 19636 66940
rect 19660 66938 19716 66940
rect 19740 66938 19796 66940
rect 19820 66938 19876 66940
rect 19580 66886 19606 66938
rect 19606 66886 19636 66938
rect 19660 66886 19670 66938
rect 19670 66886 19716 66938
rect 19740 66886 19786 66938
rect 19786 66886 19796 66938
rect 19820 66886 19850 66938
rect 19850 66886 19876 66938
rect 19580 66884 19636 66886
rect 19660 66884 19716 66886
rect 19740 66884 19796 66886
rect 19820 66884 19876 66886
rect 19580 65850 19636 65852
rect 19660 65850 19716 65852
rect 19740 65850 19796 65852
rect 19820 65850 19876 65852
rect 19580 65798 19606 65850
rect 19606 65798 19636 65850
rect 19660 65798 19670 65850
rect 19670 65798 19716 65850
rect 19740 65798 19786 65850
rect 19786 65798 19796 65850
rect 19820 65798 19850 65850
rect 19850 65798 19876 65850
rect 19580 65796 19636 65798
rect 19660 65796 19716 65798
rect 19740 65796 19796 65798
rect 19820 65796 19876 65798
rect 19580 64762 19636 64764
rect 19660 64762 19716 64764
rect 19740 64762 19796 64764
rect 19820 64762 19876 64764
rect 19580 64710 19606 64762
rect 19606 64710 19636 64762
rect 19660 64710 19670 64762
rect 19670 64710 19716 64762
rect 19740 64710 19786 64762
rect 19786 64710 19796 64762
rect 19820 64710 19850 64762
rect 19850 64710 19876 64762
rect 19580 64708 19636 64710
rect 19660 64708 19716 64710
rect 19740 64708 19796 64710
rect 19820 64708 19876 64710
rect 19580 63674 19636 63676
rect 19660 63674 19716 63676
rect 19740 63674 19796 63676
rect 19820 63674 19876 63676
rect 19580 63622 19606 63674
rect 19606 63622 19636 63674
rect 19660 63622 19670 63674
rect 19670 63622 19716 63674
rect 19740 63622 19786 63674
rect 19786 63622 19796 63674
rect 19820 63622 19850 63674
rect 19850 63622 19876 63674
rect 19580 63620 19636 63622
rect 19660 63620 19716 63622
rect 19740 63620 19796 63622
rect 19820 63620 19876 63622
rect 19580 62586 19636 62588
rect 19660 62586 19716 62588
rect 19740 62586 19796 62588
rect 19820 62586 19876 62588
rect 19580 62534 19606 62586
rect 19606 62534 19636 62586
rect 19660 62534 19670 62586
rect 19670 62534 19716 62586
rect 19740 62534 19786 62586
rect 19786 62534 19796 62586
rect 19820 62534 19850 62586
rect 19850 62534 19876 62586
rect 19580 62532 19636 62534
rect 19660 62532 19716 62534
rect 19740 62532 19796 62534
rect 19820 62532 19876 62534
rect 19580 61498 19636 61500
rect 19660 61498 19716 61500
rect 19740 61498 19796 61500
rect 19820 61498 19876 61500
rect 19580 61446 19606 61498
rect 19606 61446 19636 61498
rect 19660 61446 19670 61498
rect 19670 61446 19716 61498
rect 19740 61446 19786 61498
rect 19786 61446 19796 61498
rect 19820 61446 19850 61498
rect 19850 61446 19876 61498
rect 19580 61444 19636 61446
rect 19660 61444 19716 61446
rect 19740 61444 19796 61446
rect 19820 61444 19876 61446
rect 19580 60410 19636 60412
rect 19660 60410 19716 60412
rect 19740 60410 19796 60412
rect 19820 60410 19876 60412
rect 19580 60358 19606 60410
rect 19606 60358 19636 60410
rect 19660 60358 19670 60410
rect 19670 60358 19716 60410
rect 19740 60358 19786 60410
rect 19786 60358 19796 60410
rect 19820 60358 19850 60410
rect 19850 60358 19876 60410
rect 19580 60356 19636 60358
rect 19660 60356 19716 60358
rect 19740 60356 19796 60358
rect 19820 60356 19876 60358
rect 19580 59322 19636 59324
rect 19660 59322 19716 59324
rect 19740 59322 19796 59324
rect 19820 59322 19876 59324
rect 19580 59270 19606 59322
rect 19606 59270 19636 59322
rect 19660 59270 19670 59322
rect 19670 59270 19716 59322
rect 19740 59270 19786 59322
rect 19786 59270 19796 59322
rect 19820 59270 19850 59322
rect 19850 59270 19876 59322
rect 19580 59268 19636 59270
rect 19660 59268 19716 59270
rect 19740 59268 19796 59270
rect 19820 59268 19876 59270
rect 19580 58234 19636 58236
rect 19660 58234 19716 58236
rect 19740 58234 19796 58236
rect 19820 58234 19876 58236
rect 19580 58182 19606 58234
rect 19606 58182 19636 58234
rect 19660 58182 19670 58234
rect 19670 58182 19716 58234
rect 19740 58182 19786 58234
rect 19786 58182 19796 58234
rect 19820 58182 19850 58234
rect 19850 58182 19876 58234
rect 19580 58180 19636 58182
rect 19660 58180 19716 58182
rect 19740 58180 19796 58182
rect 19820 58180 19876 58182
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 19982 48456 20038 48512
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 19890 48184 19946 48240
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19614 28600 19670 28656
rect 19798 28620 19854 28656
rect 19798 28600 19800 28620
rect 19800 28600 19852 28620
rect 19852 28600 19854 28620
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19614 27512 19670 27568
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19798 24112 19854 24168
rect 19614 24012 19616 24032
rect 19616 24012 19668 24032
rect 19668 24012 19670 24032
rect 19614 23976 19670 24012
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19522 19216 19578 19272
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19522 18808 19578 18864
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19982 28756 20038 28792
rect 19982 28736 19984 28756
rect 19984 28736 20036 28756
rect 20036 28736 20038 28756
rect 20074 28600 20130 28656
rect 20074 27668 20130 27704
rect 20074 27648 20076 27668
rect 20076 27648 20128 27668
rect 20128 27648 20130 27668
rect 19982 23840 20038 23896
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 20810 33088 20866 33144
rect 20718 23704 20774 23760
rect 20902 24792 20958 24848
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 21270 25880 21326 25936
rect 22098 115504 22154 115560
rect 22006 115368 22062 115424
rect 22558 117136 22614 117192
rect 23202 117272 23258 117328
rect 23202 117000 23258 117056
rect 23294 115096 23350 115152
rect 23938 115776 23994 115832
rect 24490 115912 24546 115968
rect 25134 116864 25190 116920
rect 25502 116184 25558 116240
rect 26146 115368 26202 115424
rect 26422 115504 26478 115560
rect 27158 117000 27214 117056
rect 27710 114552 27766 114608
rect 28354 116864 28410 116920
rect 22098 41692 22100 41712
rect 22100 41692 22152 41712
rect 22152 41692 22154 41712
rect 22098 41656 22154 41692
rect 21638 31864 21694 31920
rect 21454 28056 21510 28112
rect 21454 24792 21510 24848
rect 21914 37884 21916 37904
rect 21916 37884 21968 37904
rect 21968 37884 21970 37904
rect 21914 37848 21970 37884
rect 21822 26968 21878 27024
rect 21730 26424 21786 26480
rect 22282 38528 22338 38584
rect 22282 38292 22284 38312
rect 22284 38292 22336 38312
rect 22336 38292 22338 38312
rect 22282 38256 22338 38292
rect 22282 37732 22338 37768
rect 22282 37712 22284 37732
rect 22284 37712 22336 37732
rect 22336 37712 22338 37732
rect 22282 34312 22338 34368
rect 22374 31048 22430 31104
rect 22282 28736 22338 28792
rect 22558 29008 22614 29064
rect 22466 28908 22468 28928
rect 22468 28908 22520 28928
rect 22520 28908 22522 28928
rect 22466 28872 22522 28908
rect 22834 38936 22890 38992
rect 22558 28620 22614 28656
rect 22558 28600 22560 28620
rect 22560 28600 22612 28620
rect 22612 28600 22614 28620
rect 22098 28212 22154 28248
rect 22098 28192 22100 28212
rect 22100 28192 22152 28212
rect 22152 28192 22154 28212
rect 22006 27784 22062 27840
rect 22006 25064 22062 25120
rect 22374 26424 22430 26480
rect 22006 24148 22008 24168
rect 22008 24148 22060 24168
rect 22060 24148 22062 24168
rect 22006 24112 22062 24148
rect 22834 32988 22836 33008
rect 22836 32988 22888 33008
rect 22888 32988 22890 33008
rect 22834 32952 22890 32988
rect 23018 38936 23074 38992
rect 23294 38936 23350 38992
rect 23110 38392 23166 38448
rect 23386 38548 23442 38584
rect 23386 38528 23388 38548
rect 23388 38528 23440 38548
rect 23440 38528 23442 38548
rect 23202 38256 23258 38312
rect 23386 37732 23442 37768
rect 23386 37712 23388 37732
rect 23388 37712 23440 37732
rect 23440 37712 23442 37732
rect 23386 32000 23442 32056
rect 23110 27512 23166 27568
rect 23570 31592 23626 31648
rect 23570 28600 23626 28656
rect 23294 22208 23350 22264
rect 22190 3476 22192 3496
rect 22192 3476 22244 3496
rect 22244 3476 22246 3496
rect 22190 3440 22246 3476
rect 24214 37884 24216 37904
rect 24216 37884 24268 37904
rect 24268 37884 24270 37904
rect 24214 37848 24270 37884
rect 24490 37712 24546 37768
rect 24398 34448 24454 34504
rect 24306 32292 24362 32328
rect 24306 32272 24308 32292
rect 24308 32272 24360 32292
rect 24360 32272 24362 32292
rect 23938 27512 23994 27568
rect 24214 27648 24270 27704
rect 24490 28872 24546 28928
rect 24214 22208 24270 22264
rect 24858 25880 24914 25936
rect 28262 115912 28318 115968
rect 28814 115232 28870 115288
rect 28998 115096 29054 115152
rect 25502 81640 25558 81696
rect 25502 79464 25558 79520
rect 25594 57024 25650 57080
rect 25226 32444 25228 32464
rect 25228 32444 25280 32464
rect 25280 32444 25282 32464
rect 25226 32408 25282 32444
rect 25410 32272 25466 32328
rect 25226 29008 25282 29064
rect 24950 23840 25006 23896
rect 25962 84224 26018 84280
rect 25870 38256 25926 38312
rect 24398 3440 24454 3496
rect 26054 79872 26110 79928
rect 26054 32408 26110 32464
rect 26514 79600 26570 79656
rect 26422 78512 26478 78568
rect 26238 56888 26294 56944
rect 26514 56908 26570 56944
rect 26514 56888 26516 56908
rect 26516 56888 26568 56908
rect 26568 56888 26570 56908
rect 26514 56752 26570 56808
rect 26238 41248 26294 41304
rect 26514 42644 26516 42664
rect 26516 42644 26568 42664
rect 26568 42644 26570 42664
rect 26514 42608 26570 42644
rect 26606 41676 26662 41712
rect 26606 41656 26608 41676
rect 26608 41656 26660 41676
rect 26660 41656 26662 41676
rect 27158 86128 27214 86184
rect 26882 34312 26938 34368
rect 26882 34176 26938 34232
rect 26698 34040 26754 34096
rect 26882 32952 26938 33008
rect 27158 41384 27214 41440
rect 26974 32564 27030 32600
rect 26974 32544 26976 32564
rect 26976 32544 27028 32564
rect 27028 32544 27030 32564
rect 26974 32428 27030 32464
rect 26974 32408 26976 32428
rect 26976 32408 27028 32428
rect 27028 32408 27030 32428
rect 26974 32272 27030 32328
rect 26974 32000 27030 32056
rect 26790 31456 26846 31512
rect 26882 31356 26884 31376
rect 26884 31356 26936 31376
rect 26936 31356 26938 31376
rect 26882 31320 26938 31356
rect 26606 28464 26662 28520
rect 27066 28192 27122 28248
rect 27526 87796 27528 87816
rect 27528 87796 27580 87816
rect 27580 87796 27582 87816
rect 27526 87760 27582 87796
rect 27618 86672 27674 86728
rect 27618 86264 27674 86320
rect 27526 84668 27528 84688
rect 27528 84668 27580 84688
rect 27580 84668 27582 84688
rect 27526 84632 27582 84668
rect 27434 81368 27490 81424
rect 27342 80824 27398 80880
rect 27434 79736 27490 79792
rect 27434 79600 27490 79656
rect 27434 57976 27490 58032
rect 27434 57160 27490 57216
rect 27526 56752 27582 56808
rect 27342 42644 27344 42664
rect 27344 42644 27396 42664
rect 27396 42644 27398 42664
rect 27342 42608 27398 42644
rect 27342 38428 27344 38448
rect 27344 38428 27396 38448
rect 27396 38428 27398 38448
rect 27342 38392 27398 38428
rect 27434 34040 27490 34096
rect 27342 32544 27398 32600
rect 27710 41520 27766 41576
rect 28170 87932 28172 87952
rect 28172 87932 28224 87952
rect 28224 87932 28226 87952
rect 28170 87896 28226 87932
rect 28170 87760 28226 87816
rect 28262 86264 28318 86320
rect 28262 83952 28318 84008
rect 28262 83408 28318 83464
rect 28170 82184 28226 82240
rect 28170 80044 28172 80064
rect 28172 80044 28224 80064
rect 28224 80044 28226 80064
rect 28170 80008 28226 80044
rect 28170 79600 28226 79656
rect 28170 79192 28226 79248
rect 28170 79056 28226 79112
rect 27894 41248 27950 41304
rect 27618 33360 27674 33416
rect 27434 31456 27490 31512
rect 27066 27784 27122 27840
rect 27710 32836 27766 32872
rect 27710 32816 27712 32836
rect 27712 32816 27764 32836
rect 27764 32816 27766 32836
rect 27986 33224 28042 33280
rect 27986 33088 28042 33144
rect 27986 32716 27988 32736
rect 27988 32716 28040 32736
rect 28040 32716 28042 32736
rect 27986 32680 28042 32716
rect 27986 32308 27988 32328
rect 27988 32308 28040 32328
rect 28040 32308 28042 32328
rect 27986 32272 28042 32308
rect 27618 29280 27674 29336
rect 27894 31592 27950 31648
rect 27894 31356 27896 31376
rect 27896 31356 27948 31376
rect 27948 31356 27950 31376
rect 27894 31320 27950 31356
rect 27802 29144 27858 29200
rect 27802 28872 27858 28928
rect 27618 28600 27674 28656
rect 27434 26968 27490 27024
rect 26146 3032 26202 3088
rect 27710 27784 27766 27840
rect 28446 84224 28502 84280
rect 28446 79872 28502 79928
rect 28354 79192 28410 79248
rect 28262 34176 28318 34232
rect 28814 87932 28816 87952
rect 28816 87932 28868 87952
rect 28868 87932 28870 87952
rect 28814 87896 28870 87932
rect 28906 86692 28962 86728
rect 28906 86672 28908 86692
rect 28908 86672 28960 86692
rect 28960 86672 28962 86692
rect 28906 86128 28962 86184
rect 28814 85448 28870 85504
rect 28630 83408 28686 83464
rect 28630 83136 28686 83192
rect 28722 82220 28724 82240
rect 28724 82220 28776 82240
rect 28776 82220 28778 82240
rect 28722 82184 28778 82220
rect 28630 80008 28686 80064
rect 28630 79464 28686 79520
rect 28630 79192 28686 79248
rect 28630 57024 28686 57080
rect 28630 43288 28686 43344
rect 28446 37712 28502 37768
rect 28630 41792 28686 41848
rect 28630 38528 28686 38584
rect 28998 84496 29054 84552
rect 29274 86284 29330 86320
rect 29274 86264 29277 86284
rect 29277 86264 29329 86284
rect 29329 86264 29330 86284
rect 29274 86148 29330 86184
rect 29274 86128 29276 86148
rect 29276 86128 29328 86148
rect 29328 86128 29330 86148
rect 29090 83988 29092 84008
rect 29092 83988 29144 84008
rect 29144 83988 29146 84008
rect 29090 83952 29146 83988
rect 29274 85448 29330 85504
rect 29366 84632 29422 84688
rect 29366 84224 29422 84280
rect 29182 81504 29238 81560
rect 28998 79636 29000 79656
rect 29000 79636 29052 79656
rect 29052 79636 29054 79656
rect 28998 79600 29054 79636
rect 29274 80280 29330 80336
rect 29090 79056 29146 79112
rect 28998 78920 29054 78976
rect 28998 51312 29054 51368
rect 28906 43288 28962 43344
rect 29642 83680 29698 83736
rect 29642 83544 29698 83600
rect 29642 81368 29698 81424
rect 29366 51584 29422 51640
rect 29182 41520 29238 41576
rect 28906 38800 28962 38856
rect 28814 38528 28870 38584
rect 28630 33632 28686 33688
rect 28262 33088 28318 33144
rect 28354 31864 28410 31920
rect 28630 33360 28686 33416
rect 28538 33224 28594 33280
rect 28538 32816 28594 32872
rect 28630 32172 28632 32192
rect 28632 32172 28684 32192
rect 28684 32172 28686 32192
rect 28630 32136 28686 32172
rect 28906 38256 28962 38312
rect 28814 34448 28870 34504
rect 28446 3032 28502 3088
rect 29458 32544 29514 32600
rect 30654 116184 30710 116240
rect 31206 114008 31262 114064
rect 29734 38120 29790 38176
rect 30102 80416 30158 80472
rect 29918 37984 29974 38040
rect 29826 37168 29882 37224
rect 30010 37440 30066 37496
rect 29734 31048 29790 31104
rect 30378 84496 30434 84552
rect 30378 83680 30434 83736
rect 30286 80012 30342 80068
rect 30378 79600 30434 79656
rect 30378 78920 30434 78976
rect 30378 39344 30434 39400
rect 30194 37032 30250 37088
rect 30654 80416 30710 80472
rect 30746 40840 30802 40896
rect 30562 39344 30618 39400
rect 30654 37848 30710 37904
rect 30930 40840 30986 40896
rect 30930 40704 30986 40760
rect 30838 37848 30894 37904
rect 31206 83816 31262 83872
rect 31114 81504 31170 81560
rect 31206 80980 31262 81016
rect 31206 80960 31208 80980
rect 31208 80960 31260 80980
rect 31260 80960 31262 80980
rect 31482 83952 31538 84008
rect 31390 80416 31446 80472
rect 31390 80316 31392 80336
rect 31392 80316 31444 80336
rect 31444 80316 31446 80336
rect 31390 80280 31446 80316
rect 31114 40704 31170 40760
rect 31114 40024 31170 40080
rect 31758 62464 31814 62520
rect 31758 43152 31814 43208
rect 31942 29144 31998 29200
rect 32494 86964 32550 87000
rect 32494 86944 32496 86964
rect 32496 86944 32548 86964
rect 32548 86944 32550 86964
rect 32770 86708 32772 86728
rect 32772 86708 32824 86728
rect 32824 86708 32826 86728
rect 32770 86672 32826 86708
rect 32402 78784 32458 78840
rect 32310 28636 32312 28656
rect 32312 28636 32364 28656
rect 32364 28636 32366 28656
rect 32310 28600 32366 28636
rect 34518 117952 34574 118008
rect 33322 44396 33378 44432
rect 33322 44376 33324 44396
rect 33324 44376 33376 44396
rect 33376 44376 33378 44396
rect 33322 35400 33378 35456
rect 33690 80960 33746 81016
rect 34702 118768 34758 118824
rect 34940 117530 34996 117532
rect 35020 117530 35076 117532
rect 35100 117530 35156 117532
rect 35180 117530 35236 117532
rect 34940 117478 34966 117530
rect 34966 117478 34996 117530
rect 35020 117478 35030 117530
rect 35030 117478 35076 117530
rect 35100 117478 35146 117530
rect 35146 117478 35156 117530
rect 35180 117478 35210 117530
rect 35210 117478 35236 117530
rect 34940 117476 34996 117478
rect 35020 117476 35076 117478
rect 35100 117476 35156 117478
rect 35180 117476 35236 117478
rect 33966 86964 34022 87000
rect 33966 86944 33968 86964
rect 33968 86944 34020 86964
rect 34020 86944 34022 86964
rect 33966 81640 34022 81696
rect 33690 2760 33746 2816
rect 34150 39480 34206 39536
rect 34334 38936 34390 38992
rect 34334 38664 34390 38720
rect 34334 35400 34390 35456
rect 34940 116442 34996 116444
rect 35020 116442 35076 116444
rect 35100 116442 35156 116444
rect 35180 116442 35236 116444
rect 34940 116390 34966 116442
rect 34966 116390 34996 116442
rect 35020 116390 35030 116442
rect 35030 116390 35076 116442
rect 35100 116390 35146 116442
rect 35146 116390 35156 116442
rect 35180 116390 35210 116442
rect 35210 116390 35236 116442
rect 34940 116388 34996 116390
rect 35020 116388 35076 116390
rect 35100 116388 35156 116390
rect 35180 116388 35236 116390
rect 35346 116184 35402 116240
rect 34940 115354 34996 115356
rect 35020 115354 35076 115356
rect 35100 115354 35156 115356
rect 35180 115354 35236 115356
rect 34940 115302 34966 115354
rect 34966 115302 34996 115354
rect 35020 115302 35030 115354
rect 35030 115302 35076 115354
rect 35100 115302 35146 115354
rect 35146 115302 35156 115354
rect 35180 115302 35210 115354
rect 35210 115302 35236 115354
rect 34940 115300 34996 115302
rect 35020 115300 35076 115302
rect 35100 115300 35156 115302
rect 35180 115300 35236 115302
rect 34702 87216 34758 87272
rect 34702 86944 34758 87000
rect 34940 114266 34996 114268
rect 35020 114266 35076 114268
rect 35100 114266 35156 114268
rect 35180 114266 35236 114268
rect 34940 114214 34966 114266
rect 34966 114214 34996 114266
rect 35020 114214 35030 114266
rect 35030 114214 35076 114266
rect 35100 114214 35146 114266
rect 35146 114214 35156 114266
rect 35180 114214 35210 114266
rect 35210 114214 35236 114266
rect 34940 114212 34996 114214
rect 35020 114212 35076 114214
rect 35100 114212 35156 114214
rect 35180 114212 35236 114214
rect 34940 113178 34996 113180
rect 35020 113178 35076 113180
rect 35100 113178 35156 113180
rect 35180 113178 35236 113180
rect 34940 113126 34966 113178
rect 34966 113126 34996 113178
rect 35020 113126 35030 113178
rect 35030 113126 35076 113178
rect 35100 113126 35146 113178
rect 35146 113126 35156 113178
rect 35180 113126 35210 113178
rect 35210 113126 35236 113178
rect 34940 113124 34996 113126
rect 35020 113124 35076 113126
rect 35100 113124 35156 113126
rect 35180 113124 35236 113126
rect 34940 112090 34996 112092
rect 35020 112090 35076 112092
rect 35100 112090 35156 112092
rect 35180 112090 35236 112092
rect 34940 112038 34966 112090
rect 34966 112038 34996 112090
rect 35020 112038 35030 112090
rect 35030 112038 35076 112090
rect 35100 112038 35146 112090
rect 35146 112038 35156 112090
rect 35180 112038 35210 112090
rect 35210 112038 35236 112090
rect 34940 112036 34996 112038
rect 35020 112036 35076 112038
rect 35100 112036 35156 112038
rect 35180 112036 35236 112038
rect 34940 111002 34996 111004
rect 35020 111002 35076 111004
rect 35100 111002 35156 111004
rect 35180 111002 35236 111004
rect 34940 110950 34966 111002
rect 34966 110950 34996 111002
rect 35020 110950 35030 111002
rect 35030 110950 35076 111002
rect 35100 110950 35146 111002
rect 35146 110950 35156 111002
rect 35180 110950 35210 111002
rect 35210 110950 35236 111002
rect 34940 110948 34996 110950
rect 35020 110948 35076 110950
rect 35100 110948 35156 110950
rect 35180 110948 35236 110950
rect 34940 109914 34996 109916
rect 35020 109914 35076 109916
rect 35100 109914 35156 109916
rect 35180 109914 35236 109916
rect 34940 109862 34966 109914
rect 34966 109862 34996 109914
rect 35020 109862 35030 109914
rect 35030 109862 35076 109914
rect 35100 109862 35146 109914
rect 35146 109862 35156 109914
rect 35180 109862 35210 109914
rect 35210 109862 35236 109914
rect 34940 109860 34996 109862
rect 35020 109860 35076 109862
rect 35100 109860 35156 109862
rect 35180 109860 35236 109862
rect 34940 108826 34996 108828
rect 35020 108826 35076 108828
rect 35100 108826 35156 108828
rect 35180 108826 35236 108828
rect 34940 108774 34966 108826
rect 34966 108774 34996 108826
rect 35020 108774 35030 108826
rect 35030 108774 35076 108826
rect 35100 108774 35146 108826
rect 35146 108774 35156 108826
rect 35180 108774 35210 108826
rect 35210 108774 35236 108826
rect 34940 108772 34996 108774
rect 35020 108772 35076 108774
rect 35100 108772 35156 108774
rect 35180 108772 35236 108774
rect 34940 107738 34996 107740
rect 35020 107738 35076 107740
rect 35100 107738 35156 107740
rect 35180 107738 35236 107740
rect 34940 107686 34966 107738
rect 34966 107686 34996 107738
rect 35020 107686 35030 107738
rect 35030 107686 35076 107738
rect 35100 107686 35146 107738
rect 35146 107686 35156 107738
rect 35180 107686 35210 107738
rect 35210 107686 35236 107738
rect 34940 107684 34996 107686
rect 35020 107684 35076 107686
rect 35100 107684 35156 107686
rect 35180 107684 35236 107686
rect 34940 106650 34996 106652
rect 35020 106650 35076 106652
rect 35100 106650 35156 106652
rect 35180 106650 35236 106652
rect 34940 106598 34966 106650
rect 34966 106598 34996 106650
rect 35020 106598 35030 106650
rect 35030 106598 35076 106650
rect 35100 106598 35146 106650
rect 35146 106598 35156 106650
rect 35180 106598 35210 106650
rect 35210 106598 35236 106650
rect 34940 106596 34996 106598
rect 35020 106596 35076 106598
rect 35100 106596 35156 106598
rect 35180 106596 35236 106598
rect 34940 105562 34996 105564
rect 35020 105562 35076 105564
rect 35100 105562 35156 105564
rect 35180 105562 35236 105564
rect 34940 105510 34966 105562
rect 34966 105510 34996 105562
rect 35020 105510 35030 105562
rect 35030 105510 35076 105562
rect 35100 105510 35146 105562
rect 35146 105510 35156 105562
rect 35180 105510 35210 105562
rect 35210 105510 35236 105562
rect 34940 105508 34996 105510
rect 35020 105508 35076 105510
rect 35100 105508 35156 105510
rect 35180 105508 35236 105510
rect 34940 104474 34996 104476
rect 35020 104474 35076 104476
rect 35100 104474 35156 104476
rect 35180 104474 35236 104476
rect 34940 104422 34966 104474
rect 34966 104422 34996 104474
rect 35020 104422 35030 104474
rect 35030 104422 35076 104474
rect 35100 104422 35146 104474
rect 35146 104422 35156 104474
rect 35180 104422 35210 104474
rect 35210 104422 35236 104474
rect 34940 104420 34996 104422
rect 35020 104420 35076 104422
rect 35100 104420 35156 104422
rect 35180 104420 35236 104422
rect 34940 103386 34996 103388
rect 35020 103386 35076 103388
rect 35100 103386 35156 103388
rect 35180 103386 35236 103388
rect 34940 103334 34966 103386
rect 34966 103334 34996 103386
rect 35020 103334 35030 103386
rect 35030 103334 35076 103386
rect 35100 103334 35146 103386
rect 35146 103334 35156 103386
rect 35180 103334 35210 103386
rect 35210 103334 35236 103386
rect 34940 103332 34996 103334
rect 35020 103332 35076 103334
rect 35100 103332 35156 103334
rect 35180 103332 35236 103334
rect 34940 102298 34996 102300
rect 35020 102298 35076 102300
rect 35100 102298 35156 102300
rect 35180 102298 35236 102300
rect 34940 102246 34966 102298
rect 34966 102246 34996 102298
rect 35020 102246 35030 102298
rect 35030 102246 35076 102298
rect 35100 102246 35146 102298
rect 35146 102246 35156 102298
rect 35180 102246 35210 102298
rect 35210 102246 35236 102298
rect 34940 102244 34996 102246
rect 35020 102244 35076 102246
rect 35100 102244 35156 102246
rect 35180 102244 35236 102246
rect 34940 101210 34996 101212
rect 35020 101210 35076 101212
rect 35100 101210 35156 101212
rect 35180 101210 35236 101212
rect 34940 101158 34966 101210
rect 34966 101158 34996 101210
rect 35020 101158 35030 101210
rect 35030 101158 35076 101210
rect 35100 101158 35146 101210
rect 35146 101158 35156 101210
rect 35180 101158 35210 101210
rect 35210 101158 35236 101210
rect 34940 101156 34996 101158
rect 35020 101156 35076 101158
rect 35100 101156 35156 101158
rect 35180 101156 35236 101158
rect 34940 100122 34996 100124
rect 35020 100122 35076 100124
rect 35100 100122 35156 100124
rect 35180 100122 35236 100124
rect 34940 100070 34966 100122
rect 34966 100070 34996 100122
rect 35020 100070 35030 100122
rect 35030 100070 35076 100122
rect 35100 100070 35146 100122
rect 35146 100070 35156 100122
rect 35180 100070 35210 100122
rect 35210 100070 35236 100122
rect 34940 100068 34996 100070
rect 35020 100068 35076 100070
rect 35100 100068 35156 100070
rect 35180 100068 35236 100070
rect 34940 99034 34996 99036
rect 35020 99034 35076 99036
rect 35100 99034 35156 99036
rect 35180 99034 35236 99036
rect 34940 98982 34966 99034
rect 34966 98982 34996 99034
rect 35020 98982 35030 99034
rect 35030 98982 35076 99034
rect 35100 98982 35146 99034
rect 35146 98982 35156 99034
rect 35180 98982 35210 99034
rect 35210 98982 35236 99034
rect 34940 98980 34996 98982
rect 35020 98980 35076 98982
rect 35100 98980 35156 98982
rect 35180 98980 35236 98982
rect 34940 97946 34996 97948
rect 35020 97946 35076 97948
rect 35100 97946 35156 97948
rect 35180 97946 35236 97948
rect 34940 97894 34966 97946
rect 34966 97894 34996 97946
rect 35020 97894 35030 97946
rect 35030 97894 35076 97946
rect 35100 97894 35146 97946
rect 35146 97894 35156 97946
rect 35180 97894 35210 97946
rect 35210 97894 35236 97946
rect 34940 97892 34996 97894
rect 35020 97892 35076 97894
rect 35100 97892 35156 97894
rect 35180 97892 35236 97894
rect 34940 96858 34996 96860
rect 35020 96858 35076 96860
rect 35100 96858 35156 96860
rect 35180 96858 35236 96860
rect 34940 96806 34966 96858
rect 34966 96806 34996 96858
rect 35020 96806 35030 96858
rect 35030 96806 35076 96858
rect 35100 96806 35146 96858
rect 35146 96806 35156 96858
rect 35180 96806 35210 96858
rect 35210 96806 35236 96858
rect 34940 96804 34996 96806
rect 35020 96804 35076 96806
rect 35100 96804 35156 96806
rect 35180 96804 35236 96806
rect 34940 95770 34996 95772
rect 35020 95770 35076 95772
rect 35100 95770 35156 95772
rect 35180 95770 35236 95772
rect 34940 95718 34966 95770
rect 34966 95718 34996 95770
rect 35020 95718 35030 95770
rect 35030 95718 35076 95770
rect 35100 95718 35146 95770
rect 35146 95718 35156 95770
rect 35180 95718 35210 95770
rect 35210 95718 35236 95770
rect 34940 95716 34996 95718
rect 35020 95716 35076 95718
rect 35100 95716 35156 95718
rect 35180 95716 35236 95718
rect 34940 94682 34996 94684
rect 35020 94682 35076 94684
rect 35100 94682 35156 94684
rect 35180 94682 35236 94684
rect 34940 94630 34966 94682
rect 34966 94630 34996 94682
rect 35020 94630 35030 94682
rect 35030 94630 35076 94682
rect 35100 94630 35146 94682
rect 35146 94630 35156 94682
rect 35180 94630 35210 94682
rect 35210 94630 35236 94682
rect 34940 94628 34996 94630
rect 35020 94628 35076 94630
rect 35100 94628 35156 94630
rect 35180 94628 35236 94630
rect 34940 93594 34996 93596
rect 35020 93594 35076 93596
rect 35100 93594 35156 93596
rect 35180 93594 35236 93596
rect 34940 93542 34966 93594
rect 34966 93542 34996 93594
rect 35020 93542 35030 93594
rect 35030 93542 35076 93594
rect 35100 93542 35146 93594
rect 35146 93542 35156 93594
rect 35180 93542 35210 93594
rect 35210 93542 35236 93594
rect 34940 93540 34996 93542
rect 35020 93540 35076 93542
rect 35100 93540 35156 93542
rect 35180 93540 35236 93542
rect 34940 92506 34996 92508
rect 35020 92506 35076 92508
rect 35100 92506 35156 92508
rect 35180 92506 35236 92508
rect 34940 92454 34966 92506
rect 34966 92454 34996 92506
rect 35020 92454 35030 92506
rect 35030 92454 35076 92506
rect 35100 92454 35146 92506
rect 35146 92454 35156 92506
rect 35180 92454 35210 92506
rect 35210 92454 35236 92506
rect 34940 92452 34996 92454
rect 35020 92452 35076 92454
rect 35100 92452 35156 92454
rect 35180 92452 35236 92454
rect 34940 91418 34996 91420
rect 35020 91418 35076 91420
rect 35100 91418 35156 91420
rect 35180 91418 35236 91420
rect 34940 91366 34966 91418
rect 34966 91366 34996 91418
rect 35020 91366 35030 91418
rect 35030 91366 35076 91418
rect 35100 91366 35146 91418
rect 35146 91366 35156 91418
rect 35180 91366 35210 91418
rect 35210 91366 35236 91418
rect 34940 91364 34996 91366
rect 35020 91364 35076 91366
rect 35100 91364 35156 91366
rect 35180 91364 35236 91366
rect 34940 90330 34996 90332
rect 35020 90330 35076 90332
rect 35100 90330 35156 90332
rect 35180 90330 35236 90332
rect 34940 90278 34966 90330
rect 34966 90278 34996 90330
rect 35020 90278 35030 90330
rect 35030 90278 35076 90330
rect 35100 90278 35146 90330
rect 35146 90278 35156 90330
rect 35180 90278 35210 90330
rect 35210 90278 35236 90330
rect 34940 90276 34996 90278
rect 35020 90276 35076 90278
rect 35100 90276 35156 90278
rect 35180 90276 35236 90278
rect 34940 89242 34996 89244
rect 35020 89242 35076 89244
rect 35100 89242 35156 89244
rect 35180 89242 35236 89244
rect 34940 89190 34966 89242
rect 34966 89190 34996 89242
rect 35020 89190 35030 89242
rect 35030 89190 35076 89242
rect 35100 89190 35146 89242
rect 35146 89190 35156 89242
rect 35180 89190 35210 89242
rect 35210 89190 35236 89242
rect 34940 89188 34996 89190
rect 35020 89188 35076 89190
rect 35100 89188 35156 89190
rect 35180 89188 35236 89190
rect 34940 88154 34996 88156
rect 35020 88154 35076 88156
rect 35100 88154 35156 88156
rect 35180 88154 35236 88156
rect 34940 88102 34966 88154
rect 34966 88102 34996 88154
rect 35020 88102 35030 88154
rect 35030 88102 35076 88154
rect 35100 88102 35146 88154
rect 35146 88102 35156 88154
rect 35180 88102 35210 88154
rect 35210 88102 35236 88154
rect 34940 88100 34996 88102
rect 35020 88100 35076 88102
rect 35100 88100 35156 88102
rect 35180 88100 35236 88102
rect 35346 114008 35402 114064
rect 35346 87216 35402 87272
rect 34940 87066 34996 87068
rect 35020 87066 35076 87068
rect 35100 87066 35156 87068
rect 35180 87066 35236 87068
rect 34940 87014 34966 87066
rect 34966 87014 34996 87066
rect 35020 87014 35030 87066
rect 35030 87014 35076 87066
rect 35100 87014 35146 87066
rect 35146 87014 35156 87066
rect 35180 87014 35210 87066
rect 35210 87014 35236 87066
rect 34940 87012 34996 87014
rect 35020 87012 35076 87014
rect 35100 87012 35156 87014
rect 35180 87012 35236 87014
rect 34940 85978 34996 85980
rect 35020 85978 35076 85980
rect 35100 85978 35156 85980
rect 35180 85978 35236 85980
rect 34940 85926 34966 85978
rect 34966 85926 34996 85978
rect 35020 85926 35030 85978
rect 35030 85926 35076 85978
rect 35100 85926 35146 85978
rect 35146 85926 35156 85978
rect 35180 85926 35210 85978
rect 35210 85926 35236 85978
rect 34940 85924 34996 85926
rect 35020 85924 35076 85926
rect 35100 85924 35156 85926
rect 35180 85924 35236 85926
rect 34940 84890 34996 84892
rect 35020 84890 35076 84892
rect 35100 84890 35156 84892
rect 35180 84890 35236 84892
rect 34940 84838 34966 84890
rect 34966 84838 34996 84890
rect 35020 84838 35030 84890
rect 35030 84838 35076 84890
rect 35100 84838 35146 84890
rect 35146 84838 35156 84890
rect 35180 84838 35210 84890
rect 35210 84838 35236 84890
rect 34940 84836 34996 84838
rect 35020 84836 35076 84838
rect 35100 84836 35156 84838
rect 35180 84836 35236 84838
rect 34940 83802 34996 83804
rect 35020 83802 35076 83804
rect 35100 83802 35156 83804
rect 35180 83802 35236 83804
rect 34940 83750 34966 83802
rect 34966 83750 34996 83802
rect 35020 83750 35030 83802
rect 35030 83750 35076 83802
rect 35100 83750 35146 83802
rect 35146 83750 35156 83802
rect 35180 83750 35210 83802
rect 35210 83750 35236 83802
rect 34940 83748 34996 83750
rect 35020 83748 35076 83750
rect 35100 83748 35156 83750
rect 35180 83748 35236 83750
rect 34940 82714 34996 82716
rect 35020 82714 35076 82716
rect 35100 82714 35156 82716
rect 35180 82714 35236 82716
rect 34940 82662 34966 82714
rect 34966 82662 34996 82714
rect 35020 82662 35030 82714
rect 35030 82662 35076 82714
rect 35100 82662 35146 82714
rect 35146 82662 35156 82714
rect 35180 82662 35210 82714
rect 35210 82662 35236 82714
rect 34940 82660 34996 82662
rect 35020 82660 35076 82662
rect 35100 82660 35156 82662
rect 35180 82660 35236 82662
rect 34940 81626 34996 81628
rect 35020 81626 35076 81628
rect 35100 81626 35156 81628
rect 35180 81626 35236 81628
rect 34940 81574 34966 81626
rect 34966 81574 34996 81626
rect 35020 81574 35030 81626
rect 35030 81574 35076 81626
rect 35100 81574 35146 81626
rect 35146 81574 35156 81626
rect 35180 81574 35210 81626
rect 35210 81574 35236 81626
rect 34940 81572 34996 81574
rect 35020 81572 35076 81574
rect 35100 81572 35156 81574
rect 35180 81572 35236 81574
rect 34940 80538 34996 80540
rect 35020 80538 35076 80540
rect 35100 80538 35156 80540
rect 35180 80538 35236 80540
rect 34940 80486 34966 80538
rect 34966 80486 34996 80538
rect 35020 80486 35030 80538
rect 35030 80486 35076 80538
rect 35100 80486 35146 80538
rect 35146 80486 35156 80538
rect 35180 80486 35210 80538
rect 35210 80486 35236 80538
rect 34940 80484 34996 80486
rect 35020 80484 35076 80486
rect 35100 80484 35156 80486
rect 35180 80484 35236 80486
rect 34940 79450 34996 79452
rect 35020 79450 35076 79452
rect 35100 79450 35156 79452
rect 35180 79450 35236 79452
rect 34940 79398 34966 79450
rect 34966 79398 34996 79450
rect 35020 79398 35030 79450
rect 35030 79398 35076 79450
rect 35100 79398 35146 79450
rect 35146 79398 35156 79450
rect 35180 79398 35210 79450
rect 35210 79398 35236 79450
rect 34940 79396 34996 79398
rect 35020 79396 35076 79398
rect 35100 79396 35156 79398
rect 35180 79396 35236 79398
rect 34940 78362 34996 78364
rect 35020 78362 35076 78364
rect 35100 78362 35156 78364
rect 35180 78362 35236 78364
rect 34940 78310 34966 78362
rect 34966 78310 34996 78362
rect 35020 78310 35030 78362
rect 35030 78310 35076 78362
rect 35100 78310 35146 78362
rect 35146 78310 35156 78362
rect 35180 78310 35210 78362
rect 35210 78310 35236 78362
rect 34940 78308 34996 78310
rect 35020 78308 35076 78310
rect 35100 78308 35156 78310
rect 35180 78308 35236 78310
rect 34940 77274 34996 77276
rect 35020 77274 35076 77276
rect 35100 77274 35156 77276
rect 35180 77274 35236 77276
rect 34940 77222 34966 77274
rect 34966 77222 34996 77274
rect 35020 77222 35030 77274
rect 35030 77222 35076 77274
rect 35100 77222 35146 77274
rect 35146 77222 35156 77274
rect 35180 77222 35210 77274
rect 35210 77222 35236 77274
rect 34940 77220 34996 77222
rect 35020 77220 35076 77222
rect 35100 77220 35156 77222
rect 35180 77220 35236 77222
rect 34940 76186 34996 76188
rect 35020 76186 35076 76188
rect 35100 76186 35156 76188
rect 35180 76186 35236 76188
rect 34940 76134 34966 76186
rect 34966 76134 34996 76186
rect 35020 76134 35030 76186
rect 35030 76134 35076 76186
rect 35100 76134 35146 76186
rect 35146 76134 35156 76186
rect 35180 76134 35210 76186
rect 35210 76134 35236 76186
rect 34940 76132 34996 76134
rect 35020 76132 35076 76134
rect 35100 76132 35156 76134
rect 35180 76132 35236 76134
rect 34940 75098 34996 75100
rect 35020 75098 35076 75100
rect 35100 75098 35156 75100
rect 35180 75098 35236 75100
rect 34940 75046 34966 75098
rect 34966 75046 34996 75098
rect 35020 75046 35030 75098
rect 35030 75046 35076 75098
rect 35100 75046 35146 75098
rect 35146 75046 35156 75098
rect 35180 75046 35210 75098
rect 35210 75046 35236 75098
rect 34940 75044 34996 75046
rect 35020 75044 35076 75046
rect 35100 75044 35156 75046
rect 35180 75044 35236 75046
rect 34940 74010 34996 74012
rect 35020 74010 35076 74012
rect 35100 74010 35156 74012
rect 35180 74010 35236 74012
rect 34940 73958 34966 74010
rect 34966 73958 34996 74010
rect 35020 73958 35030 74010
rect 35030 73958 35076 74010
rect 35100 73958 35146 74010
rect 35146 73958 35156 74010
rect 35180 73958 35210 74010
rect 35210 73958 35236 74010
rect 34940 73956 34996 73958
rect 35020 73956 35076 73958
rect 35100 73956 35156 73958
rect 35180 73956 35236 73958
rect 34940 72922 34996 72924
rect 35020 72922 35076 72924
rect 35100 72922 35156 72924
rect 35180 72922 35236 72924
rect 34940 72870 34966 72922
rect 34966 72870 34996 72922
rect 35020 72870 35030 72922
rect 35030 72870 35076 72922
rect 35100 72870 35146 72922
rect 35146 72870 35156 72922
rect 35180 72870 35210 72922
rect 35210 72870 35236 72922
rect 34940 72868 34996 72870
rect 35020 72868 35076 72870
rect 35100 72868 35156 72870
rect 35180 72868 35236 72870
rect 34940 71834 34996 71836
rect 35020 71834 35076 71836
rect 35100 71834 35156 71836
rect 35180 71834 35236 71836
rect 34940 71782 34966 71834
rect 34966 71782 34996 71834
rect 35020 71782 35030 71834
rect 35030 71782 35076 71834
rect 35100 71782 35146 71834
rect 35146 71782 35156 71834
rect 35180 71782 35210 71834
rect 35210 71782 35236 71834
rect 34940 71780 34996 71782
rect 35020 71780 35076 71782
rect 35100 71780 35156 71782
rect 35180 71780 35236 71782
rect 34940 70746 34996 70748
rect 35020 70746 35076 70748
rect 35100 70746 35156 70748
rect 35180 70746 35236 70748
rect 34940 70694 34966 70746
rect 34966 70694 34996 70746
rect 35020 70694 35030 70746
rect 35030 70694 35076 70746
rect 35100 70694 35146 70746
rect 35146 70694 35156 70746
rect 35180 70694 35210 70746
rect 35210 70694 35236 70746
rect 34940 70692 34996 70694
rect 35020 70692 35076 70694
rect 35100 70692 35156 70694
rect 35180 70692 35236 70694
rect 34940 69658 34996 69660
rect 35020 69658 35076 69660
rect 35100 69658 35156 69660
rect 35180 69658 35236 69660
rect 34940 69606 34966 69658
rect 34966 69606 34996 69658
rect 35020 69606 35030 69658
rect 35030 69606 35076 69658
rect 35100 69606 35146 69658
rect 35146 69606 35156 69658
rect 35180 69606 35210 69658
rect 35210 69606 35236 69658
rect 34940 69604 34996 69606
rect 35020 69604 35076 69606
rect 35100 69604 35156 69606
rect 35180 69604 35236 69606
rect 34940 68570 34996 68572
rect 35020 68570 35076 68572
rect 35100 68570 35156 68572
rect 35180 68570 35236 68572
rect 34940 68518 34966 68570
rect 34966 68518 34996 68570
rect 35020 68518 35030 68570
rect 35030 68518 35076 68570
rect 35100 68518 35146 68570
rect 35146 68518 35156 68570
rect 35180 68518 35210 68570
rect 35210 68518 35236 68570
rect 34940 68516 34996 68518
rect 35020 68516 35076 68518
rect 35100 68516 35156 68518
rect 35180 68516 35236 68518
rect 34940 67482 34996 67484
rect 35020 67482 35076 67484
rect 35100 67482 35156 67484
rect 35180 67482 35236 67484
rect 34940 67430 34966 67482
rect 34966 67430 34996 67482
rect 35020 67430 35030 67482
rect 35030 67430 35076 67482
rect 35100 67430 35146 67482
rect 35146 67430 35156 67482
rect 35180 67430 35210 67482
rect 35210 67430 35236 67482
rect 34940 67428 34996 67430
rect 35020 67428 35076 67430
rect 35100 67428 35156 67430
rect 35180 67428 35236 67430
rect 34940 66394 34996 66396
rect 35020 66394 35076 66396
rect 35100 66394 35156 66396
rect 35180 66394 35236 66396
rect 34940 66342 34966 66394
rect 34966 66342 34996 66394
rect 35020 66342 35030 66394
rect 35030 66342 35076 66394
rect 35100 66342 35146 66394
rect 35146 66342 35156 66394
rect 35180 66342 35210 66394
rect 35210 66342 35236 66394
rect 34940 66340 34996 66342
rect 35020 66340 35076 66342
rect 35100 66340 35156 66342
rect 35180 66340 35236 66342
rect 34940 65306 34996 65308
rect 35020 65306 35076 65308
rect 35100 65306 35156 65308
rect 35180 65306 35236 65308
rect 34940 65254 34966 65306
rect 34966 65254 34996 65306
rect 35020 65254 35030 65306
rect 35030 65254 35076 65306
rect 35100 65254 35146 65306
rect 35146 65254 35156 65306
rect 35180 65254 35210 65306
rect 35210 65254 35236 65306
rect 34940 65252 34996 65254
rect 35020 65252 35076 65254
rect 35100 65252 35156 65254
rect 35180 65252 35236 65254
rect 34940 64218 34996 64220
rect 35020 64218 35076 64220
rect 35100 64218 35156 64220
rect 35180 64218 35236 64220
rect 34940 64166 34966 64218
rect 34966 64166 34996 64218
rect 35020 64166 35030 64218
rect 35030 64166 35076 64218
rect 35100 64166 35146 64218
rect 35146 64166 35156 64218
rect 35180 64166 35210 64218
rect 35210 64166 35236 64218
rect 34940 64164 34996 64166
rect 35020 64164 35076 64166
rect 35100 64164 35156 64166
rect 35180 64164 35236 64166
rect 34940 63130 34996 63132
rect 35020 63130 35076 63132
rect 35100 63130 35156 63132
rect 35180 63130 35236 63132
rect 34940 63078 34966 63130
rect 34966 63078 34996 63130
rect 35020 63078 35030 63130
rect 35030 63078 35076 63130
rect 35100 63078 35146 63130
rect 35146 63078 35156 63130
rect 35180 63078 35210 63130
rect 35210 63078 35236 63130
rect 34940 63076 34996 63078
rect 35020 63076 35076 63078
rect 35100 63076 35156 63078
rect 35180 63076 35236 63078
rect 35438 86944 35494 87000
rect 35806 113600 35862 113656
rect 35622 87488 35678 87544
rect 35622 86944 35678 87000
rect 34940 62042 34996 62044
rect 35020 62042 35076 62044
rect 35100 62042 35156 62044
rect 35180 62042 35236 62044
rect 34940 61990 34966 62042
rect 34966 61990 34996 62042
rect 35020 61990 35030 62042
rect 35030 61990 35076 62042
rect 35100 61990 35146 62042
rect 35146 61990 35156 62042
rect 35180 61990 35210 62042
rect 35210 61990 35236 62042
rect 34940 61988 34996 61990
rect 35020 61988 35076 61990
rect 35100 61988 35156 61990
rect 35180 61988 35236 61990
rect 34518 44940 34574 44976
rect 34518 44920 34520 44940
rect 34520 44920 34572 44940
rect 34572 44920 34574 44940
rect 34610 41112 34666 41168
rect 34610 39752 34666 39808
rect 34518 39344 34574 39400
rect 34610 34584 34666 34640
rect 34940 60954 34996 60956
rect 35020 60954 35076 60956
rect 35100 60954 35156 60956
rect 35180 60954 35236 60956
rect 34940 60902 34966 60954
rect 34966 60902 34996 60954
rect 35020 60902 35030 60954
rect 35030 60902 35076 60954
rect 35100 60902 35146 60954
rect 35146 60902 35156 60954
rect 35180 60902 35210 60954
rect 35210 60902 35236 60954
rect 34940 60900 34996 60902
rect 35020 60900 35076 60902
rect 35100 60900 35156 60902
rect 35180 60900 35236 60902
rect 34940 59866 34996 59868
rect 35020 59866 35076 59868
rect 35100 59866 35156 59868
rect 35180 59866 35236 59868
rect 34940 59814 34966 59866
rect 34966 59814 34996 59866
rect 35020 59814 35030 59866
rect 35030 59814 35076 59866
rect 35100 59814 35146 59866
rect 35146 59814 35156 59866
rect 35180 59814 35210 59866
rect 35210 59814 35236 59866
rect 34940 59812 34996 59814
rect 35020 59812 35076 59814
rect 35100 59812 35156 59814
rect 35180 59812 35236 59814
rect 34940 58778 34996 58780
rect 35020 58778 35076 58780
rect 35100 58778 35156 58780
rect 35180 58778 35236 58780
rect 34940 58726 34966 58778
rect 34966 58726 34996 58778
rect 35020 58726 35030 58778
rect 35030 58726 35076 58778
rect 35100 58726 35146 58778
rect 35146 58726 35156 58778
rect 35180 58726 35210 58778
rect 35210 58726 35236 58778
rect 34940 58724 34996 58726
rect 35020 58724 35076 58726
rect 35100 58724 35156 58726
rect 35180 58724 35236 58726
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 34886 55820 34942 55856
rect 34886 55800 34888 55820
rect 34888 55800 34940 55820
rect 34940 55800 34942 55820
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 35438 55392 35494 55448
rect 36634 119176 36690 119232
rect 36542 117136 36598 117192
rect 36542 111444 36598 111480
rect 36542 111424 36544 111444
rect 36544 111424 36596 111444
rect 36596 111424 36598 111444
rect 35806 54848 35862 54904
rect 35714 54032 35770 54088
rect 35806 52808 35862 52864
rect 35806 50224 35862 50280
rect 35530 48864 35586 48920
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 35254 46280 35310 46336
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 35070 43696 35126 43752
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34978 43288 35034 43344
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34794 41928 34850 41984
rect 34794 41520 34850 41576
rect 35346 44512 35402 44568
rect 35346 43968 35402 44024
rect 35346 42336 35402 42392
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 35162 40704 35218 40760
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34794 38528 34850 38584
rect 34978 38936 35034 38992
rect 35898 47640 35954 47696
rect 35806 47540 35808 47560
rect 35808 47540 35860 47560
rect 35860 47540 35862 47560
rect 35806 47504 35862 47540
rect 35806 47116 35862 47152
rect 35806 47096 35808 47116
rect 35808 47096 35860 47116
rect 35860 47096 35862 47116
rect 35714 45872 35770 45928
rect 35714 45736 35770 45792
rect 35806 45464 35862 45520
rect 35806 45364 35808 45384
rect 35808 45364 35860 45384
rect 35860 45364 35862 45384
rect 35806 45328 35862 45364
rect 35714 45192 35770 45248
rect 35806 44648 35862 44704
rect 36818 117408 36874 117464
rect 36726 114824 36782 114880
rect 37002 118360 37058 118416
rect 37094 117000 37150 117056
rect 37186 115776 37242 115832
rect 37094 114416 37150 114472
rect 37646 116592 37702 116648
rect 37830 116048 37886 116104
rect 37646 115368 37702 115424
rect 37186 110220 37242 110256
rect 37186 110200 37188 110220
rect 37188 110200 37240 110220
rect 37240 110200 37242 110220
rect 37186 109656 37242 109712
rect 37370 114028 37426 114064
rect 37370 114008 37372 114028
rect 37372 114008 37424 114028
rect 37424 114008 37426 114028
rect 37370 113192 37426 113248
rect 37370 112804 37426 112840
rect 37370 112784 37372 112804
rect 37372 112784 37424 112804
rect 37424 112784 37426 112804
rect 37646 111832 37702 111888
rect 37370 111016 37426 111072
rect 37462 110644 37464 110664
rect 37464 110644 37516 110664
rect 37516 110644 37518 110664
rect 37462 110608 37518 110644
rect 38106 112240 38162 112296
rect 37186 108840 37242 108896
rect 37186 108044 37242 108080
rect 37186 108024 37188 108044
rect 37188 108024 37240 108044
rect 37240 108024 37242 108044
rect 37186 107480 37242 107536
rect 37186 106664 37242 106720
rect 37278 106292 37280 106312
rect 37280 106292 37332 106312
rect 37332 106292 37334 106312
rect 37278 106256 37334 106292
rect 37186 105868 37242 105904
rect 37186 105848 37188 105868
rect 37188 105848 37240 105868
rect 37240 105848 37242 105868
rect 37186 105440 37242 105496
rect 37186 104488 37242 104544
rect 37186 104100 37242 104136
rect 37186 104080 37188 104100
rect 37188 104080 37240 104100
rect 37240 104080 37242 104100
rect 37186 103264 37242 103320
rect 37278 102856 37334 102912
rect 37186 102312 37242 102368
rect 37186 101516 37242 101552
rect 37186 101496 37188 101516
rect 37188 101496 37240 101516
rect 37240 101496 37242 101516
rect 37186 100680 37242 100736
rect 37186 100272 37242 100328
rect 37186 99340 37242 99376
rect 37186 99320 37188 99340
rect 37188 99320 37240 99340
rect 37240 99320 37242 99340
rect 37186 98912 37242 98968
rect 37186 98096 37242 98152
rect 37186 97164 37242 97200
rect 37186 97144 37188 97164
rect 37188 97144 37240 97164
rect 37240 97144 37242 97164
rect 37186 96328 37242 96384
rect 37186 95920 37242 95976
rect 37278 95512 37334 95568
rect 37186 94988 37242 95024
rect 37186 94968 37188 94988
rect 37188 94968 37240 94988
rect 37240 94968 37242 94988
rect 37922 109248 37978 109304
rect 37922 108452 37978 108488
rect 37922 108432 37924 108452
rect 37924 108432 37976 108452
rect 37976 108432 37978 108452
rect 37922 107072 37978 107128
rect 37922 104896 37978 104952
rect 37922 103672 37978 103728
rect 37922 101924 37978 101960
rect 37922 101904 37924 101924
rect 37924 101904 37976 101924
rect 37976 101904 37978 101924
rect 37922 101088 37978 101144
rect 37922 99748 37978 99784
rect 37922 99728 37924 99748
rect 37924 99728 37976 99748
rect 37976 99728 37978 99748
rect 37278 94152 37334 94208
rect 37278 93336 37334 93392
rect 37186 92928 37242 92984
rect 37278 91976 37334 92032
rect 37278 91160 37334 91216
rect 37186 90752 37242 90808
rect 37278 89800 37334 89856
rect 37278 88984 37334 89040
rect 37186 88576 37242 88632
rect 37278 87796 37280 87816
rect 37280 87796 37332 87816
rect 37332 87796 37334 87816
rect 37278 87760 37334 87796
rect 37278 86808 37334 86864
rect 37186 86400 37242 86456
rect 37278 85620 37280 85640
rect 37280 85620 37332 85640
rect 37332 85620 37334 85640
rect 37278 85584 37334 85620
rect 37278 84632 37334 84688
rect 37186 84224 37242 84280
rect 37278 83444 37280 83464
rect 37280 83444 37332 83464
rect 37332 83444 37334 83464
rect 37278 83408 37334 83444
rect 37278 82456 37334 82512
rect 37186 82048 37242 82104
rect 36082 45620 36138 45656
rect 36082 45600 36084 45620
rect 36084 45600 36136 45620
rect 36136 45600 36138 45620
rect 36082 45056 36138 45112
rect 35898 44240 35954 44296
rect 35806 44104 35862 44160
rect 35714 42880 35770 42936
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34794 36080 34850 36136
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35346 38120 35402 38176
rect 35530 38936 35586 38992
rect 35806 40296 35862 40352
rect 35714 38936 35770 38992
rect 35530 37168 35586 37224
rect 35438 36352 35494 36408
rect 34794 35572 34796 35592
rect 34796 35572 34848 35592
rect 34848 35572 34850 35592
rect 34794 35536 34850 35572
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34426 2760 34482 2816
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 35530 35672 35586 35728
rect 36450 58792 36506 58848
rect 36450 57996 36506 58032
rect 36450 57976 36452 57996
rect 36452 57976 36504 57996
rect 36504 57976 36506 57996
rect 36450 57024 36506 57080
rect 36910 59200 36966 59256
rect 37278 81268 37280 81288
rect 37280 81268 37332 81288
rect 37332 81268 37334 81288
rect 37278 81232 37334 81268
rect 37278 80416 37334 80472
rect 37186 79872 37242 79928
rect 37922 98504 37978 98560
rect 37922 97688 37978 97744
rect 37922 96736 37978 96792
rect 37922 94560 37978 94616
rect 37922 93744 37978 93800
rect 37922 91568 37978 91624
rect 37922 90344 37978 90400
rect 37922 89392 37978 89448
rect 37922 88168 37978 88224
rect 37922 87216 37978 87272
rect 38014 86536 38070 86592
rect 37922 85992 37978 86048
rect 37922 85176 37978 85232
rect 37186 78684 37188 78704
rect 37188 78684 37240 78704
rect 37240 78684 37242 78704
rect 37186 78648 37242 78684
rect 37186 78240 37242 78296
rect 37186 77288 37242 77344
rect 37186 76492 37242 76528
rect 37186 76472 37188 76492
rect 37188 76472 37240 76492
rect 37240 76472 37242 76492
rect 37186 76064 37242 76120
rect 37186 75248 37242 75304
rect 37186 74316 37242 74352
rect 37186 74296 37188 74316
rect 37188 74296 37240 74316
rect 37240 74296 37242 74316
rect 37186 73888 37242 73944
rect 37186 73072 37242 73128
rect 37002 56208 37058 56264
rect 37186 72140 37242 72176
rect 37186 72120 37188 72140
rect 37188 72120 37240 72140
rect 37240 72120 37242 72140
rect 37186 71712 37242 71768
rect 37186 70896 37242 70952
rect 37186 69964 37242 70000
rect 37186 69944 37188 69964
rect 37188 69944 37240 69964
rect 37240 69944 37242 69964
rect 37186 69536 37242 69592
rect 37186 68720 37242 68776
rect 37278 68312 37334 68368
rect 37186 67904 37242 67960
rect 37278 66952 37334 67008
rect 37278 66136 37334 66192
rect 37186 65728 37242 65784
rect 37186 64776 37242 64832
rect 37278 63960 37334 64016
rect 37186 63552 37242 63608
rect 37278 62772 37280 62792
rect 37280 62772 37332 62792
rect 37332 62772 37334 62792
rect 37278 62736 37334 62772
rect 37278 61784 37334 61840
rect 37186 61376 37242 61432
rect 37278 60596 37280 60616
rect 37280 60596 37332 60616
rect 37332 60596 37334 60616
rect 37278 60560 37334 60596
rect 37186 60172 37242 60208
rect 37186 60152 37188 60172
rect 37188 60152 37240 60172
rect 37240 60152 37242 60172
rect 37186 58384 37242 58440
rect 37186 57432 37242 57488
rect 37186 56616 37242 56672
rect 36726 53644 36782 53680
rect 36726 53624 36728 53644
rect 36728 53624 36780 53644
rect 36780 53624 36782 53644
rect 36726 52964 36782 53000
rect 36726 52944 36728 52964
rect 36728 52944 36780 52964
rect 36780 52944 36782 52964
rect 36266 49716 36268 49736
rect 36268 49716 36320 49736
rect 36320 49716 36322 49736
rect 36266 49680 36322 49716
rect 36266 48728 36322 48784
rect 36266 48456 36322 48512
rect 36542 51468 36598 51504
rect 36542 51448 36544 51468
rect 36544 51448 36596 51468
rect 36596 51448 36598 51468
rect 36726 52264 36782 52320
rect 37094 54440 37150 54496
rect 36358 48048 36414 48104
rect 36358 46688 36414 46744
rect 36450 44240 36506 44296
rect 36542 43988 36598 44024
rect 36542 43968 36544 43988
rect 36544 43968 36596 43988
rect 36596 43968 36598 43988
rect 36174 40976 36230 41032
rect 36082 39924 36084 39944
rect 36084 39924 36136 39944
rect 36136 39924 36138 39944
rect 36082 39888 36138 39924
rect 36082 39616 36138 39672
rect 36174 37748 36176 37768
rect 36176 37748 36228 37768
rect 36228 37748 36230 37768
rect 36174 37712 36230 37748
rect 36174 37032 36230 37088
rect 35530 34720 35586 34776
rect 35622 34176 35678 34232
rect 35530 34076 35532 34096
rect 35532 34076 35584 34096
rect 35584 34076 35586 34096
rect 35530 34040 35586 34076
rect 35898 36236 35954 36272
rect 35898 36216 35900 36236
rect 35900 36216 35952 36236
rect 35952 36216 35954 36236
rect 35438 33360 35494 33416
rect 35530 32000 35586 32056
rect 35898 34448 35954 34504
rect 35898 33632 35954 33688
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 35806 30796 35862 30832
rect 35806 30776 35808 30796
rect 35808 30776 35860 30796
rect 35860 30776 35862 30796
rect 35806 29416 35862 29472
rect 36358 36760 36414 36816
rect 37186 51856 37242 51912
rect 37462 62464 37518 62520
rect 37922 83816 37978 83872
rect 37922 83000 37978 83056
rect 37922 81640 37978 81696
rect 37922 80824 37978 80880
rect 37922 79464 37978 79520
rect 37922 79092 37924 79112
rect 37924 79092 37976 79112
rect 37976 79092 37978 79112
rect 37922 79056 37978 79092
rect 37922 77832 37978 77888
rect 37922 76900 37978 76936
rect 37922 76880 37924 76900
rect 37924 76880 37976 76900
rect 37976 76880 37978 76900
rect 38750 86672 38806 86728
rect 38934 92384 38990 92440
rect 38842 80280 38898 80336
rect 37922 75656 37978 75712
rect 37922 74724 37978 74760
rect 37922 74704 37924 74724
rect 37924 74704 37976 74724
rect 37976 74704 37978 74724
rect 37922 73480 37978 73536
rect 37922 72664 37978 72720
rect 37370 53216 37426 53272
rect 37370 51040 37426 51096
rect 36818 43832 36874 43888
rect 37186 45736 37242 45792
rect 37186 44396 37242 44432
rect 37186 44376 37188 44396
rect 37188 44376 37240 44396
rect 37240 44376 37242 44396
rect 37370 45056 37426 45112
rect 36542 39072 36598 39128
rect 36450 35808 36506 35864
rect 36358 35672 36414 35728
rect 36174 34720 36230 34776
rect 36174 34448 36230 34504
rect 36082 33088 36138 33144
rect 35990 30232 36046 30288
rect 36174 31184 36230 31240
rect 36634 36216 36690 36272
rect 37094 40976 37150 41032
rect 36910 40024 36966 40080
rect 36910 39616 36966 39672
rect 36910 39480 36966 39536
rect 36910 38412 36966 38448
rect 36910 38392 36912 38412
rect 36912 38392 36964 38412
rect 36964 38392 36966 38412
rect 36910 38004 36966 38040
rect 36910 37984 36912 38004
rect 36912 37984 36964 38004
rect 36964 37984 36966 38004
rect 36726 34060 36782 34096
rect 36726 34040 36728 34060
rect 36728 34040 36780 34060
rect 36780 34040 36782 34060
rect 36634 33632 36690 33688
rect 35898 28952 35954 29008
rect 36082 29008 36138 29064
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 36358 28736 36414 28792
rect 36726 30368 36782 30424
rect 37554 43832 37610 43888
rect 37278 38800 37334 38856
rect 37370 36488 37426 36544
rect 37462 35808 37518 35864
rect 37462 34992 37518 35048
rect 37370 33768 37426 33824
rect 37370 32972 37426 33008
rect 37370 32952 37372 32972
rect 37372 32952 37424 32972
rect 37424 32952 37426 32972
rect 36910 31592 36966 31648
rect 35806 3576 35862 3632
rect 37186 29144 37242 29200
rect 37186 28192 37242 28248
rect 37462 30232 37518 30288
rect 37370 29824 37426 29880
rect 37922 71304 37978 71360
rect 37922 70488 37978 70544
rect 37922 69128 37978 69184
rect 37922 66544 37978 66600
rect 37922 65320 37978 65376
rect 37922 64368 37978 64424
rect 37922 63144 37978 63200
rect 37922 62192 37978 62248
rect 37922 60968 37978 61024
rect 37922 59608 37978 59664
rect 37738 52980 37740 53000
rect 37740 52980 37792 53000
rect 37792 52980 37794 53000
rect 37738 52944 37794 52980
rect 38106 50632 38162 50688
rect 38106 49272 38162 49328
rect 37738 45328 37794 45384
rect 37738 45228 37740 45248
rect 37740 45228 37792 45248
rect 37792 45228 37794 45248
rect 37738 45192 37794 45228
rect 37738 38392 37794 38448
rect 38106 45600 38162 45656
rect 38014 44648 38070 44704
rect 38106 43152 38162 43208
rect 38106 39924 38108 39944
rect 38108 39924 38160 39944
rect 38160 39924 38162 39944
rect 38106 39888 38162 39924
rect 38106 38664 38162 38720
rect 37922 37984 37978 38040
rect 37462 29044 37464 29064
rect 37464 29044 37516 29064
rect 37516 29044 37518 29064
rect 37462 29008 37518 29044
rect 37370 28600 37426 28656
rect 37462 27784 37518 27840
rect 37278 26868 37280 26888
rect 37280 26868 37332 26888
rect 37332 26868 37334 26888
rect 37278 26832 37334 26868
rect 37278 25608 37334 25664
rect 37186 25200 37242 25256
rect 37186 24268 37242 24304
rect 37186 24248 37188 24268
rect 37188 24248 37240 24268
rect 37240 24248 37242 24268
rect 37462 23840 37518 23896
rect 37186 23024 37242 23080
rect 37278 22516 37280 22536
rect 37280 22516 37332 22536
rect 37332 22516 37334 22536
rect 37278 22480 37334 22516
rect 37186 21664 37242 21720
rect 37278 21256 37334 21312
rect 37278 20440 37334 20496
rect 37278 19080 37334 19136
rect 37186 18672 37242 18728
rect 37186 17856 37242 17912
rect 37278 17312 37334 17368
rect 37186 16496 37242 16552
rect 37278 16088 37334 16144
rect 37186 15272 37242 15328
rect 37278 14728 37334 14784
rect 37186 13912 37242 13968
rect 37186 13096 37242 13152
rect 37186 12144 37242 12200
rect 37186 11736 37242 11792
rect 37186 10920 37242 10976
rect 37186 9968 37242 10024
rect 37186 9560 37242 9616
rect 37186 8744 37242 8800
rect 37186 7948 37242 7984
rect 37186 7928 37188 7948
rect 37188 7928 37240 7948
rect 37240 7928 37242 7948
rect 37186 7384 37242 7440
rect 37186 6568 37242 6624
rect 36634 3168 36690 3224
rect 36542 2760 36598 2816
rect 36450 2216 36506 2272
rect 2778 448 2834 504
rect 36818 1808 36874 1864
rect 37186 5772 37242 5808
rect 37186 5752 37188 5772
rect 37188 5752 37240 5772
rect 37240 5752 37242 5772
rect 37186 5344 37242 5400
rect 37186 4392 37242 4448
rect 37094 3984 37150 4040
rect 38106 33088 38162 33144
rect 38014 32408 38070 32464
rect 37830 28872 37886 28928
rect 37922 27240 37978 27296
rect 37922 26424 37978 26480
rect 37922 26016 37978 26072
rect 37922 24692 37924 24712
rect 37924 24692 37976 24712
rect 37976 24692 37978 24712
rect 37922 24656 37978 24692
rect 38106 28600 38162 28656
rect 38106 23432 38162 23488
rect 37922 22072 37978 22128
rect 37922 20848 37978 20904
rect 37922 19896 37978 19952
rect 37922 19488 37978 19544
rect 38934 67360 38990 67416
rect 38566 38256 38622 38312
rect 37922 18264 37978 18320
rect 37922 16904 37978 16960
rect 37922 15680 37978 15736
rect 37922 14320 37978 14376
rect 37922 13504 37978 13560
rect 37922 12708 37978 12744
rect 37922 12688 37924 12708
rect 37924 12688 37976 12708
rect 37976 12688 37978 12708
rect 37922 11328 37978 11384
rect 37922 10532 37978 10568
rect 37922 10512 37924 10532
rect 37924 10512 37976 10532
rect 37976 10512 37978 10532
rect 37922 9152 37978 9208
rect 37922 8356 37978 8392
rect 37922 8336 37924 8356
rect 37924 8336 37976 8356
rect 37976 8336 37978 8356
rect 37922 6976 37978 7032
rect 37922 6180 37978 6216
rect 37922 6160 37924 6180
rect 37924 6160 37976 6180
rect 37976 6160 37978 6180
rect 37922 4800 37978 4856
rect 37186 992 37242 1048
rect 36726 584 36782 640
rect 38106 1400 38162 1456
rect 37922 176 37978 232
<< metal3 >>
rect 36353 119642 36419 119645
rect 39200 119642 40800 119672
rect 36353 119640 40800 119642
rect 36353 119584 36358 119640
rect 36414 119584 40800 119640
rect 36353 119582 40800 119584
rect 36353 119579 36419 119582
rect 39200 119552 40800 119582
rect -800 119506 800 119536
rect 3325 119506 3391 119509
rect -800 119504 3391 119506
rect -800 119448 3330 119504
rect 3386 119448 3391 119504
rect -800 119446 3391 119448
rect -800 119416 800 119446
rect 3325 119443 3391 119446
rect 36629 119234 36695 119237
rect 39200 119234 40800 119264
rect 36629 119232 40800 119234
rect 36629 119176 36634 119232
rect 36690 119176 40800 119232
rect 36629 119174 40800 119176
rect 36629 119171 36695 119174
rect 39200 119144 40800 119174
rect 34697 118826 34763 118829
rect 39200 118826 40800 118856
rect 34697 118824 40800 118826
rect 34697 118768 34702 118824
rect 34758 118768 40800 118824
rect 34697 118766 40800 118768
rect 34697 118763 34763 118766
rect 39200 118736 40800 118766
rect -800 118690 800 118720
rect 3141 118690 3207 118693
rect -800 118688 3207 118690
rect -800 118632 3146 118688
rect 3202 118632 3207 118688
rect -800 118630 3207 118632
rect -800 118600 800 118630
rect 3141 118627 3207 118630
rect 36997 118418 37063 118421
rect 39200 118418 40800 118448
rect 36997 118416 40800 118418
rect 36997 118360 37002 118416
rect 37058 118360 40800 118416
rect 36997 118358 40800 118360
rect 36997 118355 37063 118358
rect 39200 118328 40800 118358
rect 34513 118010 34579 118013
rect 39200 118010 40800 118040
rect 34513 118008 40800 118010
rect 34513 117952 34518 118008
rect 34574 117952 40800 118008
rect 34513 117950 40800 117952
rect 34513 117947 34579 117950
rect 39200 117920 40800 117950
rect -800 117874 800 117904
rect 2957 117874 3023 117877
rect -800 117872 3023 117874
rect -800 117816 2962 117872
rect 3018 117816 3023 117872
rect -800 117814 3023 117816
rect -800 117784 800 117814
rect 2957 117811 3023 117814
rect 4208 117536 4528 117537
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 117471 4528 117472
rect 34928 117536 35248 117537
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 117471 35248 117472
rect 36813 117466 36879 117469
rect 39200 117466 40800 117496
rect 36813 117464 40800 117466
rect 36813 117408 36818 117464
rect 36874 117408 40800 117464
rect 36813 117406 40800 117408
rect 36813 117403 36879 117406
rect 39200 117376 40800 117406
rect 19885 117330 19951 117333
rect 23197 117330 23263 117333
rect 19885 117328 23263 117330
rect 19885 117272 19890 117328
rect 19946 117272 23202 117328
rect 23258 117272 23263 117328
rect 19885 117270 23263 117272
rect 19885 117267 19951 117270
rect 23197 117267 23263 117270
rect 22553 117194 22619 117197
rect 36537 117194 36603 117197
rect 22553 117192 36603 117194
rect 22553 117136 22558 117192
rect 22614 117136 36542 117192
rect 36598 117136 36603 117192
rect 22553 117134 36603 117136
rect 22553 117131 22619 117134
rect 36537 117131 36603 117134
rect -800 117058 800 117088
rect 2865 117058 2931 117061
rect -800 117056 2931 117058
rect -800 117000 2870 117056
rect 2926 117000 2931 117056
rect -800 116998 2931 117000
rect -800 116968 800 116998
rect 2865 116995 2931 116998
rect 23197 117058 23263 117061
rect 27153 117058 27219 117061
rect 23197 117056 27219 117058
rect 23197 117000 23202 117056
rect 23258 117000 27158 117056
rect 27214 117000 27219 117056
rect 23197 116998 27219 117000
rect 23197 116995 23263 116998
rect 27153 116995 27219 116998
rect 37089 117058 37155 117061
rect 39200 117058 40800 117088
rect 37089 117056 40800 117058
rect 37089 117000 37094 117056
rect 37150 117000 40800 117056
rect 37089 116998 40800 117000
rect 37089 116995 37155 116998
rect 19568 116992 19888 116993
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 39200 116968 40800 116998
rect 19568 116927 19888 116928
rect 25129 116922 25195 116925
rect 28349 116922 28415 116925
rect 25129 116920 28415 116922
rect 25129 116864 25134 116920
rect 25190 116864 28354 116920
rect 28410 116864 28415 116920
rect 25129 116862 28415 116864
rect 25129 116859 25195 116862
rect 28349 116859 28415 116862
rect 21449 116650 21515 116653
rect 22093 116650 22159 116653
rect 21449 116648 22159 116650
rect 21449 116592 21454 116648
rect 21510 116592 22098 116648
rect 22154 116592 22159 116648
rect 21449 116590 22159 116592
rect 21449 116587 21515 116590
rect 22093 116587 22159 116590
rect 37641 116650 37707 116653
rect 39200 116650 40800 116680
rect 37641 116648 40800 116650
rect 37641 116592 37646 116648
rect 37702 116592 40800 116648
rect 37641 116590 40800 116592
rect 37641 116587 37707 116590
rect 39200 116560 40800 116590
rect 4208 116448 4528 116449
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 116383 4528 116384
rect 34928 116448 35248 116449
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 34928 116383 35248 116384
rect -800 116242 800 116272
rect 1393 116242 1459 116245
rect -800 116240 1459 116242
rect -800 116184 1398 116240
rect 1454 116184 1459 116240
rect -800 116182 1459 116184
rect -800 116152 800 116182
rect 1393 116179 1459 116182
rect 21909 116242 21975 116245
rect 25497 116242 25563 116245
rect 30649 116242 30715 116245
rect 21909 116240 22110 116242
rect 21909 116184 21914 116240
rect 21970 116184 22110 116240
rect 21909 116182 22110 116184
rect 21909 116179 21975 116182
rect 22050 116106 22110 116182
rect 25497 116240 30715 116242
rect 25497 116184 25502 116240
rect 25558 116184 30654 116240
rect 30710 116184 30715 116240
rect 25497 116182 30715 116184
rect 25497 116179 25563 116182
rect 30649 116179 30715 116182
rect 35341 116242 35407 116245
rect 39200 116242 40800 116272
rect 35341 116240 40800 116242
rect 35341 116184 35346 116240
rect 35402 116184 40800 116240
rect 35341 116182 40800 116184
rect 35341 116179 35407 116182
rect 39200 116152 40800 116182
rect 37825 116106 37891 116109
rect 22050 116104 37891 116106
rect 22050 116048 37830 116104
rect 37886 116048 37891 116104
rect 22050 116046 37891 116048
rect 37825 116043 37891 116046
rect 24485 115970 24551 115973
rect 28257 115970 28323 115973
rect 24485 115968 28323 115970
rect 24485 115912 24490 115968
rect 24546 115912 28262 115968
rect 28318 115912 28323 115968
rect 24485 115910 28323 115912
rect 24485 115907 24551 115910
rect 28257 115907 28323 115910
rect 19568 115904 19888 115905
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 115839 19888 115840
rect 20253 115834 20319 115837
rect 23933 115834 23999 115837
rect 20253 115832 23999 115834
rect 20253 115776 20258 115832
rect 20314 115776 23938 115832
rect 23994 115776 23999 115832
rect 20253 115774 23999 115776
rect 20253 115771 20319 115774
rect 23933 115771 23999 115774
rect 37181 115834 37247 115837
rect 39200 115834 40800 115864
rect 37181 115832 40800 115834
rect 37181 115776 37186 115832
rect 37242 115776 40800 115832
rect 37181 115774 40800 115776
rect 37181 115771 37247 115774
rect 39200 115744 40800 115774
rect 22093 115562 22159 115565
rect 26417 115562 26483 115565
rect 22093 115560 26483 115562
rect 22093 115504 22098 115560
rect 22154 115504 26422 115560
rect 26478 115504 26483 115560
rect 22093 115502 26483 115504
rect 22093 115499 22159 115502
rect 26417 115499 26483 115502
rect -800 115426 800 115456
rect 1945 115426 2011 115429
rect -800 115424 2011 115426
rect -800 115368 1950 115424
rect 2006 115368 2011 115424
rect -800 115366 2011 115368
rect -800 115336 800 115366
rect 1945 115363 2011 115366
rect 22001 115426 22067 115429
rect 26141 115426 26207 115429
rect 22001 115424 26207 115426
rect 22001 115368 22006 115424
rect 22062 115368 26146 115424
rect 26202 115368 26207 115424
rect 22001 115366 26207 115368
rect 22001 115363 22067 115366
rect 26141 115363 26207 115366
rect 37641 115426 37707 115429
rect 39200 115426 40800 115456
rect 37641 115424 40800 115426
rect 37641 115368 37646 115424
rect 37702 115368 40800 115424
rect 37641 115366 40800 115368
rect 37641 115363 37707 115366
rect 4208 115360 4528 115361
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 115295 4528 115296
rect 34928 115360 35248 115361
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 39200 115336 40800 115366
rect 34928 115295 35248 115296
rect 20897 115290 20963 115293
rect 28809 115290 28875 115293
rect 20897 115288 28875 115290
rect 20897 115232 20902 115288
rect 20958 115232 28814 115288
rect 28870 115232 28875 115288
rect 20897 115230 28875 115232
rect 20897 115227 20963 115230
rect 28809 115227 28875 115230
rect 23289 115154 23355 115157
rect 28993 115154 29059 115157
rect 23289 115152 29059 115154
rect 23289 115096 23294 115152
rect 23350 115096 28998 115152
rect 29054 115096 29059 115152
rect 23289 115094 29059 115096
rect 23289 115091 23355 115094
rect 28993 115091 29059 115094
rect 36721 114882 36787 114885
rect 39200 114882 40800 114912
rect 36721 114880 40800 114882
rect 36721 114824 36726 114880
rect 36782 114824 40800 114880
rect 36721 114822 40800 114824
rect 36721 114819 36787 114822
rect 19568 114816 19888 114817
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 39200 114792 40800 114822
rect 19568 114751 19888 114752
rect -800 114610 800 114640
rect 2037 114610 2103 114613
rect -800 114608 2103 114610
rect -800 114552 2042 114608
rect 2098 114552 2103 114608
rect -800 114550 2103 114552
rect -800 114520 800 114550
rect 2037 114547 2103 114550
rect 20713 114610 20779 114613
rect 27705 114610 27771 114613
rect 20713 114608 27771 114610
rect 20713 114552 20718 114608
rect 20774 114552 27710 114608
rect 27766 114552 27771 114608
rect 20713 114550 27771 114552
rect 20713 114547 20779 114550
rect 27705 114547 27771 114550
rect 37089 114474 37155 114477
rect 39200 114474 40800 114504
rect 37089 114472 40800 114474
rect 37089 114416 37094 114472
rect 37150 114416 40800 114472
rect 37089 114414 40800 114416
rect 37089 114411 37155 114414
rect 39200 114384 40800 114414
rect 4208 114272 4528 114273
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 114207 4528 114208
rect 34928 114272 35248 114273
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 34928 114207 35248 114208
rect 31201 114066 31267 114069
rect 35341 114066 35407 114069
rect 31201 114064 35407 114066
rect 31201 114008 31206 114064
rect 31262 114008 35346 114064
rect 35402 114008 35407 114064
rect 31201 114006 35407 114008
rect 31201 114003 31267 114006
rect 35341 114003 35407 114006
rect 37365 114066 37431 114069
rect 39200 114066 40800 114096
rect 37365 114064 40800 114066
rect 37365 114008 37370 114064
rect 37426 114008 40800 114064
rect 37365 114006 40800 114008
rect 37365 114003 37431 114006
rect 39200 113976 40800 114006
rect -800 113794 800 113824
rect 1945 113794 2011 113797
rect -800 113792 2011 113794
rect -800 113736 1950 113792
rect 2006 113736 2011 113792
rect -800 113734 2011 113736
rect -800 113704 800 113734
rect 1945 113731 2011 113734
rect 19568 113728 19888 113729
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 19568 113663 19888 113664
rect 35801 113658 35867 113661
rect 39200 113658 40800 113688
rect 35801 113656 40800 113658
rect 35801 113600 35806 113656
rect 35862 113600 40800 113656
rect 35801 113598 40800 113600
rect 35801 113595 35867 113598
rect 39200 113568 40800 113598
rect 37365 113250 37431 113253
rect 39200 113250 40800 113280
rect 37365 113248 40800 113250
rect 37365 113192 37370 113248
rect 37426 113192 40800 113248
rect 37365 113190 40800 113192
rect 37365 113187 37431 113190
rect 4208 113184 4528 113185
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 113119 4528 113120
rect 34928 113184 35248 113185
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 39200 113160 40800 113190
rect 34928 113119 35248 113120
rect -800 112978 800 113008
rect 1853 112978 1919 112981
rect -800 112976 1919 112978
rect -800 112920 1858 112976
rect 1914 112920 1919 112976
rect -800 112918 1919 112920
rect -800 112888 800 112918
rect 1853 112915 1919 112918
rect 37365 112842 37431 112845
rect 39200 112842 40800 112872
rect 37365 112840 40800 112842
rect 37365 112784 37370 112840
rect 37426 112784 40800 112840
rect 37365 112782 40800 112784
rect 37365 112779 37431 112782
rect 39200 112752 40800 112782
rect 19568 112640 19888 112641
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 112575 19888 112576
rect 38101 112298 38167 112301
rect 39200 112298 40800 112328
rect 38101 112296 40800 112298
rect 38101 112240 38106 112296
rect 38162 112240 40800 112296
rect 38101 112238 40800 112240
rect 38101 112235 38167 112238
rect 39200 112208 40800 112238
rect -800 112162 800 112192
rect 1945 112162 2011 112165
rect -800 112160 2011 112162
rect -800 112104 1950 112160
rect 2006 112104 2011 112160
rect -800 112102 2011 112104
rect -800 112072 800 112102
rect 1945 112099 2011 112102
rect 4208 112096 4528 112097
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 112031 4528 112032
rect 34928 112096 35248 112097
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 112031 35248 112032
rect 37641 111890 37707 111893
rect 39200 111890 40800 111920
rect 37641 111888 40800 111890
rect 37641 111832 37646 111888
rect 37702 111832 40800 111888
rect 37641 111830 40800 111832
rect 37641 111827 37707 111830
rect 39200 111800 40800 111830
rect 19568 111552 19888 111553
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 19568 111487 19888 111488
rect 36537 111482 36603 111485
rect 39200 111482 40800 111512
rect 36537 111480 40800 111482
rect 36537 111424 36542 111480
rect 36598 111424 40800 111480
rect 36537 111422 40800 111424
rect 36537 111419 36603 111422
rect 39200 111392 40800 111422
rect -800 111346 800 111376
rect 1393 111346 1459 111349
rect -800 111344 1459 111346
rect -800 111288 1398 111344
rect 1454 111288 1459 111344
rect -800 111286 1459 111288
rect -800 111256 800 111286
rect 1393 111283 1459 111286
rect 37365 111074 37431 111077
rect 39200 111074 40800 111104
rect 37365 111072 40800 111074
rect 37365 111016 37370 111072
rect 37426 111016 40800 111072
rect 37365 111014 40800 111016
rect 37365 111011 37431 111014
rect 4208 111008 4528 111009
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 110943 4528 110944
rect 34928 111008 35248 111009
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 39200 110984 40800 111014
rect 34928 110943 35248 110944
rect 37457 110666 37523 110669
rect 39200 110666 40800 110696
rect 37457 110664 40800 110666
rect 37457 110608 37462 110664
rect 37518 110608 40800 110664
rect 37457 110606 40800 110608
rect 37457 110603 37523 110606
rect 39200 110576 40800 110606
rect -800 110530 800 110560
rect 1945 110530 2011 110533
rect -800 110528 2011 110530
rect -800 110472 1950 110528
rect 2006 110472 2011 110528
rect -800 110470 2011 110472
rect -800 110440 800 110470
rect 1945 110467 2011 110470
rect 19568 110464 19888 110465
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 110399 19888 110400
rect 37181 110258 37247 110261
rect 39200 110258 40800 110288
rect 37181 110256 40800 110258
rect 37181 110200 37186 110256
rect 37242 110200 40800 110256
rect 37181 110198 40800 110200
rect 37181 110195 37247 110198
rect 39200 110168 40800 110198
rect 4208 109920 4528 109921
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 109855 4528 109856
rect 34928 109920 35248 109921
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 109855 35248 109856
rect 37181 109714 37247 109717
rect 39200 109714 40800 109744
rect 37181 109712 40800 109714
rect 37181 109656 37186 109712
rect 37242 109656 40800 109712
rect 37181 109654 40800 109656
rect 37181 109651 37247 109654
rect 39200 109624 40800 109654
rect -800 109578 800 109608
rect 2037 109578 2103 109581
rect -800 109576 2103 109578
rect -800 109520 2042 109576
rect 2098 109520 2103 109576
rect -800 109518 2103 109520
rect -800 109488 800 109518
rect 2037 109515 2103 109518
rect 19568 109376 19888 109377
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 19568 109311 19888 109312
rect 37917 109306 37983 109309
rect 39200 109306 40800 109336
rect 37917 109304 40800 109306
rect 37917 109248 37922 109304
rect 37978 109248 40800 109304
rect 37917 109246 40800 109248
rect 37917 109243 37983 109246
rect 39200 109216 40800 109246
rect 37181 108898 37247 108901
rect 39200 108898 40800 108928
rect 37181 108896 40800 108898
rect 37181 108840 37186 108896
rect 37242 108840 40800 108896
rect 37181 108838 40800 108840
rect 37181 108835 37247 108838
rect 4208 108832 4528 108833
rect -800 108762 800 108792
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 108767 4528 108768
rect 34928 108832 35248 108833
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 39200 108808 40800 108838
rect 34928 108767 35248 108768
rect 1945 108762 2011 108765
rect -800 108760 2011 108762
rect -800 108704 1950 108760
rect 2006 108704 2011 108760
rect -800 108702 2011 108704
rect -800 108672 800 108702
rect 1945 108699 2011 108702
rect 37917 108490 37983 108493
rect 39200 108490 40800 108520
rect 37917 108488 40800 108490
rect 37917 108432 37922 108488
rect 37978 108432 40800 108488
rect 37917 108430 40800 108432
rect 37917 108427 37983 108430
rect 39200 108400 40800 108430
rect 19568 108288 19888 108289
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 108223 19888 108224
rect 37181 108082 37247 108085
rect 39200 108082 40800 108112
rect 37181 108080 40800 108082
rect 37181 108024 37186 108080
rect 37242 108024 40800 108080
rect 37181 108022 40800 108024
rect 37181 108019 37247 108022
rect 39200 107992 40800 108022
rect -800 107946 800 107976
rect 2037 107946 2103 107949
rect -800 107944 2103 107946
rect -800 107888 2042 107944
rect 2098 107888 2103 107944
rect -800 107886 2103 107888
rect -800 107856 800 107886
rect 2037 107883 2103 107886
rect 4208 107744 4528 107745
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 107679 4528 107680
rect 34928 107744 35248 107745
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 107679 35248 107680
rect 37181 107538 37247 107541
rect 39200 107538 40800 107568
rect 37181 107536 40800 107538
rect 37181 107480 37186 107536
rect 37242 107480 40800 107536
rect 37181 107478 40800 107480
rect 37181 107475 37247 107478
rect 39200 107448 40800 107478
rect 19568 107200 19888 107201
rect -800 107130 800 107160
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 107135 19888 107136
rect 1945 107130 2011 107133
rect -800 107128 2011 107130
rect -800 107072 1950 107128
rect 2006 107072 2011 107128
rect -800 107070 2011 107072
rect -800 107040 800 107070
rect 1945 107067 2011 107070
rect 37917 107130 37983 107133
rect 39200 107130 40800 107160
rect 37917 107128 40800 107130
rect 37917 107072 37922 107128
rect 37978 107072 40800 107128
rect 37917 107070 40800 107072
rect 37917 107067 37983 107070
rect 39200 107040 40800 107070
rect 37181 106722 37247 106725
rect 39200 106722 40800 106752
rect 37181 106720 40800 106722
rect 37181 106664 37186 106720
rect 37242 106664 40800 106720
rect 37181 106662 40800 106664
rect 37181 106659 37247 106662
rect 4208 106656 4528 106657
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 106591 4528 106592
rect 34928 106656 35248 106657
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 39200 106632 40800 106662
rect 34928 106591 35248 106592
rect -800 106314 800 106344
rect 1761 106314 1827 106317
rect -800 106312 1827 106314
rect -800 106256 1766 106312
rect 1822 106256 1827 106312
rect -800 106254 1827 106256
rect -800 106224 800 106254
rect 1761 106251 1827 106254
rect 37273 106314 37339 106317
rect 39200 106314 40800 106344
rect 37273 106312 40800 106314
rect 37273 106256 37278 106312
rect 37334 106256 40800 106312
rect 37273 106254 40800 106256
rect 37273 106251 37339 106254
rect 39200 106224 40800 106254
rect 19568 106112 19888 106113
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 19568 106047 19888 106048
rect 37181 105906 37247 105909
rect 39200 105906 40800 105936
rect 37181 105904 40800 105906
rect 37181 105848 37186 105904
rect 37242 105848 40800 105904
rect 37181 105846 40800 105848
rect 37181 105843 37247 105846
rect 39200 105816 40800 105846
rect 4208 105568 4528 105569
rect -800 105498 800 105528
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 105503 4528 105504
rect 34928 105568 35248 105569
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 105503 35248 105504
rect 1393 105498 1459 105501
rect -800 105496 1459 105498
rect -800 105440 1398 105496
rect 1454 105440 1459 105496
rect -800 105438 1459 105440
rect -800 105408 800 105438
rect 1393 105435 1459 105438
rect 37181 105498 37247 105501
rect 39200 105498 40800 105528
rect 37181 105496 40800 105498
rect 37181 105440 37186 105496
rect 37242 105440 40800 105496
rect 37181 105438 40800 105440
rect 37181 105435 37247 105438
rect 39200 105408 40800 105438
rect 19568 105024 19888 105025
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 104959 19888 104960
rect 37917 104954 37983 104957
rect 39200 104954 40800 104984
rect 37917 104952 40800 104954
rect 37917 104896 37922 104952
rect 37978 104896 40800 104952
rect 37917 104894 40800 104896
rect 37917 104891 37983 104894
rect 39200 104864 40800 104894
rect -800 104682 800 104712
rect 1853 104682 1919 104685
rect -800 104680 1919 104682
rect -800 104624 1858 104680
rect 1914 104624 1919 104680
rect -800 104622 1919 104624
rect -800 104592 800 104622
rect 1853 104619 1919 104622
rect 37181 104546 37247 104549
rect 39200 104546 40800 104576
rect 37181 104544 40800 104546
rect 37181 104488 37186 104544
rect 37242 104488 40800 104544
rect 37181 104486 40800 104488
rect 37181 104483 37247 104486
rect 4208 104480 4528 104481
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 104415 4528 104416
rect 34928 104480 35248 104481
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 39200 104456 40800 104486
rect 34928 104415 35248 104416
rect 37181 104138 37247 104141
rect 39200 104138 40800 104168
rect 37181 104136 40800 104138
rect 37181 104080 37186 104136
rect 37242 104080 40800 104136
rect 37181 104078 40800 104080
rect 37181 104075 37247 104078
rect 39200 104048 40800 104078
rect 19568 103936 19888 103937
rect -800 103866 800 103896
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 19568 103871 19888 103872
rect 1853 103866 1919 103869
rect -800 103864 1919 103866
rect -800 103808 1858 103864
rect 1914 103808 1919 103864
rect -800 103806 1919 103808
rect -800 103776 800 103806
rect 1853 103803 1919 103806
rect 37917 103730 37983 103733
rect 39200 103730 40800 103760
rect 37917 103728 40800 103730
rect 37917 103672 37922 103728
rect 37978 103672 40800 103728
rect 37917 103670 40800 103672
rect 37917 103667 37983 103670
rect 39200 103640 40800 103670
rect 4208 103392 4528 103393
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 103327 4528 103328
rect 34928 103392 35248 103393
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 103327 35248 103328
rect 37181 103322 37247 103325
rect 39200 103322 40800 103352
rect 37181 103320 40800 103322
rect 37181 103264 37186 103320
rect 37242 103264 40800 103320
rect 37181 103262 40800 103264
rect 37181 103259 37247 103262
rect 39200 103232 40800 103262
rect -800 103050 800 103080
rect 1853 103050 1919 103053
rect -800 103048 1919 103050
rect -800 102992 1858 103048
rect 1914 102992 1919 103048
rect -800 102990 1919 102992
rect -800 102960 800 102990
rect 1853 102987 1919 102990
rect 37273 102914 37339 102917
rect 39200 102914 40800 102944
rect 37273 102912 40800 102914
rect 37273 102856 37278 102912
rect 37334 102856 40800 102912
rect 37273 102854 40800 102856
rect 37273 102851 37339 102854
rect 19568 102848 19888 102849
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 39200 102824 40800 102854
rect 19568 102783 19888 102784
rect 37181 102370 37247 102373
rect 39200 102370 40800 102400
rect 37181 102368 40800 102370
rect 37181 102312 37186 102368
rect 37242 102312 40800 102368
rect 37181 102310 40800 102312
rect 37181 102307 37247 102310
rect 4208 102304 4528 102305
rect -800 102234 800 102264
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 102239 4528 102240
rect 34928 102304 35248 102305
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 39200 102280 40800 102310
rect 34928 102239 35248 102240
rect 1853 102234 1919 102237
rect -800 102232 1919 102234
rect -800 102176 1858 102232
rect 1914 102176 1919 102232
rect -800 102174 1919 102176
rect -800 102144 800 102174
rect 1853 102171 1919 102174
rect 37917 101962 37983 101965
rect 39200 101962 40800 101992
rect 37917 101960 40800 101962
rect 37917 101904 37922 101960
rect 37978 101904 40800 101960
rect 37917 101902 40800 101904
rect 37917 101899 37983 101902
rect 39200 101872 40800 101902
rect 19568 101760 19888 101761
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 19568 101695 19888 101696
rect 37181 101554 37247 101557
rect 39200 101554 40800 101584
rect 37181 101552 40800 101554
rect 37181 101496 37186 101552
rect 37242 101496 40800 101552
rect 37181 101494 40800 101496
rect 37181 101491 37247 101494
rect 39200 101464 40800 101494
rect -800 101418 800 101448
rect 1853 101418 1919 101421
rect -800 101416 1919 101418
rect -800 101360 1858 101416
rect 1914 101360 1919 101416
rect -800 101358 1919 101360
rect -800 101328 800 101358
rect 1853 101355 1919 101358
rect 4208 101216 4528 101217
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 101151 4528 101152
rect 34928 101216 35248 101217
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 34928 101151 35248 101152
rect 37917 101146 37983 101149
rect 39200 101146 40800 101176
rect 37917 101144 40800 101146
rect 37917 101088 37922 101144
rect 37978 101088 40800 101144
rect 37917 101086 40800 101088
rect 37917 101083 37983 101086
rect 39200 101056 40800 101086
rect 37181 100738 37247 100741
rect 39200 100738 40800 100768
rect 37181 100736 40800 100738
rect 37181 100680 37186 100736
rect 37242 100680 40800 100736
rect 37181 100678 40800 100680
rect 37181 100675 37247 100678
rect 19568 100672 19888 100673
rect -800 100602 800 100632
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 39200 100648 40800 100678
rect 19568 100607 19888 100608
rect 1853 100602 1919 100605
rect -800 100600 1919 100602
rect -800 100544 1858 100600
rect 1914 100544 1919 100600
rect -800 100542 1919 100544
rect -800 100512 800 100542
rect 1853 100539 1919 100542
rect 37181 100330 37247 100333
rect 39200 100330 40800 100360
rect 37181 100328 40800 100330
rect 37181 100272 37186 100328
rect 37242 100272 40800 100328
rect 37181 100270 40800 100272
rect 37181 100267 37247 100270
rect 39200 100240 40800 100270
rect 4208 100128 4528 100129
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 100063 4528 100064
rect 34928 100128 35248 100129
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 100063 35248 100064
rect 37917 99786 37983 99789
rect 39200 99786 40800 99816
rect 37917 99784 40800 99786
rect 37917 99728 37922 99784
rect 37978 99728 40800 99784
rect 37917 99726 40800 99728
rect 37917 99723 37983 99726
rect 39200 99696 40800 99726
rect -800 99650 800 99680
rect 1853 99650 1919 99653
rect -800 99648 1919 99650
rect -800 99592 1858 99648
rect 1914 99592 1919 99648
rect -800 99590 1919 99592
rect -800 99560 800 99590
rect 1853 99587 1919 99590
rect 19568 99584 19888 99585
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 99519 19888 99520
rect 37181 99378 37247 99381
rect 39200 99378 40800 99408
rect 37181 99376 40800 99378
rect 37181 99320 37186 99376
rect 37242 99320 40800 99376
rect 37181 99318 40800 99320
rect 37181 99315 37247 99318
rect 39200 99288 40800 99318
rect 4208 99040 4528 99041
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 98975 4528 98976
rect 34928 99040 35248 99041
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 34928 98975 35248 98976
rect 37181 98970 37247 98973
rect 39200 98970 40800 99000
rect 37181 98968 40800 98970
rect 37181 98912 37186 98968
rect 37242 98912 40800 98968
rect 37181 98910 40800 98912
rect 37181 98907 37247 98910
rect 39200 98880 40800 98910
rect -800 98834 800 98864
rect 1853 98834 1919 98837
rect -800 98832 1919 98834
rect -800 98776 1858 98832
rect 1914 98776 1919 98832
rect -800 98774 1919 98776
rect -800 98744 800 98774
rect 1853 98771 1919 98774
rect 37917 98562 37983 98565
rect 39200 98562 40800 98592
rect 37917 98560 40800 98562
rect 37917 98504 37922 98560
rect 37978 98504 40800 98560
rect 37917 98502 40800 98504
rect 37917 98499 37983 98502
rect 19568 98496 19888 98497
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 39200 98472 40800 98502
rect 19568 98431 19888 98432
rect 37181 98154 37247 98157
rect 39200 98154 40800 98184
rect 37181 98152 40800 98154
rect 37181 98096 37186 98152
rect 37242 98096 40800 98152
rect 37181 98094 40800 98096
rect 37181 98091 37247 98094
rect 39200 98064 40800 98094
rect -800 98018 800 98048
rect 1853 98018 1919 98021
rect -800 98016 1919 98018
rect -800 97960 1858 98016
rect 1914 97960 1919 98016
rect -800 97958 1919 97960
rect -800 97928 800 97958
rect 1853 97955 1919 97958
rect 4208 97952 4528 97953
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 97887 4528 97888
rect 34928 97952 35248 97953
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 97887 35248 97888
rect 37917 97746 37983 97749
rect 39200 97746 40800 97776
rect 37917 97744 40800 97746
rect 37917 97688 37922 97744
rect 37978 97688 40800 97744
rect 37917 97686 40800 97688
rect 37917 97683 37983 97686
rect 39200 97656 40800 97686
rect 19568 97408 19888 97409
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 97343 19888 97344
rect -800 97202 800 97232
rect 1853 97202 1919 97205
rect -800 97200 1919 97202
rect -800 97144 1858 97200
rect 1914 97144 1919 97200
rect -800 97142 1919 97144
rect -800 97112 800 97142
rect 1853 97139 1919 97142
rect 37181 97202 37247 97205
rect 39200 97202 40800 97232
rect 37181 97200 40800 97202
rect 37181 97144 37186 97200
rect 37242 97144 40800 97200
rect 37181 97142 40800 97144
rect 37181 97139 37247 97142
rect 39200 97112 40800 97142
rect 4208 96864 4528 96865
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 96799 4528 96800
rect 34928 96864 35248 96865
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 96799 35248 96800
rect 37917 96794 37983 96797
rect 39200 96794 40800 96824
rect 37917 96792 40800 96794
rect 37917 96736 37922 96792
rect 37978 96736 40800 96792
rect 37917 96734 40800 96736
rect 37917 96731 37983 96734
rect 39200 96704 40800 96734
rect -800 96386 800 96416
rect 1853 96386 1919 96389
rect -800 96384 1919 96386
rect -800 96328 1858 96384
rect 1914 96328 1919 96384
rect -800 96326 1919 96328
rect -800 96296 800 96326
rect 1853 96323 1919 96326
rect 37181 96386 37247 96389
rect 39200 96386 40800 96416
rect 37181 96384 40800 96386
rect 37181 96328 37186 96384
rect 37242 96328 40800 96384
rect 37181 96326 40800 96328
rect 37181 96323 37247 96326
rect 19568 96320 19888 96321
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 39200 96296 40800 96326
rect 19568 96255 19888 96256
rect 37181 95978 37247 95981
rect 39200 95978 40800 96008
rect 37181 95976 40800 95978
rect 37181 95920 37186 95976
rect 37242 95920 40800 95976
rect 37181 95918 40800 95920
rect 37181 95915 37247 95918
rect 39200 95888 40800 95918
rect 4208 95776 4528 95777
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 95711 4528 95712
rect 34928 95776 35248 95777
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 95711 35248 95712
rect -800 95570 800 95600
rect 1853 95570 1919 95573
rect -800 95568 1919 95570
rect -800 95512 1858 95568
rect 1914 95512 1919 95568
rect -800 95510 1919 95512
rect -800 95480 800 95510
rect 1853 95507 1919 95510
rect 37273 95570 37339 95573
rect 39200 95570 40800 95600
rect 37273 95568 40800 95570
rect 37273 95512 37278 95568
rect 37334 95512 40800 95568
rect 37273 95510 40800 95512
rect 37273 95507 37339 95510
rect 39200 95480 40800 95510
rect 19568 95232 19888 95233
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 95167 19888 95168
rect 37181 95026 37247 95029
rect 39200 95026 40800 95056
rect 37181 95024 40800 95026
rect 37181 94968 37186 95024
rect 37242 94968 40800 95024
rect 37181 94966 40800 94968
rect 37181 94963 37247 94966
rect 39200 94936 40800 94966
rect -800 94754 800 94784
rect 1853 94754 1919 94757
rect -800 94752 1919 94754
rect -800 94696 1858 94752
rect 1914 94696 1919 94752
rect -800 94694 1919 94696
rect -800 94664 800 94694
rect 1853 94691 1919 94694
rect 4208 94688 4528 94689
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 94623 4528 94624
rect 34928 94688 35248 94689
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 94623 35248 94624
rect 37917 94618 37983 94621
rect 39200 94618 40800 94648
rect 37917 94616 40800 94618
rect 37917 94560 37922 94616
rect 37978 94560 40800 94616
rect 37917 94558 40800 94560
rect 37917 94555 37983 94558
rect 39200 94528 40800 94558
rect 37273 94210 37339 94213
rect 39200 94210 40800 94240
rect 37273 94208 40800 94210
rect 37273 94152 37278 94208
rect 37334 94152 40800 94208
rect 37273 94150 40800 94152
rect 37273 94147 37339 94150
rect 19568 94144 19888 94145
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 39200 94120 40800 94150
rect 19568 94079 19888 94080
rect -800 93938 800 93968
rect 1853 93938 1919 93941
rect -800 93936 1919 93938
rect -800 93880 1858 93936
rect 1914 93880 1919 93936
rect -800 93878 1919 93880
rect -800 93848 800 93878
rect 1853 93875 1919 93878
rect 37917 93802 37983 93805
rect 39200 93802 40800 93832
rect 37917 93800 40800 93802
rect 37917 93744 37922 93800
rect 37978 93744 40800 93800
rect 37917 93742 40800 93744
rect 37917 93739 37983 93742
rect 39200 93712 40800 93742
rect 4208 93600 4528 93601
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 93535 4528 93536
rect 34928 93600 35248 93601
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 93535 35248 93536
rect 37273 93394 37339 93397
rect 39200 93394 40800 93424
rect 37273 93392 40800 93394
rect 37273 93336 37278 93392
rect 37334 93336 40800 93392
rect 37273 93334 40800 93336
rect 37273 93331 37339 93334
rect 39200 93304 40800 93334
rect -800 93122 800 93152
rect 1853 93122 1919 93125
rect -800 93120 1919 93122
rect -800 93064 1858 93120
rect 1914 93064 1919 93120
rect -800 93062 1919 93064
rect -800 93032 800 93062
rect 1853 93059 1919 93062
rect 19568 93056 19888 93057
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 92991 19888 92992
rect 37181 92986 37247 92989
rect 39200 92986 40800 93016
rect 37181 92984 40800 92986
rect 37181 92928 37186 92984
rect 37242 92928 40800 92984
rect 37181 92926 40800 92928
rect 37181 92923 37247 92926
rect 39200 92896 40800 92926
rect 4208 92512 4528 92513
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 92447 4528 92448
rect 34928 92512 35248 92513
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 92447 35248 92448
rect 38929 92442 38995 92445
rect 39200 92442 40800 92472
rect 38929 92440 40800 92442
rect 38929 92384 38934 92440
rect 38990 92384 40800 92440
rect 38929 92382 40800 92384
rect 38929 92379 38995 92382
rect 39200 92352 40800 92382
rect -800 92306 800 92336
rect 1853 92306 1919 92309
rect -800 92304 1919 92306
rect -800 92248 1858 92304
rect 1914 92248 1919 92304
rect -800 92246 1919 92248
rect -800 92216 800 92246
rect 1853 92243 1919 92246
rect 37273 92034 37339 92037
rect 39200 92034 40800 92064
rect 37273 92032 40800 92034
rect 37273 91976 37278 92032
rect 37334 91976 40800 92032
rect 37273 91974 40800 91976
rect 37273 91971 37339 91974
rect 19568 91968 19888 91969
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 39200 91944 40800 91974
rect 19568 91903 19888 91904
rect 37917 91626 37983 91629
rect 39200 91626 40800 91656
rect 37917 91624 40800 91626
rect 37917 91568 37922 91624
rect 37978 91568 40800 91624
rect 37917 91566 40800 91568
rect 37917 91563 37983 91566
rect 39200 91536 40800 91566
rect -800 91490 800 91520
rect 1853 91490 1919 91493
rect -800 91488 1919 91490
rect -800 91432 1858 91488
rect 1914 91432 1919 91488
rect -800 91430 1919 91432
rect -800 91400 800 91430
rect 1853 91427 1919 91430
rect 4208 91424 4528 91425
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 91359 4528 91360
rect 34928 91424 35248 91425
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 91359 35248 91360
rect 37273 91218 37339 91221
rect 39200 91218 40800 91248
rect 37273 91216 40800 91218
rect 37273 91160 37278 91216
rect 37334 91160 40800 91216
rect 37273 91158 40800 91160
rect 37273 91155 37339 91158
rect 39200 91128 40800 91158
rect 19568 90880 19888 90881
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 90815 19888 90816
rect 37181 90810 37247 90813
rect 39200 90810 40800 90840
rect 37181 90808 40800 90810
rect 37181 90752 37186 90808
rect 37242 90752 40800 90808
rect 37181 90750 40800 90752
rect 37181 90747 37247 90750
rect 39200 90720 40800 90750
rect -800 90674 800 90704
rect 1853 90674 1919 90677
rect -800 90672 1919 90674
rect -800 90616 1858 90672
rect 1914 90616 1919 90672
rect -800 90614 1919 90616
rect -800 90584 800 90614
rect 1853 90611 1919 90614
rect 37917 90402 37983 90405
rect 39200 90402 40800 90432
rect 37917 90400 40800 90402
rect 37917 90344 37922 90400
rect 37978 90344 40800 90400
rect 37917 90342 40800 90344
rect 37917 90339 37983 90342
rect 4208 90336 4528 90337
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 90271 4528 90272
rect 34928 90336 35248 90337
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 39200 90312 40800 90342
rect 34928 90271 35248 90272
rect 37273 89858 37339 89861
rect 39200 89858 40800 89888
rect 37273 89856 40800 89858
rect 37273 89800 37278 89856
rect 37334 89800 40800 89856
rect 37273 89798 40800 89800
rect 37273 89795 37339 89798
rect 19568 89792 19888 89793
rect -800 89722 800 89752
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 39200 89768 40800 89798
rect 19568 89727 19888 89728
rect 1853 89722 1919 89725
rect -800 89720 1919 89722
rect -800 89664 1858 89720
rect 1914 89664 1919 89720
rect -800 89662 1919 89664
rect -800 89632 800 89662
rect 1853 89659 1919 89662
rect 37917 89450 37983 89453
rect 39200 89450 40800 89480
rect 37917 89448 40800 89450
rect 37917 89392 37922 89448
rect 37978 89392 40800 89448
rect 37917 89390 40800 89392
rect 37917 89387 37983 89390
rect 39200 89360 40800 89390
rect 4208 89248 4528 89249
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 89183 4528 89184
rect 34928 89248 35248 89249
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 89183 35248 89184
rect 37273 89042 37339 89045
rect 39200 89042 40800 89072
rect 37273 89040 40800 89042
rect 37273 88984 37278 89040
rect 37334 88984 40800 89040
rect 37273 88982 40800 88984
rect 37273 88979 37339 88982
rect 39200 88952 40800 88982
rect -800 88906 800 88936
rect 1853 88906 1919 88909
rect -800 88904 1919 88906
rect -800 88848 1858 88904
rect 1914 88848 1919 88904
rect -800 88846 1919 88848
rect -800 88816 800 88846
rect 1853 88843 1919 88846
rect 19568 88704 19888 88705
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 88639 19888 88640
rect 37181 88634 37247 88637
rect 39200 88634 40800 88664
rect 37181 88632 40800 88634
rect 37181 88576 37186 88632
rect 37242 88576 40800 88632
rect 37181 88574 40800 88576
rect 37181 88571 37247 88574
rect 39200 88544 40800 88574
rect 37917 88226 37983 88229
rect 39200 88226 40800 88256
rect 37917 88224 40800 88226
rect 37917 88168 37922 88224
rect 37978 88168 40800 88224
rect 37917 88166 40800 88168
rect 37917 88163 37983 88166
rect 4208 88160 4528 88161
rect -800 88090 800 88120
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 88095 4528 88096
rect 34928 88160 35248 88161
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 39200 88136 40800 88166
rect 34928 88095 35248 88096
rect 1853 88090 1919 88093
rect -800 88088 1919 88090
rect -800 88032 1858 88088
rect 1914 88032 1919 88088
rect -800 88030 1919 88032
rect -800 88000 800 88030
rect 1853 88027 1919 88030
rect 28165 87954 28231 87957
rect 28809 87954 28875 87957
rect 28165 87952 28875 87954
rect 28165 87896 28170 87952
rect 28226 87896 28814 87952
rect 28870 87896 28875 87952
rect 28165 87894 28875 87896
rect 28165 87891 28231 87894
rect 28809 87891 28875 87894
rect 27521 87818 27587 87821
rect 28165 87818 28231 87821
rect 27521 87816 28231 87818
rect 27521 87760 27526 87816
rect 27582 87760 28170 87816
rect 28226 87760 28231 87816
rect 27521 87758 28231 87760
rect 27521 87755 27587 87758
rect 28165 87755 28231 87758
rect 37273 87818 37339 87821
rect 39200 87818 40800 87848
rect 37273 87816 40800 87818
rect 37273 87760 37278 87816
rect 37334 87760 40800 87816
rect 37273 87758 40800 87760
rect 37273 87755 37339 87758
rect 39200 87728 40800 87758
rect 19568 87616 19888 87617
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 87551 19888 87552
rect 35617 87546 35683 87549
rect 35574 87544 35683 87546
rect 35574 87488 35622 87544
rect 35678 87488 35683 87544
rect 35574 87483 35683 87488
rect -800 87274 800 87304
rect 1853 87274 1919 87277
rect 34697 87274 34763 87277
rect -800 87272 1919 87274
rect -800 87216 1858 87272
rect 1914 87216 1919 87272
rect -800 87214 1919 87216
rect -800 87184 800 87214
rect 1853 87211 1919 87214
rect 34654 87272 34763 87274
rect 34654 87216 34702 87272
rect 34758 87216 34763 87272
rect 34654 87211 34763 87216
rect 35341 87274 35407 87277
rect 35341 87272 35450 87274
rect 35341 87216 35346 87272
rect 35402 87216 35450 87272
rect 35341 87211 35450 87216
rect 4208 87072 4528 87073
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 87007 4528 87008
rect 34654 87005 34714 87211
rect 34928 87072 35248 87073
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 87007 35248 87008
rect 35390 87005 35450 87211
rect 35574 87005 35634 87483
rect 37917 87274 37983 87277
rect 39200 87274 40800 87304
rect 37917 87272 40800 87274
rect 37917 87216 37922 87272
rect 37978 87216 40800 87272
rect 37917 87214 40800 87216
rect 37917 87211 37983 87214
rect 39200 87184 40800 87214
rect 32489 87002 32555 87005
rect 33961 87002 34027 87005
rect 32489 87000 34027 87002
rect 32489 86944 32494 87000
rect 32550 86944 33966 87000
rect 34022 86944 34027 87000
rect 32489 86942 34027 86944
rect 34654 87000 34763 87005
rect 34654 86944 34702 87000
rect 34758 86944 34763 87000
rect 34654 86942 34763 86944
rect 35390 87000 35499 87005
rect 35390 86944 35438 87000
rect 35494 86944 35499 87000
rect 35390 86942 35499 86944
rect 35574 87000 35683 87005
rect 35574 86944 35622 87000
rect 35678 86944 35683 87000
rect 35574 86942 35683 86944
rect 32489 86939 32555 86942
rect 33961 86939 34027 86942
rect 34697 86939 34763 86942
rect 35433 86939 35499 86942
rect 35617 86939 35683 86942
rect 37273 86866 37339 86869
rect 39200 86866 40800 86896
rect 37273 86864 40800 86866
rect 37273 86808 37278 86864
rect 37334 86808 40800 86864
rect 37273 86806 40800 86808
rect 37273 86803 37339 86806
rect 39200 86776 40800 86806
rect 27613 86730 27679 86733
rect 28901 86730 28967 86733
rect 27613 86728 28967 86730
rect 27613 86672 27618 86728
rect 27674 86672 28906 86728
rect 28962 86672 28967 86728
rect 27613 86670 28967 86672
rect 27613 86667 27679 86670
rect 28901 86667 28967 86670
rect 32765 86730 32831 86733
rect 38745 86730 38811 86733
rect 32765 86728 38811 86730
rect 32765 86672 32770 86728
rect 32826 86672 38750 86728
rect 38806 86672 38811 86728
rect 32765 86670 38811 86672
rect 32765 86667 32831 86670
rect 38745 86667 38811 86670
rect 38009 86594 38075 86597
rect 32814 86592 38075 86594
rect 32814 86536 38014 86592
rect 38070 86536 38075 86592
rect 32814 86534 38075 86536
rect 19568 86528 19888 86529
rect -800 86458 800 86488
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 86463 19888 86464
rect 1853 86458 1919 86461
rect -800 86456 1919 86458
rect -800 86400 1858 86456
rect 1914 86400 1919 86456
rect -800 86398 1919 86400
rect -800 86368 800 86398
rect 1853 86395 1919 86398
rect 27613 86322 27679 86325
rect 28257 86322 28323 86325
rect 27613 86320 28323 86322
rect 27613 86264 27618 86320
rect 27674 86264 28262 86320
rect 28318 86264 28323 86320
rect 27613 86262 28323 86264
rect 27613 86259 27679 86262
rect 28257 86259 28323 86262
rect 29269 86322 29335 86325
rect 32814 86322 32874 86534
rect 38009 86531 38075 86534
rect 37181 86458 37247 86461
rect 39200 86458 40800 86488
rect 37181 86456 40800 86458
rect 37181 86400 37186 86456
rect 37242 86400 40800 86456
rect 37181 86398 40800 86400
rect 37181 86395 37247 86398
rect 39200 86368 40800 86398
rect 29269 86320 32874 86322
rect 29269 86264 29274 86320
rect 29330 86264 32874 86320
rect 29269 86262 32874 86264
rect 29269 86259 29335 86262
rect 27153 86186 27219 86189
rect 28901 86186 28967 86189
rect 29269 86186 29335 86189
rect 27153 86184 29335 86186
rect 27153 86128 27158 86184
rect 27214 86128 28906 86184
rect 28962 86128 29274 86184
rect 29330 86128 29335 86184
rect 27153 86126 29335 86128
rect 27153 86123 27219 86126
rect 28901 86123 28967 86126
rect 29269 86123 29335 86126
rect 37917 86050 37983 86053
rect 39200 86050 40800 86080
rect 37917 86048 40800 86050
rect 37917 85992 37922 86048
rect 37978 85992 40800 86048
rect 37917 85990 40800 85992
rect 37917 85987 37983 85990
rect 4208 85984 4528 85985
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 85919 4528 85920
rect 34928 85984 35248 85985
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 39200 85960 40800 85990
rect 34928 85919 35248 85920
rect -800 85642 800 85672
rect 1853 85642 1919 85645
rect -800 85640 1919 85642
rect -800 85584 1858 85640
rect 1914 85584 1919 85640
rect -800 85582 1919 85584
rect -800 85552 800 85582
rect 1853 85579 1919 85582
rect 37273 85642 37339 85645
rect 39200 85642 40800 85672
rect 37273 85640 40800 85642
rect 37273 85584 37278 85640
rect 37334 85584 40800 85640
rect 37273 85582 40800 85584
rect 37273 85579 37339 85582
rect 39200 85552 40800 85582
rect 28809 85506 28875 85509
rect 29269 85506 29335 85509
rect 28809 85504 29335 85506
rect 28809 85448 28814 85504
rect 28870 85448 29274 85504
rect 29330 85448 29335 85504
rect 28809 85446 29335 85448
rect 28809 85443 28875 85446
rect 29269 85443 29335 85446
rect 19568 85440 19888 85441
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 85375 19888 85376
rect 37917 85234 37983 85237
rect 39200 85234 40800 85264
rect 37917 85232 40800 85234
rect 37917 85176 37922 85232
rect 37978 85176 40800 85232
rect 37917 85174 40800 85176
rect 37917 85171 37983 85174
rect 39200 85144 40800 85174
rect 4208 84896 4528 84897
rect -800 84826 800 84856
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 84831 4528 84832
rect 34928 84896 35248 84897
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 84831 35248 84832
rect 1853 84826 1919 84829
rect -800 84824 1919 84826
rect -800 84768 1858 84824
rect 1914 84768 1919 84824
rect -800 84766 1919 84768
rect -800 84736 800 84766
rect 1853 84763 1919 84766
rect 27521 84690 27587 84693
rect 29361 84690 29427 84693
rect 27521 84688 29427 84690
rect 27521 84632 27526 84688
rect 27582 84632 29366 84688
rect 29422 84632 29427 84688
rect 27521 84630 29427 84632
rect 27521 84627 27587 84630
rect 29361 84627 29427 84630
rect 37273 84690 37339 84693
rect 39200 84690 40800 84720
rect 37273 84688 40800 84690
rect 37273 84632 37278 84688
rect 37334 84632 40800 84688
rect 37273 84630 40800 84632
rect 37273 84627 37339 84630
rect 39200 84600 40800 84630
rect 28993 84554 29059 84557
rect 30373 84554 30439 84557
rect 28993 84552 30439 84554
rect 28993 84496 28998 84552
rect 29054 84496 30378 84552
rect 30434 84496 30439 84552
rect 28993 84494 30439 84496
rect 28993 84491 29059 84494
rect 30373 84491 30439 84494
rect 19568 84352 19888 84353
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 84287 19888 84288
rect 25957 84282 26023 84285
rect 28441 84282 28507 84285
rect 25957 84280 28507 84282
rect 25957 84224 25962 84280
rect 26018 84224 28446 84280
rect 28502 84224 28507 84280
rect 25957 84222 28507 84224
rect 25957 84219 26023 84222
rect 28441 84219 28507 84222
rect 29361 84282 29427 84285
rect 37181 84282 37247 84285
rect 39200 84282 40800 84312
rect 29361 84280 29562 84282
rect 29361 84224 29366 84280
rect 29422 84224 29562 84280
rect 29361 84222 29562 84224
rect 29361 84219 29427 84222
rect -800 84010 800 84040
rect 1853 84010 1919 84013
rect -800 84008 1919 84010
rect -800 83952 1858 84008
rect 1914 83952 1919 84008
rect -800 83950 1919 83952
rect -800 83920 800 83950
rect 1853 83947 1919 83950
rect 28257 84010 28323 84013
rect 29085 84010 29151 84013
rect 28257 84008 29151 84010
rect 28257 83952 28262 84008
rect 28318 83952 29090 84008
rect 29146 83952 29151 84008
rect 28257 83950 29151 83952
rect 28257 83947 28323 83950
rect 29085 83947 29151 83950
rect 4208 83808 4528 83809
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 83743 4528 83744
rect 29502 83602 29562 84222
rect 37181 84280 40800 84282
rect 37181 84224 37186 84280
rect 37242 84224 40800 84280
rect 37181 84222 40800 84224
rect 37181 84219 37247 84222
rect 39200 84192 40800 84222
rect 31477 84008 31543 84013
rect 31477 83952 31482 84008
rect 31538 83952 31543 84008
rect 31477 83947 31543 83952
rect 31201 83874 31267 83877
rect 31480 83874 31540 83947
rect 30376 83872 31540 83874
rect 30376 83816 31206 83872
rect 31262 83816 31540 83872
rect 30376 83814 31540 83816
rect 37917 83874 37983 83877
rect 39200 83874 40800 83904
rect 37917 83872 40800 83874
rect 37917 83816 37922 83872
rect 37978 83816 40800 83872
rect 37917 83814 40800 83816
rect 30376 83741 30436 83814
rect 31201 83811 31267 83814
rect 37917 83811 37983 83814
rect 34928 83808 35248 83809
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 39200 83784 40800 83814
rect 34928 83743 35248 83744
rect 29637 83738 29703 83741
rect 29637 83736 29930 83738
rect 29637 83680 29642 83736
rect 29698 83680 29930 83736
rect 29637 83678 29930 83680
rect 29637 83675 29703 83678
rect 29637 83602 29703 83605
rect 29502 83600 29703 83602
rect 29502 83544 29642 83600
rect 29698 83544 29703 83600
rect 29502 83542 29703 83544
rect 29637 83539 29703 83542
rect 28257 83466 28323 83469
rect 28625 83466 28691 83469
rect 29870 83466 29930 83678
rect 30373 83736 30439 83741
rect 30373 83680 30378 83736
rect 30434 83680 30439 83736
rect 30373 83675 30439 83680
rect 28257 83464 28504 83466
rect 28257 83408 28262 83464
rect 28318 83408 28504 83464
rect 28257 83406 28504 83408
rect 28257 83403 28323 83406
rect 19568 83264 19888 83265
rect -800 83194 800 83224
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 83199 19888 83200
rect 1393 83194 1459 83197
rect -800 83192 1459 83194
rect -800 83136 1398 83192
rect 1454 83136 1459 83192
rect -800 83134 1459 83136
rect 28444 83194 28504 83406
rect 28625 83464 29930 83466
rect 28625 83408 28630 83464
rect 28686 83408 29930 83464
rect 28625 83406 29930 83408
rect 37273 83466 37339 83469
rect 39200 83466 40800 83496
rect 37273 83464 40800 83466
rect 37273 83408 37278 83464
rect 37334 83408 40800 83464
rect 37273 83406 40800 83408
rect 28625 83403 28691 83406
rect 37273 83403 37339 83406
rect 39200 83376 40800 83406
rect 28625 83194 28691 83197
rect 28444 83192 28691 83194
rect 28444 83136 28630 83192
rect 28686 83136 28691 83192
rect 28444 83134 28691 83136
rect -800 83104 800 83134
rect 1393 83131 1459 83134
rect 28625 83131 28691 83134
rect 37917 83058 37983 83061
rect 39200 83058 40800 83088
rect 37917 83056 40800 83058
rect 37917 83000 37922 83056
rect 37978 83000 40800 83056
rect 37917 82998 40800 83000
rect 37917 82995 37983 82998
rect 39200 82968 40800 82998
rect 4208 82720 4528 82721
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 82655 4528 82656
rect 34928 82720 35248 82721
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 82655 35248 82656
rect 37273 82514 37339 82517
rect 39200 82514 40800 82544
rect 37273 82512 40800 82514
rect 37273 82456 37278 82512
rect 37334 82456 40800 82512
rect 37273 82454 40800 82456
rect 37273 82451 37339 82454
rect 39200 82424 40800 82454
rect -800 82378 800 82408
rect 1853 82378 1919 82381
rect -800 82376 1919 82378
rect -800 82320 1858 82376
rect 1914 82320 1919 82376
rect -800 82318 1919 82320
rect -800 82288 800 82318
rect 1853 82315 1919 82318
rect 28165 82242 28231 82245
rect 28717 82242 28783 82245
rect 28165 82240 28783 82242
rect 28165 82184 28170 82240
rect 28226 82184 28722 82240
rect 28778 82184 28783 82240
rect 28165 82182 28783 82184
rect 28165 82179 28231 82182
rect 28717 82179 28783 82182
rect 19568 82176 19888 82177
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 82111 19888 82112
rect 37181 82106 37247 82109
rect 39200 82106 40800 82136
rect 37181 82104 40800 82106
rect 37181 82048 37186 82104
rect 37242 82048 40800 82104
rect 37181 82046 40800 82048
rect 37181 82043 37247 82046
rect 39200 82016 40800 82046
rect 25497 81698 25563 81701
rect 33961 81698 34027 81701
rect 25497 81696 34027 81698
rect 25497 81640 25502 81696
rect 25558 81640 33966 81696
rect 34022 81640 34027 81696
rect 25497 81638 34027 81640
rect 25497 81635 25563 81638
rect 33961 81635 34027 81638
rect 37917 81698 37983 81701
rect 39200 81698 40800 81728
rect 37917 81696 40800 81698
rect 37917 81640 37922 81696
rect 37978 81640 40800 81696
rect 37917 81638 40800 81640
rect 37917 81635 37983 81638
rect 4208 81632 4528 81633
rect -800 81562 800 81592
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 81567 4528 81568
rect 34928 81632 35248 81633
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 39200 81608 40800 81638
rect 34928 81567 35248 81568
rect 1853 81562 1919 81565
rect -800 81560 1919 81562
rect -800 81504 1858 81560
rect 1914 81504 1919 81560
rect -800 81502 1919 81504
rect -800 81472 800 81502
rect 1853 81499 1919 81502
rect 29177 81562 29243 81565
rect 31109 81562 31175 81565
rect 29177 81560 31175 81562
rect 29177 81504 29182 81560
rect 29238 81504 31114 81560
rect 31170 81504 31175 81560
rect 29177 81502 31175 81504
rect 29177 81499 29243 81502
rect 31109 81499 31175 81502
rect 27429 81424 27495 81429
rect 27429 81368 27434 81424
rect 27490 81368 27495 81424
rect 27429 81363 27495 81368
rect 29637 81426 29703 81429
rect 29637 81424 30298 81426
rect 29637 81368 29642 81424
rect 29698 81368 30298 81424
rect 29637 81366 30298 81368
rect 29637 81363 29703 81366
rect 27432 81154 27492 81363
rect 27432 81094 27538 81154
rect 19568 81088 19888 81089
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 81023 19888 81024
rect 27337 80882 27403 80885
rect 27478 80882 27538 81094
rect 27337 80880 27538 80882
rect 27337 80824 27342 80880
rect 27398 80824 27538 80880
rect 27337 80822 27538 80824
rect 27337 80819 27403 80822
rect -800 80746 800 80776
rect 1393 80746 1459 80749
rect -800 80744 1459 80746
rect -800 80688 1398 80744
rect 1454 80688 1459 80744
rect -800 80686 1459 80688
rect -800 80656 800 80686
rect 1393 80683 1459 80686
rect 4208 80544 4528 80545
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 80479 4528 80480
rect 30097 80474 30163 80477
rect 29134 80472 30163 80474
rect 29134 80416 30102 80472
rect 30158 80416 30163 80472
rect 29134 80414 30163 80416
rect 28165 80066 28231 80069
rect 28625 80066 28691 80069
rect 28165 80064 28691 80066
rect 28165 80008 28170 80064
rect 28226 80008 28630 80064
rect 28686 80008 28691 80064
rect 28165 80006 28691 80008
rect 28165 80003 28231 80006
rect 28625 80003 28691 80006
rect 19568 80000 19888 80001
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 79935 19888 79936
rect 26049 79930 26115 79933
rect 28441 79930 28507 79933
rect 26049 79928 28507 79930
rect 26049 79872 26054 79928
rect 26110 79872 28446 79928
rect 28502 79872 28507 79928
rect 26049 79870 28507 79872
rect 26049 79867 26115 79870
rect 28441 79867 28507 79870
rect -800 79794 800 79824
rect 1393 79794 1459 79797
rect 27429 79794 27495 79797
rect -800 79792 1459 79794
rect -800 79736 1398 79792
rect 1454 79736 1459 79792
rect -800 79734 1459 79736
rect -800 79704 800 79734
rect 1393 79731 1459 79734
rect 26558 79792 27495 79794
rect 26558 79736 27434 79792
rect 27490 79736 27495 79792
rect 26558 79734 27495 79736
rect 26558 79661 26618 79734
rect 27429 79731 27495 79734
rect 26509 79656 26618 79661
rect 26509 79600 26514 79656
rect 26570 79600 26618 79656
rect 26509 79598 26618 79600
rect 27429 79658 27495 79661
rect 28165 79658 28231 79661
rect 27429 79656 28231 79658
rect 27429 79600 27434 79656
rect 27490 79600 28170 79656
rect 28226 79600 28231 79656
rect 27429 79598 28231 79600
rect 26509 79595 26575 79598
rect 27429 79595 27495 79598
rect 28165 79595 28231 79598
rect 28993 79658 29059 79661
rect 29134 79658 29194 80414
rect 30097 80411 30163 80414
rect 29269 80338 29335 80341
rect 29269 80336 29378 80338
rect 29269 80280 29274 80336
rect 29330 80280 29378 80336
rect 29269 80275 29378 80280
rect 29318 80066 29378 80275
rect 28993 79656 29194 79658
rect 28993 79600 28998 79656
rect 29054 79600 29194 79656
rect 28993 79598 29194 79600
rect 28993 79595 29059 79598
rect 25497 79522 25563 79525
rect 28625 79522 28691 79525
rect 25497 79520 28691 79522
rect 25497 79464 25502 79520
rect 25558 79464 28630 79520
rect 28686 79464 28691 79520
rect 25497 79462 28691 79464
rect 25497 79459 25563 79462
rect 28625 79459 28691 79462
rect 4208 79456 4528 79457
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 79391 4528 79392
rect 29134 79386 29194 79598
rect 27570 79326 29194 79386
rect 29272 80006 29378 80066
rect 30238 80073 30298 81366
rect 37273 81290 37339 81293
rect 39200 81290 40800 81320
rect 37273 81288 40800 81290
rect 37273 81232 37278 81288
rect 37334 81232 40800 81288
rect 37273 81230 40800 81232
rect 37273 81227 37339 81230
rect 39200 81200 40800 81230
rect 31201 81018 31267 81021
rect 33685 81018 33751 81021
rect 31201 81016 33751 81018
rect 31201 80960 31206 81016
rect 31262 80960 33690 81016
rect 33746 80960 33751 81016
rect 31201 80958 33751 80960
rect 31201 80955 31267 80958
rect 33685 80955 33751 80958
rect 37917 80882 37983 80885
rect 39200 80882 40800 80912
rect 37917 80880 40800 80882
rect 37917 80824 37922 80880
rect 37978 80824 40800 80880
rect 37917 80822 40800 80824
rect 37917 80819 37983 80822
rect 39200 80792 40800 80822
rect 34928 80544 35248 80545
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 80479 35248 80480
rect 30649 80474 30715 80477
rect 31385 80474 31451 80477
rect 30649 80472 31451 80474
rect 30649 80416 30654 80472
rect 30710 80416 31390 80472
rect 31446 80416 31451 80472
rect 30649 80414 31451 80416
rect 30649 80411 30715 80414
rect 31385 80411 31451 80414
rect 37273 80474 37339 80477
rect 39200 80474 40800 80504
rect 37273 80472 40800 80474
rect 37273 80416 37278 80472
rect 37334 80416 40800 80472
rect 37273 80414 40800 80416
rect 37273 80411 37339 80414
rect 39200 80384 40800 80414
rect 31385 80338 31451 80341
rect 38837 80338 38903 80341
rect 31385 80336 38903 80338
rect 31385 80280 31390 80336
rect 31446 80280 38842 80336
rect 38898 80280 38903 80336
rect 31385 80278 38903 80280
rect 31385 80275 31451 80278
rect 38837 80275 38903 80278
rect 30238 80068 30347 80073
rect 30238 80012 30286 80068
rect 30342 80012 30347 80068
rect 30238 80010 30347 80012
rect 30281 80007 30347 80010
rect -800 78978 800 79008
rect 1853 78978 1919 78981
rect -800 78976 1919 78978
rect -800 78920 1858 78976
rect 1914 78920 1919 78976
rect -800 78918 1919 78920
rect -800 78888 800 78918
rect 1853 78915 1919 78918
rect 19568 78912 19888 78913
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 78847 19888 78848
rect 26417 78570 26483 78573
rect 27570 78570 27630 79326
rect 28165 79250 28231 79253
rect 28030 79248 28231 79250
rect 28030 79192 28170 79248
rect 28226 79192 28231 79248
rect 28030 79190 28231 79192
rect 28030 78842 28090 79190
rect 28165 79187 28231 79190
rect 28349 79250 28415 79253
rect 28625 79250 28691 79253
rect 28349 79248 28691 79250
rect 28349 79192 28354 79248
rect 28410 79192 28630 79248
rect 28686 79192 28691 79248
rect 28349 79190 28691 79192
rect 28349 79187 28415 79190
rect 28625 79187 28691 79190
rect 28165 79114 28231 79117
rect 29085 79114 29151 79117
rect 28165 79112 29151 79114
rect 28165 79056 28170 79112
rect 28226 79056 29090 79112
rect 29146 79056 29151 79112
rect 28165 79054 29151 79056
rect 28165 79051 28231 79054
rect 29085 79051 29151 79054
rect 28993 78978 29059 78981
rect 29272 78978 29332 80006
rect 37181 79930 37247 79933
rect 39200 79930 40800 79960
rect 37181 79928 40800 79930
rect 37181 79872 37186 79928
rect 37242 79872 40800 79928
rect 37181 79870 40800 79872
rect 37181 79867 37247 79870
rect 39200 79840 40800 79870
rect 30373 79658 30439 79661
rect 30373 79656 30482 79658
rect 30373 79600 30378 79656
rect 30434 79600 30482 79656
rect 30373 79595 30482 79600
rect 30422 78981 30482 79595
rect 37917 79522 37983 79525
rect 39200 79522 40800 79552
rect 37917 79520 40800 79522
rect 37917 79464 37922 79520
rect 37978 79464 40800 79520
rect 37917 79462 40800 79464
rect 37917 79459 37983 79462
rect 34928 79456 35248 79457
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 39200 79432 40800 79462
rect 34928 79391 35248 79392
rect 37917 79114 37983 79117
rect 39200 79114 40800 79144
rect 37917 79112 40800 79114
rect 37917 79056 37922 79112
rect 37978 79056 40800 79112
rect 37917 79054 40800 79056
rect 37917 79051 37983 79054
rect 39200 79024 40800 79054
rect 28993 78976 29332 78978
rect 28993 78920 28998 78976
rect 29054 78920 29332 78976
rect 28993 78918 29332 78920
rect 30373 78976 30482 78981
rect 30373 78920 30378 78976
rect 30434 78920 30482 78976
rect 30373 78918 30482 78920
rect 28993 78915 29059 78918
rect 30373 78915 30439 78918
rect 32397 78842 32463 78845
rect 28030 78840 32463 78842
rect 28030 78784 32402 78840
rect 32458 78784 32463 78840
rect 28030 78782 32463 78784
rect 32397 78779 32463 78782
rect 37181 78706 37247 78709
rect 39200 78706 40800 78736
rect 37181 78704 40800 78706
rect 37181 78648 37186 78704
rect 37242 78648 40800 78704
rect 37181 78646 40800 78648
rect 37181 78643 37247 78646
rect 39200 78616 40800 78646
rect 26417 78568 27630 78570
rect 26417 78512 26422 78568
rect 26478 78512 27630 78568
rect 26417 78510 27630 78512
rect 26417 78507 26483 78510
rect 4208 78368 4528 78369
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 78303 4528 78304
rect 34928 78368 35248 78369
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 78303 35248 78304
rect 37181 78298 37247 78301
rect 39200 78298 40800 78328
rect 37181 78296 40800 78298
rect 37181 78240 37186 78296
rect 37242 78240 40800 78296
rect 37181 78238 40800 78240
rect 37181 78235 37247 78238
rect 39200 78208 40800 78238
rect -800 78162 800 78192
rect 1853 78162 1919 78165
rect -800 78160 1919 78162
rect -800 78104 1858 78160
rect 1914 78104 1919 78160
rect -800 78102 1919 78104
rect -800 78072 800 78102
rect 1853 78099 1919 78102
rect 37917 77890 37983 77893
rect 39200 77890 40800 77920
rect 37917 77888 40800 77890
rect 37917 77832 37922 77888
rect 37978 77832 40800 77888
rect 37917 77830 40800 77832
rect 37917 77827 37983 77830
rect 19568 77824 19888 77825
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 39200 77800 40800 77830
rect 19568 77759 19888 77760
rect -800 77346 800 77376
rect 1393 77346 1459 77349
rect -800 77344 1459 77346
rect -800 77288 1398 77344
rect 1454 77288 1459 77344
rect -800 77286 1459 77288
rect -800 77256 800 77286
rect 1393 77283 1459 77286
rect 37181 77346 37247 77349
rect 39200 77346 40800 77376
rect 37181 77344 40800 77346
rect 37181 77288 37186 77344
rect 37242 77288 40800 77344
rect 37181 77286 40800 77288
rect 37181 77283 37247 77286
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 34928 77280 35248 77281
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 39200 77256 40800 77286
rect 34928 77215 35248 77216
rect 37917 76938 37983 76941
rect 39200 76938 40800 76968
rect 37917 76936 40800 76938
rect 37917 76880 37922 76936
rect 37978 76880 40800 76936
rect 37917 76878 40800 76880
rect 37917 76875 37983 76878
rect 39200 76848 40800 76878
rect 19568 76736 19888 76737
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 76671 19888 76672
rect -800 76530 800 76560
rect 1393 76530 1459 76533
rect -800 76528 1459 76530
rect -800 76472 1398 76528
rect 1454 76472 1459 76528
rect -800 76470 1459 76472
rect -800 76440 800 76470
rect 1393 76467 1459 76470
rect 37181 76530 37247 76533
rect 39200 76530 40800 76560
rect 37181 76528 40800 76530
rect 37181 76472 37186 76528
rect 37242 76472 40800 76528
rect 37181 76470 40800 76472
rect 37181 76467 37247 76470
rect 39200 76440 40800 76470
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 34928 76192 35248 76193
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 76127 35248 76128
rect 37181 76122 37247 76125
rect 39200 76122 40800 76152
rect 37181 76120 40800 76122
rect 37181 76064 37186 76120
rect 37242 76064 40800 76120
rect 37181 76062 40800 76064
rect 37181 76059 37247 76062
rect 39200 76032 40800 76062
rect -800 75714 800 75744
rect 1853 75714 1919 75717
rect -800 75712 1919 75714
rect -800 75656 1858 75712
rect 1914 75656 1919 75712
rect -800 75654 1919 75656
rect -800 75624 800 75654
rect 1853 75651 1919 75654
rect 37917 75714 37983 75717
rect 39200 75714 40800 75744
rect 37917 75712 40800 75714
rect 37917 75656 37922 75712
rect 37978 75656 40800 75712
rect 37917 75654 40800 75656
rect 37917 75651 37983 75654
rect 19568 75648 19888 75649
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 39200 75624 40800 75654
rect 19568 75583 19888 75584
rect 37181 75306 37247 75309
rect 39200 75306 40800 75336
rect 37181 75304 40800 75306
rect 37181 75248 37186 75304
rect 37242 75248 40800 75304
rect 37181 75246 40800 75248
rect 37181 75243 37247 75246
rect 39200 75216 40800 75246
rect 4208 75104 4528 75105
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 34928 75104 35248 75105
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 75039 35248 75040
rect -800 74898 800 74928
rect 1853 74898 1919 74901
rect -800 74896 1919 74898
rect -800 74840 1858 74896
rect 1914 74840 1919 74896
rect -800 74838 1919 74840
rect -800 74808 800 74838
rect 1853 74835 1919 74838
rect 37917 74762 37983 74765
rect 39200 74762 40800 74792
rect 37917 74760 40800 74762
rect 37917 74704 37922 74760
rect 37978 74704 40800 74760
rect 37917 74702 40800 74704
rect 37917 74699 37983 74702
rect 39200 74672 40800 74702
rect 19568 74560 19888 74561
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 74495 19888 74496
rect 37181 74354 37247 74357
rect 39200 74354 40800 74384
rect 37181 74352 40800 74354
rect 37181 74296 37186 74352
rect 37242 74296 40800 74352
rect 37181 74294 40800 74296
rect 37181 74291 37247 74294
rect 39200 74264 40800 74294
rect -800 74082 800 74112
rect 1853 74082 1919 74085
rect -800 74080 1919 74082
rect -800 74024 1858 74080
rect 1914 74024 1919 74080
rect -800 74022 1919 74024
rect -800 73992 800 74022
rect 1853 74019 1919 74022
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 34928 74016 35248 74017
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 73951 35248 73952
rect 37181 73946 37247 73949
rect 39200 73946 40800 73976
rect 37181 73944 40800 73946
rect 37181 73888 37186 73944
rect 37242 73888 40800 73944
rect 37181 73886 40800 73888
rect 37181 73883 37247 73886
rect 39200 73856 40800 73886
rect 37917 73538 37983 73541
rect 39200 73538 40800 73568
rect 37917 73536 40800 73538
rect 37917 73480 37922 73536
rect 37978 73480 40800 73536
rect 37917 73478 40800 73480
rect 37917 73475 37983 73478
rect 19568 73472 19888 73473
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 39200 73448 40800 73478
rect 19568 73407 19888 73408
rect -800 73266 800 73296
rect 1853 73266 1919 73269
rect -800 73264 1919 73266
rect -800 73208 1858 73264
rect 1914 73208 1919 73264
rect -800 73206 1919 73208
rect -800 73176 800 73206
rect 1853 73203 1919 73206
rect 37181 73130 37247 73133
rect 39200 73130 40800 73160
rect 37181 73128 40800 73130
rect 37181 73072 37186 73128
rect 37242 73072 40800 73128
rect 37181 73070 40800 73072
rect 37181 73067 37247 73070
rect 39200 73040 40800 73070
rect 4208 72928 4528 72929
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 34928 72928 35248 72929
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 72863 35248 72864
rect 37917 72722 37983 72725
rect 39200 72722 40800 72752
rect 37917 72720 40800 72722
rect 37917 72664 37922 72720
rect 37978 72664 40800 72720
rect 37917 72662 40800 72664
rect 37917 72659 37983 72662
rect 39200 72632 40800 72662
rect -800 72450 800 72480
rect 1853 72450 1919 72453
rect -800 72448 1919 72450
rect -800 72392 1858 72448
rect 1914 72392 1919 72448
rect -800 72390 1919 72392
rect -800 72360 800 72390
rect 1853 72387 1919 72390
rect 19568 72384 19888 72385
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 72319 19888 72320
rect 37181 72178 37247 72181
rect 39200 72178 40800 72208
rect 37181 72176 40800 72178
rect 37181 72120 37186 72176
rect 37242 72120 40800 72176
rect 37181 72118 40800 72120
rect 37181 72115 37247 72118
rect 39200 72088 40800 72118
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 34928 71840 35248 71841
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 71775 35248 71776
rect 37181 71770 37247 71773
rect 39200 71770 40800 71800
rect 37181 71768 40800 71770
rect 37181 71712 37186 71768
rect 37242 71712 40800 71768
rect 37181 71710 40800 71712
rect 37181 71707 37247 71710
rect 39200 71680 40800 71710
rect -800 71634 800 71664
rect 1853 71634 1919 71637
rect -800 71632 1919 71634
rect -800 71576 1858 71632
rect 1914 71576 1919 71632
rect -800 71574 1919 71576
rect -800 71544 800 71574
rect 1853 71571 1919 71574
rect 37917 71362 37983 71365
rect 39200 71362 40800 71392
rect 37917 71360 40800 71362
rect 37917 71304 37922 71360
rect 37978 71304 40800 71360
rect 37917 71302 40800 71304
rect 37917 71299 37983 71302
rect 19568 71296 19888 71297
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 39200 71272 40800 71302
rect 19568 71231 19888 71232
rect 37181 70954 37247 70957
rect 39200 70954 40800 70984
rect 37181 70952 40800 70954
rect 37181 70896 37186 70952
rect 37242 70896 40800 70952
rect 37181 70894 40800 70896
rect 37181 70891 37247 70894
rect 39200 70864 40800 70894
rect -800 70818 800 70848
rect 1853 70818 1919 70821
rect -800 70816 1919 70818
rect -800 70760 1858 70816
rect 1914 70760 1919 70816
rect -800 70758 1919 70760
rect -800 70728 800 70758
rect 1853 70755 1919 70758
rect 4208 70752 4528 70753
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 34928 70752 35248 70753
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 70687 35248 70688
rect 37917 70546 37983 70549
rect 39200 70546 40800 70576
rect 37917 70544 40800 70546
rect 37917 70488 37922 70544
rect 37978 70488 40800 70544
rect 37917 70486 40800 70488
rect 37917 70483 37983 70486
rect 39200 70456 40800 70486
rect 19568 70208 19888 70209
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 70143 19888 70144
rect 37181 70002 37247 70005
rect 39200 70002 40800 70032
rect 37181 70000 40800 70002
rect 37181 69944 37186 70000
rect 37242 69944 40800 70000
rect 37181 69942 40800 69944
rect 37181 69939 37247 69942
rect 39200 69912 40800 69942
rect -800 69866 800 69896
rect 1853 69866 1919 69869
rect -800 69864 1919 69866
rect -800 69808 1858 69864
rect 1914 69808 1919 69864
rect -800 69806 1919 69808
rect -800 69776 800 69806
rect 1853 69803 1919 69806
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 34928 69664 35248 69665
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 69599 35248 69600
rect 37181 69594 37247 69597
rect 39200 69594 40800 69624
rect 37181 69592 40800 69594
rect 37181 69536 37186 69592
rect 37242 69536 40800 69592
rect 37181 69534 40800 69536
rect 37181 69531 37247 69534
rect 39200 69504 40800 69534
rect 37917 69186 37983 69189
rect 39200 69186 40800 69216
rect 37917 69184 40800 69186
rect 37917 69128 37922 69184
rect 37978 69128 40800 69184
rect 37917 69126 40800 69128
rect 37917 69123 37983 69126
rect 19568 69120 19888 69121
rect -800 69050 800 69080
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 39200 69096 40800 69126
rect 19568 69055 19888 69056
rect 1853 69050 1919 69053
rect -800 69048 1919 69050
rect -800 68992 1858 69048
rect 1914 68992 1919 69048
rect -800 68990 1919 68992
rect -800 68960 800 68990
rect 1853 68987 1919 68990
rect 37181 68778 37247 68781
rect 39200 68778 40800 68808
rect 37181 68776 40800 68778
rect 37181 68720 37186 68776
rect 37242 68720 40800 68776
rect 37181 68718 40800 68720
rect 37181 68715 37247 68718
rect 39200 68688 40800 68718
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 34928 68576 35248 68577
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 68511 35248 68512
rect 37273 68370 37339 68373
rect 39200 68370 40800 68400
rect 37273 68368 40800 68370
rect 37273 68312 37278 68368
rect 37334 68312 40800 68368
rect 37273 68310 40800 68312
rect 37273 68307 37339 68310
rect 39200 68280 40800 68310
rect -800 68234 800 68264
rect 1853 68234 1919 68237
rect -800 68232 1919 68234
rect -800 68176 1858 68232
rect 1914 68176 1919 68232
rect -800 68174 1919 68176
rect -800 68144 800 68174
rect 1853 68171 1919 68174
rect 19568 68032 19888 68033
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 67967 19888 67968
rect 37181 67962 37247 67965
rect 39200 67962 40800 67992
rect 37181 67960 40800 67962
rect 37181 67904 37186 67960
rect 37242 67904 40800 67960
rect 37181 67902 40800 67904
rect 37181 67899 37247 67902
rect 39200 67872 40800 67902
rect 4208 67488 4528 67489
rect -800 67418 800 67448
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 34928 67488 35248 67489
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 67423 35248 67424
rect 1393 67418 1459 67421
rect -800 67416 1459 67418
rect -800 67360 1398 67416
rect 1454 67360 1459 67416
rect -800 67358 1459 67360
rect -800 67328 800 67358
rect 1393 67355 1459 67358
rect 38929 67418 38995 67421
rect 39200 67418 40800 67448
rect 38929 67416 40800 67418
rect 38929 67360 38934 67416
rect 38990 67360 40800 67416
rect 38929 67358 40800 67360
rect 38929 67355 38995 67358
rect 39200 67328 40800 67358
rect 37273 67010 37339 67013
rect 39200 67010 40800 67040
rect 37273 67008 40800 67010
rect 37273 66952 37278 67008
rect 37334 66952 40800 67008
rect 37273 66950 40800 66952
rect 37273 66947 37339 66950
rect 19568 66944 19888 66945
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 39200 66920 40800 66950
rect 19568 66879 19888 66880
rect -800 66602 800 66632
rect 1393 66602 1459 66605
rect -800 66600 1459 66602
rect -800 66544 1398 66600
rect 1454 66544 1459 66600
rect -800 66542 1459 66544
rect -800 66512 800 66542
rect 1393 66539 1459 66542
rect 37917 66602 37983 66605
rect 39200 66602 40800 66632
rect 37917 66600 40800 66602
rect 37917 66544 37922 66600
rect 37978 66544 40800 66600
rect 37917 66542 40800 66544
rect 37917 66539 37983 66542
rect 39200 66512 40800 66542
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 34928 66400 35248 66401
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 66335 35248 66336
rect 37273 66194 37339 66197
rect 39200 66194 40800 66224
rect 37273 66192 40800 66194
rect 37273 66136 37278 66192
rect 37334 66136 40800 66192
rect 37273 66134 40800 66136
rect 37273 66131 37339 66134
rect 39200 66104 40800 66134
rect 19568 65856 19888 65857
rect -800 65786 800 65816
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 65791 19888 65792
rect 1393 65786 1459 65789
rect -800 65784 1459 65786
rect -800 65728 1398 65784
rect 1454 65728 1459 65784
rect -800 65726 1459 65728
rect -800 65696 800 65726
rect 1393 65723 1459 65726
rect 37181 65786 37247 65789
rect 39200 65786 40800 65816
rect 37181 65784 40800 65786
rect 37181 65728 37186 65784
rect 37242 65728 40800 65784
rect 37181 65726 40800 65728
rect 37181 65723 37247 65726
rect 39200 65696 40800 65726
rect 37917 65378 37983 65381
rect 39200 65378 40800 65408
rect 37917 65376 40800 65378
rect 37917 65320 37922 65376
rect 37978 65320 40800 65376
rect 37917 65318 40800 65320
rect 37917 65315 37983 65318
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 34928 65312 35248 65313
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 39200 65288 40800 65318
rect 34928 65247 35248 65248
rect -800 64970 800 65000
rect 1393 64970 1459 64973
rect -800 64968 1459 64970
rect -800 64912 1398 64968
rect 1454 64912 1459 64968
rect -800 64910 1459 64912
rect -800 64880 800 64910
rect 1393 64907 1459 64910
rect 37181 64834 37247 64837
rect 39200 64834 40800 64864
rect 37181 64832 40800 64834
rect 37181 64776 37186 64832
rect 37242 64776 40800 64832
rect 37181 64774 40800 64776
rect 37181 64771 37247 64774
rect 19568 64768 19888 64769
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 39200 64744 40800 64774
rect 19568 64703 19888 64704
rect 37917 64426 37983 64429
rect 39200 64426 40800 64456
rect 37917 64424 40800 64426
rect 37917 64368 37922 64424
rect 37978 64368 40800 64424
rect 37917 64366 40800 64368
rect 37917 64363 37983 64366
rect 39200 64336 40800 64366
rect 4208 64224 4528 64225
rect -800 64154 800 64184
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 34928 64224 35248 64225
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 64159 35248 64160
rect 1393 64154 1459 64157
rect -800 64152 1459 64154
rect -800 64096 1398 64152
rect 1454 64096 1459 64152
rect -800 64094 1459 64096
rect -800 64064 800 64094
rect 1393 64091 1459 64094
rect 37273 64018 37339 64021
rect 39200 64018 40800 64048
rect 37273 64016 40800 64018
rect 37273 63960 37278 64016
rect 37334 63960 40800 64016
rect 37273 63958 40800 63960
rect 37273 63955 37339 63958
rect 39200 63928 40800 63958
rect 19568 63680 19888 63681
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 63615 19888 63616
rect 37181 63610 37247 63613
rect 39200 63610 40800 63640
rect 37181 63608 40800 63610
rect 37181 63552 37186 63608
rect 37242 63552 40800 63608
rect 37181 63550 40800 63552
rect 37181 63547 37247 63550
rect 39200 63520 40800 63550
rect -800 63338 800 63368
rect 1393 63338 1459 63341
rect -800 63336 1459 63338
rect -800 63280 1398 63336
rect 1454 63280 1459 63336
rect -800 63278 1459 63280
rect -800 63248 800 63278
rect 1393 63275 1459 63278
rect 37917 63202 37983 63205
rect 39200 63202 40800 63232
rect 37917 63200 40800 63202
rect 37917 63144 37922 63200
rect 37978 63144 40800 63200
rect 37917 63142 40800 63144
rect 37917 63139 37983 63142
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 34928 63136 35248 63137
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 39200 63112 40800 63142
rect 34928 63071 35248 63072
rect 37273 62794 37339 62797
rect 39200 62794 40800 62824
rect 37273 62792 40800 62794
rect 37273 62736 37278 62792
rect 37334 62736 40800 62792
rect 37273 62734 40800 62736
rect 37273 62731 37339 62734
rect 39200 62704 40800 62734
rect 19568 62592 19888 62593
rect -800 62522 800 62552
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 62527 19888 62528
rect 1393 62522 1459 62525
rect -800 62520 1459 62522
rect -800 62464 1398 62520
rect 1454 62464 1459 62520
rect -800 62462 1459 62464
rect -800 62432 800 62462
rect 1393 62459 1459 62462
rect 31753 62522 31819 62525
rect 37457 62522 37523 62525
rect 31753 62520 37523 62522
rect 31753 62464 31758 62520
rect 31814 62464 37462 62520
rect 37518 62464 37523 62520
rect 31753 62462 37523 62464
rect 31753 62459 31819 62462
rect 37457 62459 37523 62462
rect 37917 62250 37983 62253
rect 39200 62250 40800 62280
rect 37917 62248 40800 62250
rect 37917 62192 37922 62248
rect 37978 62192 40800 62248
rect 37917 62190 40800 62192
rect 37917 62187 37983 62190
rect 39200 62160 40800 62190
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 34928 62048 35248 62049
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 61983 35248 61984
rect 37273 61842 37339 61845
rect 39200 61842 40800 61872
rect 37273 61840 40800 61842
rect 37273 61784 37278 61840
rect 37334 61784 40800 61840
rect 37273 61782 40800 61784
rect 37273 61779 37339 61782
rect 39200 61752 40800 61782
rect -800 61706 800 61736
rect 1393 61706 1459 61709
rect -800 61704 1459 61706
rect -800 61648 1398 61704
rect 1454 61648 1459 61704
rect -800 61646 1459 61648
rect -800 61616 800 61646
rect 1393 61643 1459 61646
rect 19568 61504 19888 61505
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 61439 19888 61440
rect 37181 61434 37247 61437
rect 39200 61434 40800 61464
rect 37181 61432 40800 61434
rect 37181 61376 37186 61432
rect 37242 61376 40800 61432
rect 37181 61374 40800 61376
rect 37181 61371 37247 61374
rect 39200 61344 40800 61374
rect 37917 61026 37983 61029
rect 39200 61026 40800 61056
rect 37917 61024 40800 61026
rect 37917 60968 37922 61024
rect 37978 60968 40800 61024
rect 37917 60966 40800 60968
rect 37917 60963 37983 60966
rect 4208 60960 4528 60961
rect -800 60890 800 60920
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 34928 60960 35248 60961
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 39200 60936 40800 60966
rect 34928 60895 35248 60896
rect 1393 60890 1459 60893
rect -800 60888 1459 60890
rect -800 60832 1398 60888
rect 1454 60832 1459 60888
rect -800 60830 1459 60832
rect -800 60800 800 60830
rect 1393 60827 1459 60830
rect 37273 60618 37339 60621
rect 39200 60618 40800 60648
rect 37273 60616 40800 60618
rect 37273 60560 37278 60616
rect 37334 60560 40800 60616
rect 37273 60558 40800 60560
rect 37273 60555 37339 60558
rect 39200 60528 40800 60558
rect 19568 60416 19888 60417
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 60351 19888 60352
rect 37181 60210 37247 60213
rect 39200 60210 40800 60240
rect 37181 60208 40800 60210
rect 37181 60152 37186 60208
rect 37242 60152 40800 60208
rect 37181 60150 40800 60152
rect 37181 60147 37247 60150
rect 39200 60120 40800 60150
rect -800 59938 800 59968
rect 1393 59938 1459 59941
rect -800 59936 1459 59938
rect -800 59880 1398 59936
rect 1454 59880 1459 59936
rect -800 59878 1459 59880
rect -800 59848 800 59878
rect 1393 59875 1459 59878
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 34928 59872 35248 59873
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 59807 35248 59808
rect 37917 59666 37983 59669
rect 39200 59666 40800 59696
rect 37917 59664 40800 59666
rect 37917 59608 37922 59664
rect 37978 59608 40800 59664
rect 37917 59606 40800 59608
rect 37917 59603 37983 59606
rect 39200 59576 40800 59606
rect 19568 59328 19888 59329
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 59263 19888 59264
rect 36905 59258 36971 59261
rect 39200 59258 40800 59288
rect 36905 59256 40800 59258
rect 36905 59200 36910 59256
rect 36966 59200 40800 59256
rect 36905 59198 40800 59200
rect 36905 59195 36971 59198
rect 39200 59168 40800 59198
rect -800 59122 800 59152
rect 1393 59122 1459 59125
rect -800 59120 1459 59122
rect -800 59064 1398 59120
rect 1454 59064 1459 59120
rect -800 59062 1459 59064
rect -800 59032 800 59062
rect 1393 59059 1459 59062
rect 36445 58850 36511 58853
rect 39200 58850 40800 58880
rect 36445 58848 40800 58850
rect 36445 58792 36450 58848
rect 36506 58792 40800 58848
rect 36445 58790 40800 58792
rect 36445 58787 36511 58790
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 34928 58784 35248 58785
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 39200 58760 40800 58790
rect 34928 58719 35248 58720
rect 37181 58442 37247 58445
rect 39200 58442 40800 58472
rect 37181 58440 40800 58442
rect 37181 58384 37186 58440
rect 37242 58384 40800 58440
rect 37181 58382 40800 58384
rect 37181 58379 37247 58382
rect 39200 58352 40800 58382
rect -800 58306 800 58336
rect 1393 58306 1459 58309
rect -800 58304 1459 58306
rect -800 58248 1398 58304
rect 1454 58248 1459 58304
rect -800 58246 1459 58248
rect -800 58216 800 58246
rect 1393 58243 1459 58246
rect 19568 58240 19888 58241
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 58175 19888 58176
rect 27429 58034 27495 58037
rect 36445 58034 36511 58037
rect 39200 58034 40800 58064
rect 27429 58032 27538 58034
rect 27429 57976 27434 58032
rect 27490 57976 27538 58032
rect 27429 57971 27538 57976
rect 36445 58032 40800 58034
rect 36445 57976 36450 58032
rect 36506 57976 40800 58032
rect 36445 57974 40800 57976
rect 36445 57971 36511 57974
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect -800 57490 800 57520
rect 1393 57490 1459 57493
rect -800 57488 1459 57490
rect -800 57432 1398 57488
rect 1454 57432 1459 57488
rect -800 57430 1459 57432
rect -800 57400 800 57430
rect 1393 57427 1459 57430
rect 27478 57221 27538 57971
rect 39200 57944 40800 57974
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 37181 57490 37247 57493
rect 39200 57490 40800 57520
rect 37181 57488 40800 57490
rect 37181 57432 37186 57488
rect 37242 57432 40800 57488
rect 37181 57430 40800 57432
rect 37181 57427 37247 57430
rect 39200 57400 40800 57430
rect 27429 57216 27538 57221
rect 27429 57160 27434 57216
rect 27490 57160 27538 57216
rect 27429 57158 27538 57160
rect 27429 57155 27495 57158
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 25589 57082 25655 57085
rect 28625 57082 28691 57085
rect 25589 57080 28691 57082
rect 25589 57024 25594 57080
rect 25650 57024 28630 57080
rect 28686 57024 28691 57080
rect 25589 57022 28691 57024
rect 25589 57019 25655 57022
rect 28625 57019 28691 57022
rect 36445 57082 36511 57085
rect 39200 57082 40800 57112
rect 36445 57080 40800 57082
rect 36445 57024 36450 57080
rect 36506 57024 40800 57080
rect 36445 57022 40800 57024
rect 36445 57019 36511 57022
rect 39200 56992 40800 57022
rect 26233 56946 26299 56949
rect 26509 56946 26575 56949
rect 26233 56944 26575 56946
rect 26233 56888 26238 56944
rect 26294 56888 26514 56944
rect 26570 56888 26575 56944
rect 26233 56886 26575 56888
rect 26233 56883 26299 56886
rect 26509 56883 26575 56886
rect 26509 56810 26575 56813
rect 27521 56810 27587 56813
rect 26509 56808 27587 56810
rect 26509 56752 26514 56808
rect 26570 56752 27526 56808
rect 27582 56752 27587 56808
rect 26509 56750 27587 56752
rect 26509 56747 26575 56750
rect 27521 56747 27587 56750
rect -800 56674 800 56704
rect 1393 56674 1459 56677
rect -800 56672 1459 56674
rect -800 56616 1398 56672
rect 1454 56616 1459 56672
rect -800 56614 1459 56616
rect -800 56584 800 56614
rect 1393 56611 1459 56614
rect 37181 56674 37247 56677
rect 39200 56674 40800 56704
rect 37181 56672 40800 56674
rect 37181 56616 37186 56672
rect 37242 56616 40800 56672
rect 37181 56614 40800 56616
rect 37181 56611 37247 56614
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 39200 56584 40800 56614
rect 34928 56543 35248 56544
rect 36997 56266 37063 56269
rect 39200 56266 40800 56296
rect 36997 56264 40800 56266
rect 36997 56208 37002 56264
rect 37058 56208 40800 56264
rect 36997 56206 40800 56208
rect 36997 56203 37063 56206
rect 39200 56176 40800 56206
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect -800 55858 800 55888
rect 1393 55858 1459 55861
rect -800 55856 1459 55858
rect -800 55800 1398 55856
rect 1454 55800 1459 55856
rect -800 55798 1459 55800
rect -800 55768 800 55798
rect 1393 55795 1459 55798
rect 34881 55858 34947 55861
rect 39200 55858 40800 55888
rect 34881 55856 40800 55858
rect 34881 55800 34886 55856
rect 34942 55800 40800 55856
rect 34881 55798 40800 55800
rect 34881 55795 34947 55798
rect 39200 55768 40800 55798
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 35433 55450 35499 55453
rect 39200 55450 40800 55480
rect 35433 55448 40800 55450
rect 35433 55392 35438 55448
rect 35494 55392 40800 55448
rect 35433 55390 40800 55392
rect 35433 55387 35499 55390
rect 39200 55360 40800 55390
rect -800 55042 800 55072
rect 1393 55042 1459 55045
rect -800 55040 1459 55042
rect -800 54984 1398 55040
rect 1454 54984 1459 55040
rect -800 54982 1459 54984
rect -800 54952 800 54982
rect 1393 54979 1459 54982
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 35801 54906 35867 54909
rect 39200 54906 40800 54936
rect 35801 54904 40800 54906
rect 35801 54848 35806 54904
rect 35862 54848 40800 54904
rect 35801 54846 40800 54848
rect 35801 54843 35867 54846
rect 39200 54816 40800 54846
rect 37089 54498 37155 54501
rect 39200 54498 40800 54528
rect 37089 54496 40800 54498
rect 37089 54440 37094 54496
rect 37150 54440 40800 54496
rect 37089 54438 40800 54440
rect 37089 54435 37155 54438
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 39200 54408 40800 54438
rect 34928 54367 35248 54368
rect -800 54226 800 54256
rect 1393 54226 1459 54229
rect -800 54224 1459 54226
rect -800 54168 1398 54224
rect 1454 54168 1459 54224
rect -800 54166 1459 54168
rect -800 54136 800 54166
rect 1393 54163 1459 54166
rect 35709 54090 35775 54093
rect 39200 54090 40800 54120
rect 35709 54088 40800 54090
rect 35709 54032 35714 54088
rect 35770 54032 40800 54088
rect 35709 54030 40800 54032
rect 35709 54027 35775 54030
rect 39200 54000 40800 54030
rect 19568 53888 19888 53889
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 36721 53682 36787 53685
rect 39200 53682 40800 53712
rect 36721 53680 40800 53682
rect 36721 53624 36726 53680
rect 36782 53624 40800 53680
rect 36721 53622 40800 53624
rect 36721 53619 36787 53622
rect 39200 53592 40800 53622
rect -800 53410 800 53440
rect 1393 53410 1459 53413
rect -800 53408 1459 53410
rect -800 53352 1398 53408
rect 1454 53352 1459 53408
rect -800 53350 1459 53352
rect -800 53320 800 53350
rect 1393 53347 1459 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 53279 35248 53280
rect 37365 53274 37431 53277
rect 39200 53274 40800 53304
rect 37365 53272 40800 53274
rect 37365 53216 37370 53272
rect 37426 53216 40800 53272
rect 37365 53214 40800 53216
rect 37365 53211 37431 53214
rect 39200 53184 40800 53214
rect 36721 53002 36787 53005
rect 37733 53002 37799 53005
rect 36721 53000 37799 53002
rect 36721 52944 36726 53000
rect 36782 52944 37738 53000
rect 37794 52944 37799 53000
rect 36721 52942 37799 52944
rect 36721 52939 36787 52942
rect 37733 52939 37799 52942
rect 35801 52866 35867 52869
rect 39200 52866 40800 52896
rect 35801 52864 40800 52866
rect 35801 52808 35806 52864
rect 35862 52808 40800 52864
rect 35801 52806 40800 52808
rect 35801 52803 35867 52806
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 39200 52776 40800 52806
rect 19568 52735 19888 52736
rect -800 52594 800 52624
rect 1853 52594 1919 52597
rect -800 52592 1919 52594
rect -800 52536 1858 52592
rect 1914 52536 1919 52592
rect -800 52534 1919 52536
rect -800 52504 800 52534
rect 1853 52531 1919 52534
rect 36721 52322 36787 52325
rect 39200 52322 40800 52352
rect 36721 52320 40800 52322
rect 36721 52264 36726 52320
rect 36782 52264 40800 52320
rect 36721 52262 40800 52264
rect 36721 52259 36787 52262
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 39200 52232 40800 52262
rect 34928 52191 35248 52192
rect 37181 51914 37247 51917
rect 39200 51914 40800 51944
rect 37181 51912 40800 51914
rect 37181 51856 37186 51912
rect 37242 51856 40800 51912
rect 37181 51854 40800 51856
rect 37181 51851 37247 51854
rect 39200 51824 40800 51854
rect -800 51778 800 51808
rect 1853 51778 1919 51781
rect -800 51776 1919 51778
rect -800 51720 1858 51776
rect 1914 51720 1919 51776
rect -800 51718 1919 51720
rect -800 51688 800 51718
rect 1853 51715 1919 51718
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 29361 51642 29427 51645
rect 29318 51640 29427 51642
rect 29318 51584 29366 51640
rect 29422 51584 29427 51640
rect 29318 51579 29427 51584
rect 28993 51370 29059 51373
rect 29318 51370 29378 51579
rect 36537 51506 36603 51509
rect 39200 51506 40800 51536
rect 36537 51504 40800 51506
rect 36537 51448 36542 51504
rect 36598 51448 40800 51504
rect 36537 51446 40800 51448
rect 36537 51443 36603 51446
rect 39200 51416 40800 51446
rect 28993 51368 29378 51370
rect 28993 51312 28998 51368
rect 29054 51312 29378 51368
rect 28993 51310 29378 51312
rect 28993 51307 29059 51310
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 51103 35248 51104
rect 37365 51098 37431 51101
rect 39200 51098 40800 51128
rect 37365 51096 40800 51098
rect 37365 51040 37370 51096
rect 37426 51040 40800 51096
rect 37365 51038 40800 51040
rect 37365 51035 37431 51038
rect 39200 51008 40800 51038
rect -800 50962 800 50992
rect 1853 50962 1919 50965
rect -800 50960 1919 50962
rect -800 50904 1858 50960
rect 1914 50904 1919 50960
rect -800 50902 1919 50904
rect -800 50872 800 50902
rect 1853 50899 1919 50902
rect 38101 50690 38167 50693
rect 39200 50690 40800 50720
rect 38101 50688 40800 50690
rect 38101 50632 38106 50688
rect 38162 50632 40800 50688
rect 38101 50630 40800 50632
rect 38101 50627 38167 50630
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 39200 50600 40800 50630
rect 19568 50559 19888 50560
rect 35801 50282 35867 50285
rect 39200 50282 40800 50312
rect 35801 50280 40800 50282
rect 35801 50224 35806 50280
rect 35862 50224 40800 50280
rect 35801 50222 40800 50224
rect 35801 50219 35867 50222
rect 39200 50192 40800 50222
rect 4208 50080 4528 50081
rect -800 50010 800 50040
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 1853 50010 1919 50013
rect -800 50008 1919 50010
rect -800 49952 1858 50008
rect 1914 49952 1919 50008
rect -800 49950 1919 49952
rect -800 49920 800 49950
rect 1853 49947 1919 49950
rect 36261 49738 36327 49741
rect 39200 49738 40800 49768
rect 36261 49736 40800 49738
rect 36261 49680 36266 49736
rect 36322 49680 40800 49736
rect 36261 49678 40800 49680
rect 36261 49675 36327 49678
rect 39200 49648 40800 49678
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 38101 49330 38167 49333
rect 39200 49330 40800 49360
rect 38101 49328 40800 49330
rect 38101 49272 38106 49328
rect 38162 49272 40800 49328
rect 38101 49270 40800 49272
rect 38101 49267 38167 49270
rect 39200 49240 40800 49270
rect -800 49194 800 49224
rect 1853 49194 1919 49197
rect -800 49192 1919 49194
rect -800 49136 1858 49192
rect 1914 49136 1919 49192
rect -800 49134 1919 49136
rect -800 49104 800 49134
rect 1853 49131 1919 49134
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 35525 48922 35591 48925
rect 39200 48922 40800 48952
rect 35525 48920 40800 48922
rect 35525 48864 35530 48920
rect 35586 48864 40800 48920
rect 35525 48862 40800 48864
rect 35525 48859 35591 48862
rect 39200 48832 40800 48862
rect 36261 48786 36327 48789
rect 36126 48784 36327 48786
rect 36126 48728 36266 48784
rect 36322 48728 36327 48784
rect 36126 48726 36327 48728
rect 19977 48514 20043 48517
rect 19977 48512 20178 48514
rect 19977 48456 19982 48512
rect 20038 48456 20178 48512
rect 19977 48454 20178 48456
rect 19977 48451 20043 48454
rect 19568 48448 19888 48449
rect -800 48378 800 48408
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 1853 48378 1919 48381
rect -800 48376 1919 48378
rect -800 48320 1858 48376
rect 1914 48320 1919 48376
rect -800 48318 1919 48320
rect -800 48288 800 48318
rect 1853 48315 1919 48318
rect 19885 48242 19951 48245
rect 20118 48242 20178 48454
rect 19885 48240 20178 48242
rect 19885 48184 19890 48240
rect 19946 48184 20178 48240
rect 19885 48182 20178 48184
rect 19885 48179 19951 48182
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 35893 47698 35959 47701
rect 36126 47698 36186 48726
rect 36261 48723 36327 48726
rect 36261 48514 36327 48517
rect 39200 48514 40800 48544
rect 36261 48512 40800 48514
rect 36261 48456 36266 48512
rect 36322 48456 40800 48512
rect 36261 48454 40800 48456
rect 36261 48451 36327 48454
rect 39200 48424 40800 48454
rect 36353 48106 36419 48109
rect 39200 48106 40800 48136
rect 36353 48104 40800 48106
rect 36353 48048 36358 48104
rect 36414 48048 40800 48104
rect 36353 48046 40800 48048
rect 36353 48043 36419 48046
rect 39200 48016 40800 48046
rect 35893 47696 36186 47698
rect 35893 47640 35898 47696
rect 35954 47640 36186 47696
rect 35893 47638 36186 47640
rect 35893 47635 35959 47638
rect -800 47562 800 47592
rect 1393 47562 1459 47565
rect -800 47560 1459 47562
rect -800 47504 1398 47560
rect 1454 47504 1459 47560
rect -800 47502 1459 47504
rect -800 47472 800 47502
rect 1393 47499 1459 47502
rect 35801 47562 35867 47565
rect 39200 47562 40800 47592
rect 35801 47560 40800 47562
rect 35801 47504 35806 47560
rect 35862 47504 40800 47560
rect 35801 47502 40800 47504
rect 35801 47499 35867 47502
rect 39200 47472 40800 47502
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 35801 47154 35867 47157
rect 39200 47154 40800 47184
rect 35801 47152 40800 47154
rect 35801 47096 35806 47152
rect 35862 47096 40800 47152
rect 35801 47094 40800 47096
rect 35801 47091 35867 47094
rect 39200 47064 40800 47094
rect 4208 46816 4528 46817
rect -800 46746 800 46776
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 1393 46746 1459 46749
rect -800 46744 1459 46746
rect -800 46688 1398 46744
rect 1454 46688 1459 46744
rect -800 46686 1459 46688
rect -800 46656 800 46686
rect 1393 46683 1459 46686
rect 36353 46746 36419 46749
rect 39200 46746 40800 46776
rect 36353 46744 40800 46746
rect 36353 46688 36358 46744
rect 36414 46688 40800 46744
rect 36353 46686 40800 46688
rect 36353 46683 36419 46686
rect 39200 46656 40800 46686
rect 35249 46338 35315 46341
rect 39200 46338 40800 46368
rect 35249 46336 40800 46338
rect 35249 46280 35254 46336
rect 35310 46280 40800 46336
rect 35249 46278 40800 46280
rect 35249 46275 35315 46278
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 39200 46248 40800 46278
rect 19568 46207 19888 46208
rect -800 45930 800 45960
rect 1853 45930 1919 45933
rect -800 45928 1919 45930
rect -800 45872 1858 45928
rect 1914 45872 1919 45928
rect -800 45870 1919 45872
rect -800 45840 800 45870
rect 1853 45867 1919 45870
rect 35709 45930 35775 45933
rect 39200 45930 40800 45960
rect 35709 45928 40800 45930
rect 35709 45872 35714 45928
rect 35770 45872 40800 45928
rect 35709 45870 40800 45872
rect 35709 45867 35775 45870
rect 39200 45840 40800 45870
rect 35709 45794 35775 45797
rect 37181 45794 37247 45797
rect 35709 45792 37247 45794
rect 35709 45736 35714 45792
rect 35770 45736 37186 45792
rect 37242 45736 37247 45792
rect 35709 45734 37247 45736
rect 35709 45731 35775 45734
rect 37181 45731 37247 45734
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 36077 45658 36143 45661
rect 38101 45658 38167 45661
rect 36077 45656 38167 45658
rect 36077 45600 36082 45656
rect 36138 45600 38106 45656
rect 38162 45600 38167 45656
rect 36077 45598 38167 45600
rect 36077 45595 36143 45598
rect 38101 45595 38167 45598
rect 35801 45522 35867 45525
rect 39200 45522 40800 45552
rect 35801 45520 40800 45522
rect 35801 45464 35806 45520
rect 35862 45464 40800 45520
rect 35801 45462 40800 45464
rect 35801 45459 35867 45462
rect 39200 45432 40800 45462
rect 35801 45386 35867 45389
rect 37733 45386 37799 45389
rect 35801 45384 37799 45386
rect 35801 45328 35806 45384
rect 35862 45328 37738 45384
rect 37794 45328 37799 45384
rect 35801 45326 37799 45328
rect 35801 45323 35867 45326
rect 37733 45323 37799 45326
rect 35709 45250 35775 45253
rect 37733 45250 37799 45253
rect 35709 45248 37799 45250
rect 35709 45192 35714 45248
rect 35770 45192 37738 45248
rect 37794 45192 37799 45248
rect 35709 45190 37799 45192
rect 35709 45187 35775 45190
rect 37733 45187 37799 45190
rect 19568 45184 19888 45185
rect -800 45114 800 45144
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 1853 45114 1919 45117
rect -800 45112 1919 45114
rect -800 45056 1858 45112
rect 1914 45056 1919 45112
rect -800 45054 1919 45056
rect -800 45024 800 45054
rect 1853 45051 1919 45054
rect 36077 45114 36143 45117
rect 37365 45114 37431 45117
rect 36077 45112 37431 45114
rect 36077 45056 36082 45112
rect 36138 45056 37370 45112
rect 37426 45056 37431 45112
rect 36077 45054 37431 45056
rect 36077 45051 36143 45054
rect 37365 45051 37431 45054
rect 34513 44978 34579 44981
rect 39200 44978 40800 45008
rect 34513 44976 40800 44978
rect 34513 44920 34518 44976
rect 34574 44920 40800 44976
rect 34513 44918 40800 44920
rect 34513 44915 34579 44918
rect 39200 44888 40800 44918
rect 35801 44706 35867 44709
rect 38009 44706 38075 44709
rect 35801 44704 38075 44706
rect 35801 44648 35806 44704
rect 35862 44648 38014 44704
rect 38070 44648 38075 44704
rect 35801 44646 38075 44648
rect 35801 44643 35867 44646
rect 38009 44643 38075 44646
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 35341 44570 35407 44573
rect 39200 44570 40800 44600
rect 35341 44568 40800 44570
rect 35341 44512 35346 44568
rect 35402 44512 40800 44568
rect 35341 44510 40800 44512
rect 35341 44507 35407 44510
rect 39200 44480 40800 44510
rect 33317 44434 33383 44437
rect 37181 44434 37247 44437
rect 33317 44432 37247 44434
rect 33317 44376 33322 44432
rect 33378 44376 37186 44432
rect 37242 44376 37247 44432
rect 33317 44374 37247 44376
rect 33317 44371 33383 44374
rect 37181 44371 37247 44374
rect -800 44298 800 44328
rect 1853 44298 1919 44301
rect -800 44296 1919 44298
rect -800 44240 1858 44296
rect 1914 44240 1919 44296
rect -800 44238 1919 44240
rect -800 44208 800 44238
rect 1853 44235 1919 44238
rect 35893 44298 35959 44301
rect 36445 44298 36511 44301
rect 35893 44296 36511 44298
rect 35893 44240 35898 44296
rect 35954 44240 36450 44296
rect 36506 44240 36511 44296
rect 35893 44238 36511 44240
rect 35893 44235 35959 44238
rect 36445 44235 36511 44238
rect 35801 44162 35867 44165
rect 39200 44162 40800 44192
rect 35801 44160 40800 44162
rect 35801 44104 35806 44160
rect 35862 44104 40800 44160
rect 35801 44102 40800 44104
rect 35801 44099 35867 44102
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 39200 44072 40800 44102
rect 19568 44031 19888 44032
rect 35341 44026 35407 44029
rect 36537 44026 36603 44029
rect 35341 44024 36603 44026
rect 35341 43968 35346 44024
rect 35402 43968 36542 44024
rect 36598 43968 36603 44024
rect 35341 43966 36603 43968
rect 35341 43963 35407 43966
rect 36537 43963 36603 43966
rect 36813 43890 36879 43893
rect 37549 43890 37615 43893
rect 36813 43888 37615 43890
rect 36813 43832 36818 43888
rect 36874 43832 37554 43888
rect 37610 43832 37615 43888
rect 36813 43830 37615 43832
rect 36813 43827 36879 43830
rect 37549 43827 37615 43830
rect 35065 43754 35131 43757
rect 39200 43754 40800 43784
rect 35065 43752 40800 43754
rect 35065 43696 35070 43752
rect 35126 43696 40800 43752
rect 35065 43694 40800 43696
rect 35065 43691 35131 43694
rect 39200 43664 40800 43694
rect 4208 43552 4528 43553
rect -800 43482 800 43512
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 1853 43482 1919 43485
rect -800 43480 1919 43482
rect -800 43424 1858 43480
rect 1914 43424 1919 43480
rect -800 43422 1919 43424
rect -800 43392 800 43422
rect 1853 43419 1919 43422
rect 28625 43346 28691 43349
rect 28901 43346 28967 43349
rect 28625 43344 28967 43346
rect 28625 43288 28630 43344
rect 28686 43288 28906 43344
rect 28962 43288 28967 43344
rect 28625 43286 28967 43288
rect 28625 43283 28691 43286
rect 28901 43283 28967 43286
rect 34973 43346 35039 43349
rect 39200 43346 40800 43376
rect 34973 43344 40800 43346
rect 34973 43288 34978 43344
rect 35034 43288 40800 43344
rect 34973 43286 40800 43288
rect 34973 43283 35039 43286
rect 39200 43256 40800 43286
rect 31753 43210 31819 43213
rect 38101 43210 38167 43213
rect 31753 43208 38167 43210
rect 31753 43152 31758 43208
rect 31814 43152 38106 43208
rect 38162 43152 38167 43208
rect 31753 43150 38167 43152
rect 31753 43147 31819 43150
rect 38101 43147 38167 43150
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 35709 42938 35775 42941
rect 39200 42938 40800 42968
rect 35709 42936 40800 42938
rect 35709 42880 35714 42936
rect 35770 42880 40800 42936
rect 35709 42878 40800 42880
rect 35709 42875 35775 42878
rect 39200 42848 40800 42878
rect -800 42666 800 42696
rect 1853 42666 1919 42669
rect -800 42664 1919 42666
rect -800 42608 1858 42664
rect 1914 42608 1919 42664
rect -800 42606 1919 42608
rect -800 42576 800 42606
rect 1853 42603 1919 42606
rect 26509 42666 26575 42669
rect 27337 42666 27403 42669
rect 26509 42664 27403 42666
rect 26509 42608 26514 42664
rect 26570 42608 27342 42664
rect 27398 42608 27403 42664
rect 26509 42606 27403 42608
rect 26509 42603 26575 42606
rect 27337 42603 27403 42606
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 35341 42394 35407 42397
rect 39200 42394 40800 42424
rect 35341 42392 40800 42394
rect 35341 42336 35346 42392
rect 35402 42336 40800 42392
rect 35341 42334 40800 42336
rect 35341 42331 35407 42334
rect 39200 42304 40800 42334
rect 34789 41986 34855 41989
rect 39200 41986 40800 42016
rect 34789 41984 40800 41986
rect 34789 41928 34794 41984
rect 34850 41928 40800 41984
rect 34789 41926 40800 41928
rect 34789 41923 34855 41926
rect 19568 41920 19888 41921
rect -800 41850 800 41880
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 39200 41896 40800 41926
rect 19568 41855 19888 41856
rect 1853 41850 1919 41853
rect 28625 41850 28691 41853
rect -800 41848 1919 41850
rect -800 41792 1858 41848
rect 1914 41792 1919 41848
rect -800 41790 1919 41792
rect -800 41760 800 41790
rect 1853 41787 1919 41790
rect 28398 41848 28691 41850
rect 28398 41792 28630 41848
rect 28686 41792 28691 41848
rect 28398 41790 28691 41792
rect 22093 41714 22159 41717
rect 26601 41714 26667 41717
rect 22093 41712 26667 41714
rect 22093 41656 22098 41712
rect 22154 41656 26606 41712
rect 26662 41656 26667 41712
rect 22093 41654 26667 41656
rect 22093 41651 22159 41654
rect 26601 41651 26667 41654
rect 27705 41578 27771 41581
rect 28398 41578 28458 41790
rect 28625 41787 28691 41790
rect 29177 41578 29243 41581
rect 27705 41576 28458 41578
rect 27705 41520 27710 41576
rect 27766 41520 28458 41576
rect 27705 41518 28458 41520
rect 28950 41576 29243 41578
rect 28950 41520 29182 41576
rect 29238 41520 29243 41576
rect 28950 41518 29243 41520
rect 27705 41515 27771 41518
rect 27153 41442 27219 41445
rect 28950 41442 29010 41518
rect 29177 41515 29243 41518
rect 34789 41578 34855 41581
rect 39200 41578 40800 41608
rect 34789 41576 40800 41578
rect 34789 41520 34794 41576
rect 34850 41520 40800 41576
rect 34789 41518 40800 41520
rect 34789 41515 34855 41518
rect 39200 41488 40800 41518
rect 27153 41440 29010 41442
rect 27153 41384 27158 41440
rect 27214 41384 29010 41440
rect 27153 41382 29010 41384
rect 27153 41379 27219 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 26233 41306 26299 41309
rect 27889 41306 27955 41309
rect 26233 41304 27955 41306
rect 26233 41248 26238 41304
rect 26294 41248 27894 41304
rect 27950 41248 27955 41304
rect 26233 41246 27955 41248
rect 26233 41243 26299 41246
rect 27889 41243 27955 41246
rect 34605 41170 34671 41173
rect 39200 41170 40800 41200
rect 34605 41168 40800 41170
rect 34605 41112 34610 41168
rect 34666 41112 40800 41168
rect 34605 41110 40800 41112
rect 34605 41107 34671 41110
rect 39200 41080 40800 41110
rect -800 41034 800 41064
rect 1853 41034 1919 41037
rect -800 41032 1919 41034
rect -800 40976 1858 41032
rect 1914 40976 1919 41032
rect -800 40974 1919 40976
rect -800 40944 800 40974
rect 1853 40971 1919 40974
rect 36169 41034 36235 41037
rect 37089 41034 37155 41037
rect 36169 41032 37155 41034
rect 36169 40976 36174 41032
rect 36230 40976 37094 41032
rect 37150 40976 37155 41032
rect 36169 40974 37155 40976
rect 36169 40971 36235 40974
rect 37089 40971 37155 40974
rect 30741 40898 30807 40901
rect 30925 40898 30991 40901
rect 30741 40896 30991 40898
rect 30741 40840 30746 40896
rect 30802 40840 30930 40896
rect 30986 40840 30991 40896
rect 30741 40838 30991 40840
rect 30741 40835 30807 40838
rect 30925 40835 30991 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 30925 40762 30991 40765
rect 31109 40762 31175 40765
rect 30925 40760 31175 40762
rect 30925 40704 30930 40760
rect 30986 40704 31114 40760
rect 31170 40704 31175 40760
rect 30925 40702 31175 40704
rect 30925 40699 30991 40702
rect 31109 40699 31175 40702
rect 35157 40762 35223 40765
rect 39200 40762 40800 40792
rect 35157 40760 40800 40762
rect 35157 40704 35162 40760
rect 35218 40704 40800 40760
rect 35157 40702 40800 40704
rect 35157 40699 35223 40702
rect 39200 40672 40800 40702
rect 35801 40354 35867 40357
rect 39200 40354 40800 40384
rect 35801 40352 40800 40354
rect 35801 40296 35806 40352
rect 35862 40296 40800 40352
rect 35801 40294 40800 40296
rect 35801 40291 35867 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 39200 40264 40800 40294
rect 34928 40223 35248 40224
rect -800 40082 800 40112
rect 1853 40082 1919 40085
rect -800 40080 1919 40082
rect -800 40024 1858 40080
rect 1914 40024 1919 40080
rect -800 40022 1919 40024
rect -800 39992 800 40022
rect 1853 40019 1919 40022
rect 31109 40082 31175 40085
rect 36905 40082 36971 40085
rect 31109 40080 36971 40082
rect 31109 40024 31114 40080
rect 31170 40024 36910 40080
rect 36966 40024 36971 40080
rect 31109 40022 36971 40024
rect 31109 40019 31175 40022
rect 36905 40019 36971 40022
rect 36077 39946 36143 39949
rect 38101 39946 38167 39949
rect 36077 39944 38167 39946
rect 36077 39888 36082 39944
rect 36138 39888 38106 39944
rect 38162 39888 38167 39944
rect 36077 39886 38167 39888
rect 36077 39883 36143 39886
rect 38101 39883 38167 39886
rect 34605 39810 34671 39813
rect 39200 39810 40800 39840
rect 34605 39808 40800 39810
rect 34605 39752 34610 39808
rect 34666 39752 40800 39808
rect 34605 39750 40800 39752
rect 34605 39747 34671 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 39200 39720 40800 39750
rect 19568 39679 19888 39680
rect 36077 39674 36143 39677
rect 36905 39674 36971 39677
rect 36077 39672 36971 39674
rect 36077 39616 36082 39672
rect 36138 39616 36910 39672
rect 36966 39616 36971 39672
rect 36077 39614 36971 39616
rect 36077 39611 36143 39614
rect 36905 39611 36971 39614
rect 34145 39538 34211 39541
rect 36905 39538 36971 39541
rect 34145 39536 36971 39538
rect 34145 39480 34150 39536
rect 34206 39480 36910 39536
rect 36966 39480 36971 39536
rect 34145 39478 36971 39480
rect 34145 39475 34211 39478
rect 36905 39475 36971 39478
rect 30373 39402 30439 39405
rect 30557 39402 30623 39405
rect 30373 39400 30623 39402
rect 30373 39344 30378 39400
rect 30434 39344 30562 39400
rect 30618 39344 30623 39400
rect 30373 39342 30623 39344
rect 30373 39339 30439 39342
rect 30557 39339 30623 39342
rect 34513 39402 34579 39405
rect 39200 39402 40800 39432
rect 34513 39400 40800 39402
rect 34513 39344 34518 39400
rect 34574 39344 40800 39400
rect 34513 39342 40800 39344
rect 34513 39339 34579 39342
rect 39200 39312 40800 39342
rect -800 39266 800 39296
rect 1853 39266 1919 39269
rect -800 39264 1919 39266
rect -800 39208 1858 39264
rect 1914 39208 1919 39264
rect -800 39206 1919 39208
rect -800 39176 800 39206
rect 1853 39203 1919 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 36537 39130 36603 39133
rect 35574 39128 36603 39130
rect 35574 39072 36542 39128
rect 36598 39072 36603 39128
rect 35574 39070 36603 39072
rect 35574 38997 35634 39070
rect 36537 39067 36603 39070
rect 22829 38994 22895 38997
rect 23013 38994 23079 38997
rect 23289 38994 23355 38997
rect 22829 38992 23355 38994
rect 22829 38936 22834 38992
rect 22890 38936 23018 38992
rect 23074 38936 23294 38992
rect 23350 38936 23355 38992
rect 22829 38934 23355 38936
rect 22829 38931 22895 38934
rect 23013 38931 23079 38934
rect 23289 38931 23355 38934
rect 34329 38994 34395 38997
rect 34973 38994 35039 38997
rect 34329 38992 35039 38994
rect 34329 38936 34334 38992
rect 34390 38936 34978 38992
rect 35034 38936 35039 38992
rect 34329 38934 35039 38936
rect 34329 38931 34395 38934
rect 34973 38931 35039 38934
rect 35525 38992 35634 38997
rect 35525 38936 35530 38992
rect 35586 38936 35634 38992
rect 35525 38934 35634 38936
rect 35709 38994 35775 38997
rect 39200 38994 40800 39024
rect 35709 38992 40800 38994
rect 35709 38936 35714 38992
rect 35770 38936 40800 38992
rect 35709 38934 40800 38936
rect 35525 38931 35591 38934
rect 35709 38931 35775 38934
rect 39200 38904 40800 38934
rect 28901 38858 28967 38861
rect 37273 38858 37339 38861
rect 28901 38856 37339 38858
rect 28901 38800 28906 38856
rect 28962 38800 37278 38856
rect 37334 38800 37339 38856
rect 28901 38798 37339 38800
rect 28901 38795 28967 38798
rect 37273 38795 37339 38798
rect 34329 38722 34395 38725
rect 38101 38722 38167 38725
rect 34329 38720 38167 38722
rect 34329 38664 34334 38720
rect 34390 38664 38106 38720
rect 38162 38664 38167 38720
rect 34329 38662 38167 38664
rect 34329 38659 34395 38662
rect 38101 38659 38167 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 22277 38586 22343 38589
rect 23381 38586 23447 38589
rect 22277 38584 23447 38586
rect 22277 38528 22282 38584
rect 22338 38528 23386 38584
rect 23442 38528 23447 38584
rect 22277 38526 23447 38528
rect 22277 38523 22343 38526
rect 23381 38523 23447 38526
rect 28625 38586 28691 38589
rect 28809 38586 28875 38589
rect 28625 38584 28875 38586
rect 28625 38528 28630 38584
rect 28686 38528 28814 38584
rect 28870 38528 28875 38584
rect 28625 38526 28875 38528
rect 28625 38523 28691 38526
rect 28809 38523 28875 38526
rect 34789 38586 34855 38589
rect 39200 38586 40800 38616
rect 34789 38584 40800 38586
rect 34789 38528 34794 38584
rect 34850 38528 40800 38584
rect 34789 38526 40800 38528
rect 34789 38523 34855 38526
rect 39200 38496 40800 38526
rect -800 38450 800 38480
rect 1853 38450 1919 38453
rect -800 38448 1919 38450
rect -800 38392 1858 38448
rect 1914 38392 1919 38448
rect -800 38390 1919 38392
rect -800 38360 800 38390
rect 1853 38387 1919 38390
rect 23105 38450 23171 38453
rect 27337 38450 27403 38453
rect 23105 38448 27403 38450
rect 23105 38392 23110 38448
rect 23166 38392 27342 38448
rect 27398 38392 27403 38448
rect 23105 38390 27403 38392
rect 23105 38387 23171 38390
rect 27337 38387 27403 38390
rect 36905 38450 36971 38453
rect 37733 38450 37799 38453
rect 36905 38448 37799 38450
rect 36905 38392 36910 38448
rect 36966 38392 37738 38448
rect 37794 38392 37799 38448
rect 36905 38390 37799 38392
rect 36905 38387 36971 38390
rect 37733 38387 37799 38390
rect 22277 38314 22343 38317
rect 23197 38314 23263 38317
rect 22277 38312 23263 38314
rect 22277 38256 22282 38312
rect 22338 38256 23202 38312
rect 23258 38256 23263 38312
rect 22277 38254 23263 38256
rect 22277 38251 22343 38254
rect 23197 38251 23263 38254
rect 25865 38314 25931 38317
rect 28901 38314 28967 38317
rect 38561 38314 38627 38317
rect 25865 38312 28967 38314
rect 25865 38256 25870 38312
rect 25926 38256 28906 38312
rect 28962 38256 28967 38312
rect 25865 38254 28967 38256
rect 25865 38251 25931 38254
rect 28901 38251 28967 38254
rect 29686 38312 38627 38314
rect 29686 38256 38566 38312
rect 38622 38256 38627 38312
rect 29686 38254 38627 38256
rect 29686 38181 29746 38254
rect 38561 38251 38627 38254
rect 29686 38176 29795 38181
rect 29686 38120 29734 38176
rect 29790 38120 29795 38176
rect 29686 38118 29795 38120
rect 29729 38115 29795 38118
rect 35341 38178 35407 38181
rect 39200 38178 40800 38208
rect 35341 38176 40800 38178
rect 35341 38120 35346 38176
rect 35402 38120 40800 38176
rect 35341 38118 40800 38120
rect 35341 38115 35407 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 39200 38088 40800 38118
rect 34928 38047 35248 38048
rect 29913 38042 29979 38045
rect 36905 38042 36971 38045
rect 37917 38042 37983 38045
rect 29913 38040 30298 38042
rect 29913 37984 29918 38040
rect 29974 37984 30298 38040
rect 29913 37982 30298 37984
rect 29913 37979 29979 37982
rect 21909 37906 21975 37909
rect 24209 37906 24275 37909
rect 21909 37904 24275 37906
rect 21909 37848 21914 37904
rect 21970 37848 24214 37904
rect 24270 37848 24275 37904
rect 21909 37846 24275 37848
rect 21909 37843 21975 37846
rect 24209 37843 24275 37846
rect 22277 37770 22343 37773
rect 23381 37770 23447 37773
rect 22277 37768 23447 37770
rect 22277 37712 22282 37768
rect 22338 37712 23386 37768
rect 23442 37712 23447 37768
rect 22277 37710 23447 37712
rect 22277 37707 22343 37710
rect 23381 37707 23447 37710
rect 24485 37770 24551 37773
rect 28441 37770 28507 37773
rect 24485 37768 28507 37770
rect 24485 37712 24490 37768
rect 24546 37712 28446 37768
rect 28502 37712 28507 37768
rect 24485 37710 28507 37712
rect 24485 37707 24551 37710
rect 28441 37707 28507 37710
rect -800 37634 800 37664
rect 1853 37634 1919 37637
rect -800 37632 1919 37634
rect -800 37576 1858 37632
rect 1914 37576 1919 37632
rect -800 37574 1919 37576
rect -800 37544 800 37574
rect 1853 37571 1919 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 30005 37498 30071 37501
rect 29870 37496 30071 37498
rect 29870 37440 30010 37496
rect 30066 37440 30071 37496
rect 29870 37438 30071 37440
rect 29870 37229 29930 37438
rect 30005 37435 30071 37438
rect 29821 37224 29930 37229
rect 29821 37168 29826 37224
rect 29882 37168 29930 37224
rect 29821 37166 29930 37168
rect 29821 37163 29887 37166
rect 30238 37093 30298 37982
rect 36905 38040 37983 38042
rect 36905 37984 36910 38040
rect 36966 37984 37922 38040
rect 37978 37984 37983 38040
rect 36905 37982 37983 37984
rect 36905 37979 36971 37982
rect 37917 37979 37983 37982
rect 30649 37906 30715 37909
rect 30833 37906 30899 37909
rect 30649 37904 30899 37906
rect 30649 37848 30654 37904
rect 30710 37848 30838 37904
rect 30894 37848 30899 37904
rect 30649 37846 30899 37848
rect 30649 37843 30715 37846
rect 30833 37843 30899 37846
rect 36169 37770 36235 37773
rect 39200 37770 40800 37800
rect 36169 37768 40800 37770
rect 36169 37712 36174 37768
rect 36230 37712 40800 37768
rect 36169 37710 40800 37712
rect 36169 37707 36235 37710
rect 39200 37680 40800 37710
rect 35525 37226 35591 37229
rect 39200 37226 40800 37256
rect 35525 37224 40800 37226
rect 35525 37168 35530 37224
rect 35586 37168 40800 37224
rect 35525 37166 40800 37168
rect 35525 37163 35591 37166
rect 39200 37136 40800 37166
rect 30189 37088 30298 37093
rect 36169 37090 36235 37093
rect 30189 37032 30194 37088
rect 30250 37032 30298 37088
rect 30189 37030 30298 37032
rect 36126 37088 36235 37090
rect 36126 37032 36174 37088
rect 36230 37032 36235 37088
rect 30189 37027 30255 37030
rect 36126 37027 36235 37032
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect -800 36818 800 36848
rect 1393 36818 1459 36821
rect -800 36816 1459 36818
rect -800 36760 1398 36816
rect 1454 36760 1459 36816
rect -800 36758 1459 36760
rect -800 36728 800 36758
rect 1393 36755 1459 36758
rect 36126 36546 36186 37027
rect 36353 36818 36419 36821
rect 39200 36818 40800 36848
rect 36353 36816 40800 36818
rect 36353 36760 36358 36816
rect 36414 36760 40800 36816
rect 36353 36758 40800 36760
rect 36353 36755 36419 36758
rect 39200 36728 40800 36758
rect 37365 36546 37431 36549
rect 36126 36544 37431 36546
rect 36126 36488 37370 36544
rect 37426 36488 37431 36544
rect 36126 36486 37431 36488
rect 37365 36483 37431 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 35433 36410 35499 36413
rect 39200 36410 40800 36440
rect 35433 36408 40800 36410
rect 35433 36352 35438 36408
rect 35494 36352 40800 36408
rect 35433 36350 40800 36352
rect 35433 36347 35499 36350
rect 39200 36320 40800 36350
rect 35893 36274 35959 36277
rect 36629 36274 36695 36277
rect 35893 36272 36695 36274
rect 35893 36216 35898 36272
rect 35954 36216 36634 36272
rect 36690 36216 36695 36272
rect 35893 36214 36695 36216
rect 35893 36211 35959 36214
rect 36629 36211 36695 36214
rect 34789 36138 34855 36141
rect 34789 36136 36002 36138
rect 34789 36080 34794 36136
rect 34850 36080 36002 36136
rect 34789 36078 36002 36080
rect 34789 36075 34855 36078
rect -800 36002 800 36032
rect 1393 36002 1459 36005
rect -800 36000 1459 36002
rect -800 35944 1398 36000
rect 1454 35944 1459 36000
rect -800 35942 1459 35944
rect 35942 36002 36002 36078
rect 39200 36002 40800 36032
rect 35942 35942 40800 36002
rect -800 35912 800 35942
rect 1393 35939 1459 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 39200 35912 40800 35942
rect 34928 35871 35248 35872
rect 36445 35866 36511 35869
rect 37457 35866 37523 35869
rect 36445 35864 37523 35866
rect 36445 35808 36450 35864
rect 36506 35808 37462 35864
rect 37518 35808 37523 35864
rect 36445 35806 37523 35808
rect 36445 35803 36511 35806
rect 37457 35803 37523 35806
rect 35525 35730 35591 35733
rect 36353 35730 36419 35733
rect 35525 35728 36419 35730
rect 35525 35672 35530 35728
rect 35586 35672 36358 35728
rect 36414 35672 36419 35728
rect 35525 35670 36419 35672
rect 35525 35667 35591 35670
rect 36353 35667 36419 35670
rect 34789 35594 34855 35597
rect 39200 35594 40800 35624
rect 34789 35592 40800 35594
rect 34789 35536 34794 35592
rect 34850 35536 40800 35592
rect 34789 35534 40800 35536
rect 34789 35531 34855 35534
rect 39200 35504 40800 35534
rect 33317 35458 33383 35461
rect 34329 35458 34395 35461
rect 33317 35456 34395 35458
rect 33317 35400 33322 35456
rect 33378 35400 34334 35456
rect 34390 35400 34395 35456
rect 33317 35398 34395 35400
rect 33317 35395 33383 35398
rect 34329 35395 34395 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect -800 35186 800 35216
rect 1393 35186 1459 35189
rect -800 35184 1459 35186
rect -800 35128 1398 35184
rect 1454 35128 1459 35184
rect -800 35126 1459 35128
rect -800 35096 800 35126
rect 1393 35123 1459 35126
rect 37457 35050 37523 35053
rect 39200 35050 40800 35080
rect 37457 35048 40800 35050
rect 37457 34992 37462 35048
rect 37518 34992 40800 35048
rect 37457 34990 40800 34992
rect 37457 34987 37523 34990
rect 39200 34960 40800 34990
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 35525 34778 35591 34781
rect 36169 34778 36235 34781
rect 35525 34776 36235 34778
rect 35525 34720 35530 34776
rect 35586 34720 36174 34776
rect 36230 34720 36235 34776
rect 35525 34718 36235 34720
rect 35525 34715 35591 34718
rect 36169 34715 36235 34718
rect 34605 34642 34671 34645
rect 39200 34642 40800 34672
rect 34605 34640 40800 34642
rect 34605 34584 34610 34640
rect 34666 34584 40800 34640
rect 34605 34582 40800 34584
rect 34605 34579 34671 34582
rect 39200 34552 40800 34582
rect 24393 34506 24459 34509
rect 28809 34506 28875 34509
rect 24393 34504 28875 34506
rect 24393 34448 24398 34504
rect 24454 34448 28814 34504
rect 28870 34448 28875 34504
rect 24393 34446 28875 34448
rect 24393 34443 24459 34446
rect 28809 34443 28875 34446
rect 35893 34506 35959 34509
rect 36169 34506 36235 34509
rect 35893 34504 36235 34506
rect 35893 34448 35898 34504
rect 35954 34448 36174 34504
rect 36230 34448 36235 34504
rect 35893 34446 36235 34448
rect 35893 34443 35959 34446
rect 36169 34443 36235 34446
rect -800 34370 800 34400
rect 1393 34370 1459 34373
rect -800 34368 1459 34370
rect -800 34312 1398 34368
rect 1454 34312 1459 34368
rect -800 34310 1459 34312
rect -800 34280 800 34310
rect 1393 34307 1459 34310
rect 22277 34370 22343 34373
rect 26877 34370 26943 34373
rect 22277 34368 26943 34370
rect 22277 34312 22282 34368
rect 22338 34312 26882 34368
rect 26938 34312 26943 34368
rect 22277 34310 26943 34312
rect 22277 34307 22343 34310
rect 26877 34307 26943 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 26877 34234 26943 34237
rect 28257 34234 28323 34237
rect 26877 34232 28323 34234
rect 26877 34176 26882 34232
rect 26938 34176 28262 34232
rect 28318 34176 28323 34232
rect 26877 34174 28323 34176
rect 26877 34171 26943 34174
rect 28257 34171 28323 34174
rect 35617 34234 35683 34237
rect 39200 34234 40800 34264
rect 35617 34232 40800 34234
rect 35617 34176 35622 34232
rect 35678 34176 40800 34232
rect 35617 34174 40800 34176
rect 35617 34171 35683 34174
rect 39200 34144 40800 34174
rect 26693 34098 26759 34101
rect 27429 34098 27495 34101
rect 26693 34096 27495 34098
rect 26693 34040 26698 34096
rect 26754 34040 27434 34096
rect 27490 34040 27495 34096
rect 26693 34038 27495 34040
rect 26693 34035 26759 34038
rect 27429 34035 27495 34038
rect 35525 34098 35591 34101
rect 36721 34098 36787 34101
rect 35525 34096 36787 34098
rect 35525 34040 35530 34096
rect 35586 34040 36726 34096
rect 36782 34040 36787 34096
rect 35525 34038 36787 34040
rect 35525 34035 35591 34038
rect 36721 34035 36787 34038
rect 37365 33826 37431 33829
rect 39200 33826 40800 33856
rect 37365 33824 40800 33826
rect 37365 33768 37370 33824
rect 37426 33768 40800 33824
rect 37365 33766 40800 33768
rect 37365 33763 37431 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 39200 33736 40800 33766
rect 34928 33695 35248 33696
rect 28625 33690 28691 33693
rect 28582 33688 28691 33690
rect 28582 33632 28630 33688
rect 28686 33632 28691 33688
rect 28582 33627 28691 33632
rect 35893 33690 35959 33693
rect 36629 33690 36695 33693
rect 35893 33688 36695 33690
rect 35893 33632 35898 33688
rect 35954 33632 36634 33688
rect 36690 33632 36695 33688
rect 35893 33630 36695 33632
rect 35893 33627 35959 33630
rect 36629 33627 36695 33630
rect -800 33554 800 33584
rect 1853 33554 1919 33557
rect -800 33552 1919 33554
rect -800 33496 1858 33552
rect 1914 33496 1919 33552
rect -800 33494 1919 33496
rect -800 33464 800 33494
rect 1853 33491 1919 33494
rect 28582 33421 28642 33627
rect 27613 33418 27679 33421
rect 27613 33416 28458 33418
rect 27613 33360 27618 33416
rect 27674 33360 28458 33416
rect 27613 33358 28458 33360
rect 28582 33416 28691 33421
rect 28582 33360 28630 33416
rect 28686 33360 28691 33416
rect 28582 33358 28691 33360
rect 27613 33355 27679 33358
rect 27981 33282 28047 33285
rect 28398 33282 28458 33358
rect 28625 33355 28691 33358
rect 35433 33418 35499 33421
rect 39200 33418 40800 33448
rect 35433 33416 40800 33418
rect 35433 33360 35438 33416
rect 35494 33360 40800 33416
rect 35433 33358 40800 33360
rect 35433 33355 35499 33358
rect 39200 33328 40800 33358
rect 28533 33282 28599 33285
rect 27981 33280 28320 33282
rect 27981 33224 27986 33280
rect 28042 33224 28320 33280
rect 27981 33222 28320 33224
rect 28398 33280 28599 33282
rect 28398 33224 28538 33280
rect 28594 33224 28599 33280
rect 28398 33222 28599 33224
rect 27981 33219 28047 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 28260 33149 28320 33222
rect 28533 33219 28599 33222
rect 20805 33146 20871 33149
rect 27981 33146 28047 33149
rect 20805 33144 28047 33146
rect 20805 33088 20810 33144
rect 20866 33088 27986 33144
rect 28042 33088 28047 33144
rect 20805 33086 28047 33088
rect 20805 33083 20871 33086
rect 27981 33083 28047 33086
rect 28257 33144 28323 33149
rect 28257 33088 28262 33144
rect 28318 33088 28323 33144
rect 28257 33083 28323 33088
rect 36077 33146 36143 33149
rect 38101 33146 38167 33149
rect 36077 33144 38167 33146
rect 36077 33088 36082 33144
rect 36138 33088 38106 33144
rect 38162 33088 38167 33144
rect 36077 33086 38167 33088
rect 36077 33083 36143 33086
rect 38101 33083 38167 33086
rect 22829 33010 22895 33013
rect 26877 33010 26943 33013
rect 22829 33008 26943 33010
rect 22829 32952 22834 33008
rect 22890 32952 26882 33008
rect 26938 32952 26943 33008
rect 22829 32950 26943 32952
rect 22829 32947 22895 32950
rect 26877 32947 26943 32950
rect 37365 33010 37431 33013
rect 39200 33010 40800 33040
rect 37365 33008 40800 33010
rect 37365 32952 37370 33008
rect 37426 32952 40800 33008
rect 37365 32950 40800 32952
rect 37365 32947 37431 32950
rect 39200 32920 40800 32950
rect 27705 32874 27771 32877
rect 28533 32874 28599 32877
rect 27705 32872 28599 32874
rect 27705 32816 27710 32872
rect 27766 32816 28538 32872
rect 28594 32816 28599 32872
rect 27705 32814 28599 32816
rect 27705 32811 27771 32814
rect 28533 32811 28599 32814
rect -800 32738 800 32768
rect 1393 32738 1459 32741
rect 27981 32738 28047 32741
rect -800 32736 1459 32738
rect -800 32680 1398 32736
rect 1454 32680 1459 32736
rect -800 32678 1459 32680
rect -800 32648 800 32678
rect 1393 32675 1459 32678
rect 27110 32736 28047 32738
rect 27110 32680 27986 32736
rect 28042 32680 28047 32736
rect 27110 32678 28047 32680
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 26969 32602 27035 32605
rect 27110 32602 27170 32678
rect 27981 32675 28047 32678
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 26969 32600 27170 32602
rect 26969 32544 26974 32600
rect 27030 32544 27170 32600
rect 26969 32542 27170 32544
rect 27337 32602 27403 32605
rect 29453 32602 29519 32605
rect 27337 32600 29519 32602
rect 27337 32544 27342 32600
rect 27398 32544 29458 32600
rect 29514 32544 29519 32600
rect 27337 32542 29519 32544
rect 26969 32539 27035 32542
rect 27337 32539 27403 32542
rect 29453 32539 29519 32542
rect 25221 32466 25287 32469
rect 26049 32466 26115 32469
rect 26969 32466 27035 32469
rect 25221 32464 25698 32466
rect 25221 32408 25226 32464
rect 25282 32408 25698 32464
rect 25221 32406 25698 32408
rect 25221 32403 25287 32406
rect 24301 32330 24367 32333
rect 25405 32330 25471 32333
rect 24301 32328 25471 32330
rect 24301 32272 24306 32328
rect 24362 32272 25410 32328
rect 25466 32272 25471 32328
rect 24301 32270 25471 32272
rect 24301 32267 24367 32270
rect 25405 32267 25471 32270
rect 25638 32194 25698 32406
rect 26049 32464 27035 32466
rect 26049 32408 26054 32464
rect 26110 32408 26974 32464
rect 27030 32408 27035 32464
rect 26049 32406 27035 32408
rect 26049 32403 26115 32406
rect 26969 32403 27035 32406
rect 38009 32466 38075 32469
rect 39200 32466 40800 32496
rect 38009 32464 40800 32466
rect 38009 32408 38014 32464
rect 38070 32408 40800 32464
rect 38009 32406 40800 32408
rect 38009 32403 38075 32406
rect 39200 32376 40800 32406
rect 26969 32330 27035 32333
rect 27981 32330 28047 32333
rect 26969 32328 28047 32330
rect 26969 32272 26974 32328
rect 27030 32272 27986 32328
rect 28042 32272 28047 32328
rect 26969 32270 28047 32272
rect 26969 32267 27035 32270
rect 27981 32267 28047 32270
rect 28625 32194 28691 32197
rect 25638 32192 28691 32194
rect 25638 32136 28630 32192
rect 28686 32136 28691 32192
rect 25638 32134 28691 32136
rect 28625 32131 28691 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 23381 32058 23447 32061
rect 26969 32058 27035 32061
rect 23381 32056 27035 32058
rect 23381 32000 23386 32056
rect 23442 32000 26974 32056
rect 27030 32000 27035 32056
rect 23381 31998 27035 32000
rect 23381 31995 23447 31998
rect 26969 31995 27035 31998
rect 35525 32058 35591 32061
rect 39200 32058 40800 32088
rect 35525 32056 40800 32058
rect 35525 32000 35530 32056
rect 35586 32000 40800 32056
rect 35525 31998 40800 32000
rect 35525 31995 35591 31998
rect 39200 31968 40800 31998
rect -800 31922 800 31952
rect 1393 31922 1459 31925
rect -800 31920 1459 31922
rect -800 31864 1398 31920
rect 1454 31864 1459 31920
rect -800 31862 1459 31864
rect -800 31832 800 31862
rect 1393 31859 1459 31862
rect 21633 31922 21699 31925
rect 28349 31922 28415 31925
rect 21633 31920 28415 31922
rect 21633 31864 21638 31920
rect 21694 31864 28354 31920
rect 28410 31864 28415 31920
rect 21633 31862 28415 31864
rect 21633 31859 21699 31862
rect 28349 31859 28415 31862
rect 23565 31650 23631 31653
rect 27889 31650 27955 31653
rect 23565 31648 27955 31650
rect 23565 31592 23570 31648
rect 23626 31592 27894 31648
rect 27950 31592 27955 31648
rect 23565 31590 27955 31592
rect 23565 31587 23631 31590
rect 27889 31587 27955 31590
rect 36905 31650 36971 31653
rect 39200 31650 40800 31680
rect 36905 31648 40800 31650
rect 36905 31592 36910 31648
rect 36966 31592 40800 31648
rect 36905 31590 40800 31592
rect 36905 31587 36971 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 39200 31560 40800 31590
rect 34928 31519 35248 31520
rect 26785 31514 26851 31517
rect 27429 31514 27495 31517
rect 26785 31512 27495 31514
rect 26785 31456 26790 31512
rect 26846 31456 27434 31512
rect 27490 31456 27495 31512
rect 26785 31454 27495 31456
rect 26785 31451 26851 31454
rect 27429 31451 27495 31454
rect 26877 31378 26943 31381
rect 27889 31378 27955 31381
rect 26877 31376 27955 31378
rect 26877 31320 26882 31376
rect 26938 31320 27894 31376
rect 27950 31320 27955 31376
rect 26877 31318 27955 31320
rect 26877 31315 26943 31318
rect 27889 31315 27955 31318
rect 36169 31242 36235 31245
rect 39200 31242 40800 31272
rect 36169 31240 40800 31242
rect 36169 31184 36174 31240
rect 36230 31184 40800 31240
rect 36169 31182 40800 31184
rect 36169 31179 36235 31182
rect 39200 31152 40800 31182
rect -800 31106 800 31136
rect 1393 31106 1459 31109
rect -800 31104 1459 31106
rect -800 31048 1398 31104
rect 1454 31048 1459 31104
rect -800 31046 1459 31048
rect -800 31016 800 31046
rect 1393 31043 1459 31046
rect 22369 31106 22435 31109
rect 29729 31106 29795 31109
rect 22369 31104 29795 31106
rect 22369 31048 22374 31104
rect 22430 31048 29734 31104
rect 29790 31048 29795 31104
rect 22369 31046 29795 31048
rect 22369 31043 22435 31046
rect 29729 31043 29795 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 35801 30834 35867 30837
rect 39200 30834 40800 30864
rect 35801 30832 40800 30834
rect 35801 30776 35806 30832
rect 35862 30776 40800 30832
rect 35801 30774 40800 30776
rect 35801 30771 35867 30774
rect 39200 30744 40800 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 36721 30426 36787 30429
rect 39200 30426 40800 30456
rect 36721 30424 40800 30426
rect 36721 30368 36726 30424
rect 36782 30368 40800 30424
rect 36721 30366 40800 30368
rect 36721 30363 36787 30366
rect 39200 30336 40800 30366
rect 35985 30290 36051 30293
rect 37457 30290 37523 30293
rect 35985 30288 37523 30290
rect 35985 30232 35990 30288
rect 36046 30232 37462 30288
rect 37518 30232 37523 30288
rect 35985 30230 37523 30232
rect 35985 30227 36051 30230
rect 37457 30227 37523 30230
rect -800 30154 800 30184
rect 1393 30154 1459 30157
rect -800 30152 1459 30154
rect -800 30096 1398 30152
rect 1454 30096 1459 30152
rect -800 30094 1459 30096
rect -800 30064 800 30094
rect 1393 30091 1459 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 37365 29882 37431 29885
rect 39200 29882 40800 29912
rect 37365 29880 40800 29882
rect 37365 29824 37370 29880
rect 37426 29824 40800 29880
rect 37365 29822 40800 29824
rect 37365 29819 37431 29822
rect 39200 29792 40800 29822
rect 35801 29474 35867 29477
rect 39200 29474 40800 29504
rect 35801 29472 40800 29474
rect 35801 29416 35806 29472
rect 35862 29416 40800 29472
rect 35801 29414 40800 29416
rect 35801 29411 35867 29414
rect 4208 29408 4528 29409
rect -800 29338 800 29368
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 39200 29384 40800 29414
rect 34928 29343 35248 29344
rect 1393 29338 1459 29341
rect 27613 29338 27679 29341
rect -800 29336 1459 29338
rect -800 29280 1398 29336
rect 1454 29280 1459 29336
rect -800 29278 1459 29280
rect -800 29248 800 29278
rect 1393 29275 1459 29278
rect 27570 29336 27679 29338
rect 27570 29280 27618 29336
rect 27674 29280 27679 29336
rect 27570 29275 27679 29280
rect 22553 29066 22619 29069
rect 25221 29066 25287 29069
rect 22553 29064 25287 29066
rect 22553 29008 22558 29064
rect 22614 29008 25226 29064
rect 25282 29008 25287 29064
rect 22553 29006 25287 29008
rect 22553 29003 22619 29006
rect 25221 29003 25287 29006
rect 22461 28930 22527 28933
rect 24485 28930 24551 28933
rect 22461 28928 24551 28930
rect 22461 28872 22466 28928
rect 22522 28872 24490 28928
rect 24546 28872 24551 28928
rect 22461 28870 24551 28872
rect 22461 28867 22527 28870
rect 24485 28867 24551 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 14457 28794 14523 28797
rect 19977 28794 20043 28797
rect 22277 28794 22343 28797
rect 14457 28792 17970 28794
rect 14457 28736 14462 28792
rect 14518 28736 17970 28792
rect 14457 28734 17970 28736
rect 14457 28731 14523 28734
rect 17910 28658 17970 28734
rect 19977 28792 22343 28794
rect 19977 28736 19982 28792
rect 20038 28736 22282 28792
rect 22338 28736 22343 28792
rect 19977 28734 22343 28736
rect 19977 28731 20043 28734
rect 22277 28731 22343 28734
rect 27570 28661 27630 29275
rect 27797 29202 27863 29205
rect 31937 29202 32003 29205
rect 37181 29202 37247 29205
rect 27797 29200 27906 29202
rect 27797 29144 27802 29200
rect 27858 29144 27906 29200
rect 27797 29139 27906 29144
rect 31937 29200 37247 29202
rect 31937 29144 31942 29200
rect 31998 29144 37186 29200
rect 37242 29144 37247 29200
rect 31937 29142 37247 29144
rect 31937 29139 32003 29142
rect 37181 29139 37247 29142
rect 27846 28933 27906 29139
rect 36077 29066 36143 29069
rect 37457 29066 37523 29069
rect 39200 29066 40800 29096
rect 36077 29064 36186 29066
rect 35893 29010 35959 29013
rect 35893 29008 36002 29010
rect 35893 28952 35898 29008
rect 35954 28952 36002 29008
rect 36077 29008 36082 29064
rect 36138 29008 36186 29064
rect 36077 29003 36186 29008
rect 37457 29064 40800 29066
rect 37457 29008 37462 29064
rect 37518 29008 40800 29064
rect 37457 29006 40800 29008
rect 37457 29003 37523 29006
rect 35893 28947 36002 28952
rect 27797 28928 27906 28933
rect 27797 28872 27802 28928
rect 27858 28872 27906 28928
rect 27797 28870 27906 28872
rect 27797 28867 27863 28870
rect 35942 28794 36002 28947
rect 36126 28930 36186 29003
rect 39200 28976 40800 29006
rect 37825 28930 37891 28933
rect 36126 28928 37891 28930
rect 36126 28872 37830 28928
rect 37886 28872 37891 28928
rect 36126 28870 37891 28872
rect 37825 28867 37891 28870
rect 36353 28794 36419 28797
rect 35942 28792 36419 28794
rect 35942 28736 36358 28792
rect 36414 28736 36419 28792
rect 35942 28734 36419 28736
rect 36353 28731 36419 28734
rect 19609 28658 19675 28661
rect 17910 28656 19675 28658
rect 17910 28600 19614 28656
rect 19670 28600 19675 28656
rect 17910 28598 19675 28600
rect 19609 28595 19675 28598
rect 19793 28658 19859 28661
rect 20069 28658 20135 28661
rect 19793 28656 20135 28658
rect 19793 28600 19798 28656
rect 19854 28600 20074 28656
rect 20130 28600 20135 28656
rect 19793 28598 20135 28600
rect 19793 28595 19859 28598
rect 20069 28595 20135 28598
rect 22553 28658 22619 28661
rect 23565 28658 23631 28661
rect 22553 28656 23631 28658
rect 22553 28600 22558 28656
rect 22614 28600 23570 28656
rect 23626 28600 23631 28656
rect 22553 28598 23631 28600
rect 27570 28656 27679 28661
rect 27570 28600 27618 28656
rect 27674 28600 27679 28656
rect 27570 28598 27679 28600
rect 22553 28595 22619 28598
rect 23565 28595 23631 28598
rect 27613 28595 27679 28598
rect 32305 28658 32371 28661
rect 37365 28658 37431 28661
rect 32305 28656 37431 28658
rect 32305 28600 32310 28656
rect 32366 28600 37370 28656
rect 37426 28600 37431 28656
rect 32305 28598 37431 28600
rect 32305 28595 32371 28598
rect 37365 28595 37431 28598
rect 38101 28658 38167 28661
rect 39200 28658 40800 28688
rect 38101 28656 40800 28658
rect 38101 28600 38106 28656
rect 38162 28600 40800 28656
rect 38101 28598 40800 28600
rect 38101 28595 38167 28598
rect 39200 28568 40800 28598
rect -800 28522 800 28552
rect 1393 28522 1459 28525
rect -800 28520 1459 28522
rect -800 28464 1398 28520
rect 1454 28464 1459 28520
rect -800 28462 1459 28464
rect -800 28432 800 28462
rect 1393 28459 1459 28462
rect 26601 28522 26667 28525
rect 26601 28520 26986 28522
rect 26601 28464 26606 28520
rect 26662 28464 26986 28520
rect 26601 28462 26986 28464
rect 26601 28459 26667 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 18229 28250 18295 28253
rect 22093 28250 22159 28253
rect 18229 28248 22159 28250
rect 18229 28192 18234 28248
rect 18290 28192 22098 28248
rect 22154 28192 22159 28248
rect 18229 28190 22159 28192
rect 26926 28250 26986 28462
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 27061 28250 27127 28253
rect 26926 28248 27127 28250
rect 26926 28192 27066 28248
rect 27122 28192 27127 28248
rect 26926 28190 27127 28192
rect 18229 28187 18295 28190
rect 22093 28187 22159 28190
rect 27061 28187 27127 28190
rect 37181 28250 37247 28253
rect 39200 28250 40800 28280
rect 37181 28248 40800 28250
rect 37181 28192 37186 28248
rect 37242 28192 40800 28248
rect 37181 28190 40800 28192
rect 37181 28187 37247 28190
rect 39200 28160 40800 28190
rect 21449 28114 21515 28117
rect 21449 28112 21650 28114
rect 21449 28056 21454 28112
rect 21510 28056 21650 28112
rect 21449 28054 21650 28056
rect 21449 28051 21515 28054
rect 21590 27842 21650 28054
rect 22001 27842 22067 27845
rect 21590 27840 22067 27842
rect 21590 27784 22006 27840
rect 22062 27784 22067 27840
rect 21590 27782 22067 27784
rect 22001 27779 22067 27782
rect 27061 27842 27127 27845
rect 27705 27842 27771 27845
rect 27061 27840 27771 27842
rect 27061 27784 27066 27840
rect 27122 27784 27710 27840
rect 27766 27784 27771 27840
rect 27061 27782 27771 27784
rect 27061 27779 27127 27782
rect 27705 27779 27771 27782
rect 37457 27842 37523 27845
rect 39200 27842 40800 27872
rect 37457 27840 40800 27842
rect 37457 27784 37462 27840
rect 37518 27784 40800 27840
rect 37457 27782 40800 27784
rect 37457 27779 37523 27782
rect 19568 27776 19888 27777
rect -800 27706 800 27736
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 39200 27752 40800 27782
rect 19568 27711 19888 27712
rect 1853 27706 1919 27709
rect -800 27704 1919 27706
rect -800 27648 1858 27704
rect 1914 27648 1919 27704
rect -800 27646 1919 27648
rect -800 27616 800 27646
rect 1853 27643 1919 27646
rect 20069 27706 20135 27709
rect 24209 27706 24275 27709
rect 20069 27704 24275 27706
rect 20069 27648 20074 27704
rect 20130 27648 24214 27704
rect 24270 27648 24275 27704
rect 20069 27646 24275 27648
rect 20069 27643 20135 27646
rect 24209 27643 24275 27646
rect 19609 27570 19675 27573
rect 23105 27570 23171 27573
rect 23933 27570 23999 27573
rect 19609 27568 23999 27570
rect 19609 27512 19614 27568
rect 19670 27512 23110 27568
rect 23166 27512 23938 27568
rect 23994 27512 23999 27568
rect 19609 27510 23999 27512
rect 19609 27507 19675 27510
rect 23105 27507 23171 27510
rect 23933 27507 23999 27510
rect 37917 27298 37983 27301
rect 39200 27298 40800 27328
rect 37917 27296 40800 27298
rect 37917 27240 37922 27296
rect 37978 27240 40800 27296
rect 37917 27238 40800 27240
rect 37917 27235 37983 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 39200 27208 40800 27238
rect 34928 27167 35248 27168
rect 21817 27026 21883 27029
rect 27429 27026 27495 27029
rect 21817 27024 27495 27026
rect 21817 26968 21822 27024
rect 21878 26968 27434 27024
rect 27490 26968 27495 27024
rect 21817 26966 27495 26968
rect 21817 26963 21883 26966
rect 27429 26963 27495 26966
rect -800 26890 800 26920
rect 1853 26890 1919 26893
rect -800 26888 1919 26890
rect -800 26832 1858 26888
rect 1914 26832 1919 26888
rect -800 26830 1919 26832
rect -800 26800 800 26830
rect 1853 26827 1919 26830
rect 37273 26890 37339 26893
rect 39200 26890 40800 26920
rect 37273 26888 40800 26890
rect 37273 26832 37278 26888
rect 37334 26832 40800 26888
rect 37273 26830 40800 26832
rect 37273 26827 37339 26830
rect 39200 26800 40800 26830
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 21725 26482 21791 26485
rect 22369 26482 22435 26485
rect 21725 26480 22435 26482
rect 21725 26424 21730 26480
rect 21786 26424 22374 26480
rect 22430 26424 22435 26480
rect 21725 26422 22435 26424
rect 21725 26419 21791 26422
rect 22369 26419 22435 26422
rect 37917 26482 37983 26485
rect 39200 26482 40800 26512
rect 37917 26480 40800 26482
rect 37917 26424 37922 26480
rect 37978 26424 40800 26480
rect 37917 26422 40800 26424
rect 37917 26419 37983 26422
rect 39200 26392 40800 26422
rect 4208 26144 4528 26145
rect -800 26074 800 26104
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 1853 26074 1919 26077
rect -800 26072 1919 26074
rect -800 26016 1858 26072
rect 1914 26016 1919 26072
rect -800 26014 1919 26016
rect -800 25984 800 26014
rect 1853 26011 1919 26014
rect 37917 26074 37983 26077
rect 39200 26074 40800 26104
rect 37917 26072 40800 26074
rect 37917 26016 37922 26072
rect 37978 26016 40800 26072
rect 37917 26014 40800 26016
rect 37917 26011 37983 26014
rect 39200 25984 40800 26014
rect 21265 25938 21331 25941
rect 24853 25938 24919 25941
rect 21265 25936 24919 25938
rect 21265 25880 21270 25936
rect 21326 25880 24858 25936
rect 24914 25880 24919 25936
rect 21265 25878 24919 25880
rect 21265 25875 21331 25878
rect 24853 25875 24919 25878
rect 37273 25666 37339 25669
rect 39200 25666 40800 25696
rect 37273 25664 40800 25666
rect 37273 25608 37278 25664
rect 37334 25608 40800 25664
rect 37273 25606 40800 25608
rect 37273 25603 37339 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 39200 25576 40800 25606
rect 19568 25535 19888 25536
rect -800 25258 800 25288
rect 1853 25258 1919 25261
rect -800 25256 1919 25258
rect -800 25200 1858 25256
rect 1914 25200 1919 25256
rect -800 25198 1919 25200
rect -800 25168 800 25198
rect 1853 25195 1919 25198
rect 37181 25258 37247 25261
rect 39200 25258 40800 25288
rect 37181 25256 40800 25258
rect 37181 25200 37186 25256
rect 37242 25200 40800 25256
rect 37181 25198 40800 25200
rect 37181 25195 37247 25198
rect 39200 25168 40800 25198
rect 22001 25122 22067 25125
rect 21590 25120 22067 25122
rect 21590 25064 22006 25120
rect 22062 25064 22067 25120
rect 21590 25062 22067 25064
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 20897 24850 20963 24853
rect 21449 24850 21515 24853
rect 20897 24848 21515 24850
rect 20897 24792 20902 24848
rect 20958 24792 21454 24848
rect 21510 24792 21515 24848
rect 20897 24790 21515 24792
rect 20897 24787 20963 24790
rect 21449 24787 21515 24790
rect 19568 24512 19888 24513
rect -800 24442 800 24472
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 1853 24442 1919 24445
rect -800 24440 1919 24442
rect -800 24384 1858 24440
rect 1914 24384 1919 24440
rect -800 24382 1919 24384
rect -800 24352 800 24382
rect 1853 24379 1919 24382
rect 21590 24306 21650 25062
rect 22001 25059 22067 25062
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 37917 24714 37983 24717
rect 39200 24714 40800 24744
rect 37917 24712 40800 24714
rect 37917 24656 37922 24712
rect 37978 24656 40800 24712
rect 37917 24654 40800 24656
rect 37917 24651 37983 24654
rect 39200 24624 40800 24654
rect 19566 24246 21650 24306
rect 37181 24306 37247 24309
rect 39200 24306 40800 24336
rect 37181 24304 40800 24306
rect 37181 24248 37186 24304
rect 37242 24248 40800 24304
rect 37181 24246 40800 24248
rect 19566 24037 19626 24246
rect 37181 24243 37247 24246
rect 39200 24216 40800 24246
rect 19793 24170 19859 24173
rect 22001 24170 22067 24173
rect 19793 24168 22067 24170
rect 19793 24112 19798 24168
rect 19854 24112 22006 24168
rect 22062 24112 22067 24168
rect 19793 24110 22067 24112
rect 19793 24107 19859 24110
rect 22001 24107 22067 24110
rect 18045 24034 18111 24037
rect 19566 24034 19675 24037
rect 18045 24032 19675 24034
rect 18045 23976 18050 24032
rect 18106 23976 19614 24032
rect 19670 23976 19675 24032
rect 18045 23974 19675 23976
rect 18045 23971 18111 23974
rect 19609 23971 19675 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 18873 23898 18939 23901
rect 19241 23898 19307 23901
rect 18873 23896 19307 23898
rect 18873 23840 18878 23896
rect 18934 23840 19246 23896
rect 19302 23840 19307 23896
rect 18873 23838 19307 23840
rect 18873 23835 18939 23838
rect 19241 23835 19307 23838
rect 19977 23898 20043 23901
rect 24945 23898 25011 23901
rect 19977 23896 25011 23898
rect 19977 23840 19982 23896
rect 20038 23840 24950 23896
rect 25006 23840 25011 23896
rect 19977 23838 25011 23840
rect 19977 23835 20043 23838
rect 24945 23835 25011 23838
rect 37457 23898 37523 23901
rect 39200 23898 40800 23928
rect 37457 23896 40800 23898
rect 37457 23840 37462 23896
rect 37518 23840 40800 23896
rect 37457 23838 40800 23840
rect 37457 23835 37523 23838
rect 39200 23808 40800 23838
rect 17309 23762 17375 23765
rect 20713 23762 20779 23765
rect 17309 23760 20779 23762
rect 17309 23704 17314 23760
rect 17370 23704 20718 23760
rect 20774 23704 20779 23760
rect 17309 23702 20779 23704
rect 17309 23699 17375 23702
rect 20713 23699 20779 23702
rect -800 23626 800 23656
rect 1853 23626 1919 23629
rect -800 23624 1919 23626
rect -800 23568 1858 23624
rect 1914 23568 1919 23624
rect -800 23566 1919 23568
rect -800 23536 800 23566
rect 1853 23563 1919 23566
rect 38101 23490 38167 23493
rect 39200 23490 40800 23520
rect 38101 23488 40800 23490
rect 38101 23432 38106 23488
rect 38162 23432 40800 23488
rect 38101 23430 40800 23432
rect 38101 23427 38167 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 39200 23400 40800 23430
rect 19568 23359 19888 23360
rect 37181 23082 37247 23085
rect 39200 23082 40800 23112
rect 37181 23080 40800 23082
rect 37181 23024 37186 23080
rect 37242 23024 40800 23080
rect 37181 23022 40800 23024
rect 37181 23019 37247 23022
rect 39200 22992 40800 23022
rect 4208 22880 4528 22881
rect -800 22810 800 22840
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 1393 22810 1459 22813
rect -800 22808 1459 22810
rect -800 22752 1398 22808
rect 1454 22752 1459 22808
rect -800 22750 1459 22752
rect -800 22720 800 22750
rect 1393 22747 1459 22750
rect 37273 22538 37339 22541
rect 39200 22538 40800 22568
rect 37273 22536 40800 22538
rect 37273 22480 37278 22536
rect 37334 22480 40800 22536
rect 37273 22478 40800 22480
rect 37273 22475 37339 22478
rect 39200 22448 40800 22478
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 23289 22266 23355 22269
rect 24209 22266 24275 22269
rect 23289 22264 24275 22266
rect 23289 22208 23294 22264
rect 23350 22208 24214 22264
rect 24270 22208 24275 22264
rect 23289 22206 24275 22208
rect 23289 22203 23355 22206
rect 24209 22203 24275 22206
rect 37917 22130 37983 22133
rect 39200 22130 40800 22160
rect 37917 22128 40800 22130
rect 37917 22072 37922 22128
rect 37978 22072 40800 22128
rect 37917 22070 40800 22072
rect 37917 22067 37983 22070
rect 39200 22040 40800 22070
rect -800 21994 800 22024
rect 1393 21994 1459 21997
rect -800 21992 1459 21994
rect -800 21936 1398 21992
rect 1454 21936 1459 21992
rect -800 21934 1459 21936
rect -800 21904 800 21934
rect 1393 21931 1459 21934
rect 17125 21994 17191 21997
rect 18873 21994 18939 21997
rect 17125 21992 18939 21994
rect 17125 21936 17130 21992
rect 17186 21936 18878 21992
rect 18934 21936 18939 21992
rect 17125 21934 18939 21936
rect 17125 21931 17191 21934
rect 18873 21931 18939 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 37181 21722 37247 21725
rect 39200 21722 40800 21752
rect 37181 21720 40800 21722
rect 37181 21664 37186 21720
rect 37242 21664 40800 21720
rect 37181 21662 40800 21664
rect 37181 21659 37247 21662
rect 39200 21632 40800 21662
rect 17677 21586 17743 21589
rect 18597 21586 18663 21589
rect 17677 21584 18663 21586
rect 17677 21528 17682 21584
rect 17738 21528 18602 21584
rect 18658 21528 18663 21584
rect 17677 21526 18663 21528
rect 17677 21523 17743 21526
rect 18597 21523 18663 21526
rect 18781 21586 18847 21589
rect 19241 21586 19307 21589
rect 18781 21584 19307 21586
rect 18781 21528 18786 21584
rect 18842 21528 19246 21584
rect 19302 21528 19307 21584
rect 18781 21526 19307 21528
rect 18781 21523 18847 21526
rect 19241 21523 19307 21526
rect 17125 21450 17191 21453
rect 18505 21450 18571 21453
rect 17125 21448 18571 21450
rect 17125 21392 17130 21448
rect 17186 21392 18510 21448
rect 18566 21392 18571 21448
rect 17125 21390 18571 21392
rect 17125 21387 17191 21390
rect 18505 21387 18571 21390
rect 37273 21314 37339 21317
rect 39200 21314 40800 21344
rect 37273 21312 40800 21314
rect 37273 21256 37278 21312
rect 37334 21256 40800 21312
rect 37273 21254 40800 21256
rect 37273 21251 37339 21254
rect 19568 21248 19888 21249
rect -800 21178 800 21208
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 39200 21224 40800 21254
rect 19568 21183 19888 21184
rect 1393 21178 1459 21181
rect -800 21176 1459 21178
rect -800 21120 1398 21176
rect 1454 21120 1459 21176
rect -800 21118 1459 21120
rect -800 21088 800 21118
rect 1393 21115 1459 21118
rect 37917 20906 37983 20909
rect 39200 20906 40800 20936
rect 37917 20904 40800 20906
rect 37917 20848 37922 20904
rect 37978 20848 40800 20904
rect 37917 20846 40800 20848
rect 37917 20843 37983 20846
rect 39200 20816 40800 20846
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 37273 20498 37339 20501
rect 39200 20498 40800 20528
rect 37273 20496 40800 20498
rect 37273 20440 37278 20496
rect 37334 20440 40800 20496
rect 37273 20438 40800 20440
rect 37273 20435 37339 20438
rect 39200 20408 40800 20438
rect -800 20226 800 20256
rect 1393 20226 1459 20229
rect -800 20224 1459 20226
rect -800 20168 1398 20224
rect 1454 20168 1459 20224
rect -800 20166 1459 20168
rect -800 20136 800 20166
rect 1393 20163 1459 20166
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 37917 19954 37983 19957
rect 39200 19954 40800 19984
rect 37917 19952 40800 19954
rect 37917 19896 37922 19952
rect 37978 19896 40800 19952
rect 37917 19894 40800 19896
rect 37917 19891 37983 19894
rect 39200 19864 40800 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 37917 19546 37983 19549
rect 39200 19546 40800 19576
rect 37917 19544 40800 19546
rect 37917 19488 37922 19544
rect 37978 19488 40800 19544
rect 37917 19486 40800 19488
rect 37917 19483 37983 19486
rect 39200 19456 40800 19486
rect -800 19410 800 19440
rect 1393 19410 1459 19413
rect -800 19408 1459 19410
rect -800 19352 1398 19408
rect 1454 19352 1459 19408
rect -800 19350 1459 19352
rect -800 19320 800 19350
rect 1393 19347 1459 19350
rect 17217 19308 17283 19311
rect 17217 19306 17418 19308
rect 17217 19250 17222 19306
rect 17278 19250 17418 19306
rect 19517 19274 19583 19277
rect 17217 19248 17418 19250
rect 17217 19245 17283 19248
rect 13445 19138 13511 19141
rect 17217 19138 17283 19141
rect 13445 19136 17283 19138
rect 13445 19080 13450 19136
rect 13506 19080 17222 19136
rect 17278 19080 17283 19136
rect 13445 19078 17283 19080
rect 13445 19075 13511 19078
rect 17217 19075 17283 19078
rect 17358 19005 17418 19248
rect 17309 19000 17418 19005
rect 17309 18944 17314 19000
rect 17370 18944 17418 19000
rect 17309 18942 17418 18944
rect 19382 19272 19583 19274
rect 19382 19216 19522 19272
rect 19578 19216 19583 19272
rect 19382 19214 19583 19216
rect 17309 18939 17375 18942
rect 10317 18866 10383 18869
rect 18413 18866 18479 18869
rect 10317 18864 18479 18866
rect 10317 18808 10322 18864
rect 10378 18808 18418 18864
rect 18474 18808 18479 18864
rect 10317 18806 18479 18808
rect 19382 18866 19442 19214
rect 19517 19211 19583 19214
rect 37273 19138 37339 19141
rect 39200 19138 40800 19168
rect 37273 19136 40800 19138
rect 37273 19080 37278 19136
rect 37334 19080 40800 19136
rect 37273 19078 40800 19080
rect 37273 19075 37339 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 39200 19048 40800 19078
rect 19568 19007 19888 19008
rect 19517 18866 19583 18869
rect 19382 18864 19583 18866
rect 19382 18808 19522 18864
rect 19578 18808 19583 18864
rect 19382 18806 19583 18808
rect 10317 18803 10383 18806
rect 18413 18803 18479 18806
rect 19517 18803 19583 18806
rect 37181 18730 37247 18733
rect 39200 18730 40800 18760
rect 37181 18728 40800 18730
rect 37181 18672 37186 18728
rect 37242 18672 40800 18728
rect 37181 18670 40800 18672
rect 37181 18667 37247 18670
rect 39200 18640 40800 18670
rect -800 18594 800 18624
rect 1393 18594 1459 18597
rect -800 18592 1459 18594
rect -800 18536 1398 18592
rect 1454 18536 1459 18592
rect -800 18534 1459 18536
rect -800 18504 800 18534
rect 1393 18531 1459 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 37917 18322 37983 18325
rect 39200 18322 40800 18352
rect 37917 18320 40800 18322
rect 37917 18264 37922 18320
rect 37978 18264 40800 18320
rect 37917 18262 40800 18264
rect 37917 18259 37983 18262
rect 39200 18232 40800 18262
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 37181 17914 37247 17917
rect 39200 17914 40800 17944
rect 37181 17912 40800 17914
rect 37181 17856 37186 17912
rect 37242 17856 40800 17912
rect 37181 17854 40800 17856
rect 37181 17851 37247 17854
rect 39200 17824 40800 17854
rect -800 17778 800 17808
rect 1393 17778 1459 17781
rect -800 17776 1459 17778
rect -800 17720 1398 17776
rect 1454 17720 1459 17776
rect -800 17718 1459 17720
rect -800 17688 800 17718
rect 1393 17715 1459 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 37273 17370 37339 17373
rect 39200 17370 40800 17400
rect 37273 17368 40800 17370
rect 37273 17312 37278 17368
rect 37334 17312 40800 17368
rect 37273 17310 40800 17312
rect 37273 17307 37339 17310
rect 39200 17280 40800 17310
rect -800 16962 800 16992
rect 1393 16962 1459 16965
rect -800 16960 1459 16962
rect -800 16904 1398 16960
rect 1454 16904 1459 16960
rect -800 16902 1459 16904
rect -800 16872 800 16902
rect 1393 16899 1459 16902
rect 37917 16962 37983 16965
rect 39200 16962 40800 16992
rect 37917 16960 40800 16962
rect 37917 16904 37922 16960
rect 37978 16904 40800 16960
rect 37917 16902 40800 16904
rect 37917 16899 37983 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 39200 16872 40800 16902
rect 19568 16831 19888 16832
rect 37181 16554 37247 16557
rect 39200 16554 40800 16584
rect 37181 16552 40800 16554
rect 37181 16496 37186 16552
rect 37242 16496 40800 16552
rect 37181 16494 40800 16496
rect 37181 16491 37247 16494
rect 39200 16464 40800 16494
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect -800 16146 800 16176
rect 1393 16146 1459 16149
rect -800 16144 1459 16146
rect -800 16088 1398 16144
rect 1454 16088 1459 16144
rect -800 16086 1459 16088
rect -800 16056 800 16086
rect 1393 16083 1459 16086
rect 37273 16146 37339 16149
rect 39200 16146 40800 16176
rect 37273 16144 40800 16146
rect 37273 16088 37278 16144
rect 37334 16088 40800 16144
rect 37273 16086 40800 16088
rect 37273 16083 37339 16086
rect 39200 16056 40800 16086
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 37917 15738 37983 15741
rect 39200 15738 40800 15768
rect 37917 15736 40800 15738
rect 37917 15680 37922 15736
rect 37978 15680 40800 15736
rect 37917 15678 40800 15680
rect 37917 15675 37983 15678
rect 39200 15648 40800 15678
rect -800 15330 800 15360
rect 1393 15330 1459 15333
rect -800 15328 1459 15330
rect -800 15272 1398 15328
rect 1454 15272 1459 15328
rect -800 15270 1459 15272
rect -800 15240 800 15270
rect 1393 15267 1459 15270
rect 37181 15330 37247 15333
rect 39200 15330 40800 15360
rect 37181 15328 40800 15330
rect 37181 15272 37186 15328
rect 37242 15272 40800 15328
rect 37181 15270 40800 15272
rect 37181 15267 37247 15270
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 39200 15240 40800 15270
rect 34928 15199 35248 15200
rect 37273 14786 37339 14789
rect 39200 14786 40800 14816
rect 37273 14784 40800 14786
rect 37273 14728 37278 14784
rect 37334 14728 40800 14784
rect 37273 14726 40800 14728
rect 37273 14723 37339 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 39200 14696 40800 14726
rect 19568 14655 19888 14656
rect -800 14514 800 14544
rect 1393 14514 1459 14517
rect -800 14512 1459 14514
rect -800 14456 1398 14512
rect 1454 14456 1459 14512
rect -800 14454 1459 14456
rect -800 14424 800 14454
rect 1393 14451 1459 14454
rect 37917 14378 37983 14381
rect 39200 14378 40800 14408
rect 37917 14376 40800 14378
rect 37917 14320 37922 14376
rect 37978 14320 40800 14376
rect 37917 14318 40800 14320
rect 37917 14315 37983 14318
rect 39200 14288 40800 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 37181 13970 37247 13973
rect 39200 13970 40800 14000
rect 37181 13968 40800 13970
rect 37181 13912 37186 13968
rect 37242 13912 40800 13968
rect 37181 13910 40800 13912
rect 37181 13907 37247 13910
rect 39200 13880 40800 13910
rect -800 13698 800 13728
rect 1393 13698 1459 13701
rect -800 13696 1459 13698
rect -800 13640 1398 13696
rect 1454 13640 1459 13696
rect -800 13638 1459 13640
rect -800 13608 800 13638
rect 1393 13635 1459 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 37917 13562 37983 13565
rect 39200 13562 40800 13592
rect 37917 13560 40800 13562
rect 37917 13504 37922 13560
rect 37978 13504 40800 13560
rect 37917 13502 40800 13504
rect 37917 13499 37983 13502
rect 39200 13472 40800 13502
rect 37181 13154 37247 13157
rect 39200 13154 40800 13184
rect 37181 13152 40800 13154
rect 37181 13096 37186 13152
rect 37242 13096 40800 13152
rect 37181 13094 40800 13096
rect 37181 13091 37247 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 39200 13064 40800 13094
rect 34928 13023 35248 13024
rect -800 12882 800 12912
rect 1393 12882 1459 12885
rect -800 12880 1459 12882
rect -800 12824 1398 12880
rect 1454 12824 1459 12880
rect -800 12822 1459 12824
rect -800 12792 800 12822
rect 1393 12819 1459 12822
rect 37917 12746 37983 12749
rect 39200 12746 40800 12776
rect 37917 12744 40800 12746
rect 37917 12688 37922 12744
rect 37978 12688 40800 12744
rect 37917 12686 40800 12688
rect 37917 12683 37983 12686
rect 39200 12656 40800 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 37181 12202 37247 12205
rect 39200 12202 40800 12232
rect 37181 12200 40800 12202
rect 37181 12144 37186 12200
rect 37242 12144 40800 12200
rect 37181 12142 40800 12144
rect 37181 12139 37247 12142
rect 39200 12112 40800 12142
rect -800 12066 800 12096
rect 1393 12066 1459 12069
rect -800 12064 1459 12066
rect -800 12008 1398 12064
rect 1454 12008 1459 12064
rect -800 12006 1459 12008
rect -800 11976 800 12006
rect 1393 12003 1459 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 37181 11794 37247 11797
rect 39200 11794 40800 11824
rect 37181 11792 40800 11794
rect 37181 11736 37186 11792
rect 37242 11736 40800 11792
rect 37181 11734 40800 11736
rect 37181 11731 37247 11734
rect 39200 11704 40800 11734
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 37917 11386 37983 11389
rect 39200 11386 40800 11416
rect 37917 11384 40800 11386
rect 37917 11328 37922 11384
rect 37978 11328 40800 11384
rect 37917 11326 40800 11328
rect 37917 11323 37983 11326
rect 39200 11296 40800 11326
rect -800 11250 800 11280
rect 1393 11250 1459 11253
rect -800 11248 1459 11250
rect -800 11192 1398 11248
rect 1454 11192 1459 11248
rect -800 11190 1459 11192
rect -800 11160 800 11190
rect 1393 11187 1459 11190
rect 37181 10978 37247 10981
rect 39200 10978 40800 11008
rect 37181 10976 40800 10978
rect 37181 10920 37186 10976
rect 37242 10920 40800 10976
rect 37181 10918 40800 10920
rect 37181 10915 37247 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 39200 10888 40800 10918
rect 34928 10847 35248 10848
rect 37917 10570 37983 10573
rect 39200 10570 40800 10600
rect 37917 10568 40800 10570
rect 37917 10512 37922 10568
rect 37978 10512 40800 10568
rect 37917 10510 40800 10512
rect 37917 10507 37983 10510
rect 39200 10480 40800 10510
rect 19568 10368 19888 10369
rect -800 10298 800 10328
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 1393 10298 1459 10301
rect -800 10296 1459 10298
rect -800 10240 1398 10296
rect 1454 10240 1459 10296
rect -800 10238 1459 10240
rect -800 10208 800 10238
rect 1393 10235 1459 10238
rect 37181 10026 37247 10029
rect 39200 10026 40800 10056
rect 37181 10024 40800 10026
rect 37181 9968 37186 10024
rect 37242 9968 40800 10024
rect 37181 9966 40800 9968
rect 37181 9963 37247 9966
rect 39200 9936 40800 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 37181 9618 37247 9621
rect 39200 9618 40800 9648
rect 37181 9616 40800 9618
rect 37181 9560 37186 9616
rect 37242 9560 40800 9616
rect 37181 9558 40800 9560
rect 37181 9555 37247 9558
rect 39200 9528 40800 9558
rect -800 9482 800 9512
rect 1393 9482 1459 9485
rect -800 9480 1459 9482
rect -800 9424 1398 9480
rect 1454 9424 1459 9480
rect -800 9422 1459 9424
rect -800 9392 800 9422
rect 1393 9419 1459 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 37917 9210 37983 9213
rect 39200 9210 40800 9240
rect 37917 9208 40800 9210
rect 37917 9152 37922 9208
rect 37978 9152 40800 9208
rect 37917 9150 40800 9152
rect 37917 9147 37983 9150
rect 39200 9120 40800 9150
rect 37181 8802 37247 8805
rect 39200 8802 40800 8832
rect 37181 8800 40800 8802
rect 37181 8744 37186 8800
rect 37242 8744 40800 8800
rect 37181 8742 40800 8744
rect 37181 8739 37247 8742
rect 4208 8736 4528 8737
rect -800 8666 800 8696
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 39200 8712 40800 8742
rect 34928 8671 35248 8672
rect 1393 8666 1459 8669
rect -800 8664 1459 8666
rect -800 8608 1398 8664
rect 1454 8608 1459 8664
rect -800 8606 1459 8608
rect -800 8576 800 8606
rect 1393 8603 1459 8606
rect 37917 8394 37983 8397
rect 39200 8394 40800 8424
rect 37917 8392 40800 8394
rect 37917 8336 37922 8392
rect 37978 8336 40800 8392
rect 37917 8334 40800 8336
rect 37917 8331 37983 8334
rect 39200 8304 40800 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 37181 7986 37247 7989
rect 39200 7986 40800 8016
rect 37181 7984 40800 7986
rect 37181 7928 37186 7984
rect 37242 7928 40800 7984
rect 37181 7926 40800 7928
rect 37181 7923 37247 7926
rect 39200 7896 40800 7926
rect -800 7850 800 7880
rect 1393 7850 1459 7853
rect -800 7848 1459 7850
rect -800 7792 1398 7848
rect 1454 7792 1459 7848
rect -800 7790 1459 7792
rect -800 7760 800 7790
rect 1393 7787 1459 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 37181 7442 37247 7445
rect 39200 7442 40800 7472
rect 37181 7440 40800 7442
rect 37181 7384 37186 7440
rect 37242 7384 40800 7440
rect 37181 7382 40800 7384
rect 37181 7379 37247 7382
rect 39200 7352 40800 7382
rect 19568 7104 19888 7105
rect -800 7034 800 7064
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 1393 7034 1459 7037
rect -800 7032 1459 7034
rect -800 6976 1398 7032
rect 1454 6976 1459 7032
rect -800 6974 1459 6976
rect -800 6944 800 6974
rect 1393 6971 1459 6974
rect 37917 7034 37983 7037
rect 39200 7034 40800 7064
rect 37917 7032 40800 7034
rect 37917 6976 37922 7032
rect 37978 6976 40800 7032
rect 37917 6974 40800 6976
rect 37917 6971 37983 6974
rect 39200 6944 40800 6974
rect 37181 6626 37247 6629
rect 39200 6626 40800 6656
rect 37181 6624 40800 6626
rect 37181 6568 37186 6624
rect 37242 6568 40800 6624
rect 37181 6566 40800 6568
rect 37181 6563 37247 6566
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 39200 6536 40800 6566
rect 34928 6495 35248 6496
rect -800 6218 800 6248
rect 1393 6218 1459 6221
rect -800 6216 1459 6218
rect -800 6160 1398 6216
rect 1454 6160 1459 6216
rect -800 6158 1459 6160
rect -800 6128 800 6158
rect 1393 6155 1459 6158
rect 37917 6218 37983 6221
rect 39200 6218 40800 6248
rect 37917 6216 40800 6218
rect 37917 6160 37922 6216
rect 37978 6160 40800 6216
rect 37917 6158 40800 6160
rect 37917 6155 37983 6158
rect 39200 6128 40800 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 37181 5810 37247 5813
rect 39200 5810 40800 5840
rect 37181 5808 40800 5810
rect 37181 5752 37186 5808
rect 37242 5752 40800 5808
rect 37181 5750 40800 5752
rect 37181 5747 37247 5750
rect 39200 5720 40800 5750
rect 4208 5472 4528 5473
rect -800 5402 800 5432
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 2037 5402 2103 5405
rect -800 5400 2103 5402
rect -800 5344 2042 5400
rect 2098 5344 2103 5400
rect -800 5342 2103 5344
rect -800 5312 800 5342
rect 2037 5339 2103 5342
rect 37181 5402 37247 5405
rect 39200 5402 40800 5432
rect 37181 5400 40800 5402
rect 37181 5344 37186 5400
rect 37242 5344 40800 5400
rect 37181 5342 40800 5344
rect 37181 5339 37247 5342
rect 39200 5312 40800 5342
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 37917 4858 37983 4861
rect 39200 4858 40800 4888
rect 37917 4856 40800 4858
rect 37917 4800 37922 4856
rect 37978 4800 40800 4856
rect 37917 4798 40800 4800
rect 37917 4795 37983 4798
rect 39200 4768 40800 4798
rect -800 4586 800 4616
rect 1393 4586 1459 4589
rect -800 4584 1459 4586
rect -800 4528 1398 4584
rect 1454 4528 1459 4584
rect -800 4526 1459 4528
rect -800 4496 800 4526
rect 1393 4523 1459 4526
rect 37181 4450 37247 4453
rect 39200 4450 40800 4480
rect 37181 4448 40800 4450
rect 37181 4392 37186 4448
rect 37242 4392 40800 4448
rect 37181 4390 40800 4392
rect 37181 4387 37247 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 39200 4360 40800 4390
rect 34928 4319 35248 4320
rect 37089 4042 37155 4045
rect 39200 4042 40800 4072
rect 37089 4040 40800 4042
rect 37089 3984 37094 4040
rect 37150 3984 40800 4040
rect 37089 3982 40800 3984
rect 37089 3979 37155 3982
rect 39200 3952 40800 3982
rect 19568 3840 19888 3841
rect -800 3770 800 3800
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 2773 3770 2839 3773
rect -800 3768 2839 3770
rect -800 3712 2778 3768
rect 2834 3712 2839 3768
rect -800 3710 2839 3712
rect -800 3680 800 3710
rect 2773 3707 2839 3710
rect 35801 3634 35867 3637
rect 39200 3634 40800 3664
rect 35801 3632 40800 3634
rect 35801 3576 35806 3632
rect 35862 3576 40800 3632
rect 35801 3574 40800 3576
rect 35801 3571 35867 3574
rect 39200 3544 40800 3574
rect 22185 3498 22251 3501
rect 24393 3498 24459 3501
rect 22185 3496 24459 3498
rect 22185 3440 22190 3496
rect 22246 3440 24398 3496
rect 24454 3440 24459 3496
rect 22185 3438 24459 3440
rect 22185 3435 22251 3438
rect 24393 3435 24459 3438
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 36629 3226 36695 3229
rect 39200 3226 40800 3256
rect 36629 3224 40800 3226
rect 36629 3168 36634 3224
rect 36690 3168 40800 3224
rect 36629 3166 40800 3168
rect 36629 3163 36695 3166
rect 39200 3136 40800 3166
rect 26141 3090 26207 3093
rect 28441 3090 28507 3093
rect 26141 3088 28507 3090
rect 26141 3032 26146 3088
rect 26202 3032 28446 3088
rect 28502 3032 28507 3088
rect 26141 3030 28507 3032
rect 26141 3027 26207 3030
rect 28441 3027 28507 3030
rect -800 2954 800 2984
rect 1301 2954 1367 2957
rect -800 2952 1367 2954
rect -800 2896 1306 2952
rect 1362 2896 1367 2952
rect -800 2894 1367 2896
rect -800 2864 800 2894
rect 1301 2891 1367 2894
rect 33685 2818 33751 2821
rect 34421 2818 34487 2821
rect 33685 2816 34487 2818
rect 33685 2760 33690 2816
rect 33746 2760 34426 2816
rect 34482 2760 34487 2816
rect 33685 2758 34487 2760
rect 33685 2755 33751 2758
rect 34421 2755 34487 2758
rect 36537 2818 36603 2821
rect 39200 2818 40800 2848
rect 36537 2816 40800 2818
rect 36537 2760 36542 2816
rect 36598 2760 40800 2816
rect 36537 2758 40800 2760
rect 36537 2755 36603 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 39200 2728 40800 2758
rect 19568 2687 19888 2688
rect 36445 2274 36511 2277
rect 39200 2274 40800 2304
rect 36445 2272 40800 2274
rect 36445 2216 36450 2272
rect 36506 2216 40800 2272
rect 36445 2214 40800 2216
rect 36445 2211 36511 2214
rect 4208 2208 4528 2209
rect -800 2138 800 2168
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 39200 2184 40800 2214
rect 34928 2143 35248 2144
rect 3325 2138 3391 2141
rect -800 2136 3391 2138
rect -800 2080 3330 2136
rect 3386 2080 3391 2136
rect -800 2078 3391 2080
rect -800 2048 800 2078
rect 3325 2075 3391 2078
rect 36813 1866 36879 1869
rect 39200 1866 40800 1896
rect 36813 1864 40800 1866
rect 36813 1808 36818 1864
rect 36874 1808 40800 1864
rect 36813 1806 40800 1808
rect 36813 1803 36879 1806
rect 39200 1776 40800 1806
rect 38101 1458 38167 1461
rect 39200 1458 40800 1488
rect 38101 1456 40800 1458
rect 38101 1400 38106 1456
rect 38162 1400 40800 1456
rect 38101 1398 40800 1400
rect 38101 1395 38167 1398
rect 39200 1368 40800 1398
rect -800 1322 800 1352
rect 3049 1322 3115 1325
rect -800 1320 3115 1322
rect -800 1264 3054 1320
rect 3110 1264 3115 1320
rect -800 1262 3115 1264
rect -800 1232 800 1262
rect 3049 1259 3115 1262
rect 37181 1050 37247 1053
rect 39200 1050 40800 1080
rect 37181 1048 40800 1050
rect 37181 992 37186 1048
rect 37242 992 40800 1048
rect 37181 990 40800 992
rect 37181 987 37247 990
rect 39200 960 40800 990
rect 36721 642 36787 645
rect 39200 642 40800 672
rect 36721 640 40800 642
rect 36721 584 36726 640
rect 36782 584 40800 640
rect 36721 582 40800 584
rect 36721 579 36787 582
rect 39200 552 40800 582
rect -800 506 800 536
rect 2773 506 2839 509
rect -800 504 2839 506
rect -800 448 2778 504
rect 2834 448 2839 504
rect -800 446 2839 448
rect -800 416 800 446
rect 2773 443 2839 446
rect 37917 234 37983 237
rect 39200 234 40800 264
rect 37917 232 40800 234
rect 37917 176 37922 232
rect 37978 176 40800 232
rect 37917 174 40800 176
rect 37917 171 37983 174
rect 39200 144 40800 174
<< via3 >>
rect 4216 117532 4280 117536
rect 4216 117476 4220 117532
rect 4220 117476 4276 117532
rect 4276 117476 4280 117532
rect 4216 117472 4280 117476
rect 4296 117532 4360 117536
rect 4296 117476 4300 117532
rect 4300 117476 4356 117532
rect 4356 117476 4360 117532
rect 4296 117472 4360 117476
rect 4376 117532 4440 117536
rect 4376 117476 4380 117532
rect 4380 117476 4436 117532
rect 4436 117476 4440 117532
rect 4376 117472 4440 117476
rect 4456 117532 4520 117536
rect 4456 117476 4460 117532
rect 4460 117476 4516 117532
rect 4516 117476 4520 117532
rect 4456 117472 4520 117476
rect 34936 117532 35000 117536
rect 34936 117476 34940 117532
rect 34940 117476 34996 117532
rect 34996 117476 35000 117532
rect 34936 117472 35000 117476
rect 35016 117532 35080 117536
rect 35016 117476 35020 117532
rect 35020 117476 35076 117532
rect 35076 117476 35080 117532
rect 35016 117472 35080 117476
rect 35096 117532 35160 117536
rect 35096 117476 35100 117532
rect 35100 117476 35156 117532
rect 35156 117476 35160 117532
rect 35096 117472 35160 117476
rect 35176 117532 35240 117536
rect 35176 117476 35180 117532
rect 35180 117476 35236 117532
rect 35236 117476 35240 117532
rect 35176 117472 35240 117476
rect 19576 116988 19640 116992
rect 19576 116932 19580 116988
rect 19580 116932 19636 116988
rect 19636 116932 19640 116988
rect 19576 116928 19640 116932
rect 19656 116988 19720 116992
rect 19656 116932 19660 116988
rect 19660 116932 19716 116988
rect 19716 116932 19720 116988
rect 19656 116928 19720 116932
rect 19736 116988 19800 116992
rect 19736 116932 19740 116988
rect 19740 116932 19796 116988
rect 19796 116932 19800 116988
rect 19736 116928 19800 116932
rect 19816 116988 19880 116992
rect 19816 116932 19820 116988
rect 19820 116932 19876 116988
rect 19876 116932 19880 116988
rect 19816 116928 19880 116932
rect 4216 116444 4280 116448
rect 4216 116388 4220 116444
rect 4220 116388 4276 116444
rect 4276 116388 4280 116444
rect 4216 116384 4280 116388
rect 4296 116444 4360 116448
rect 4296 116388 4300 116444
rect 4300 116388 4356 116444
rect 4356 116388 4360 116444
rect 4296 116384 4360 116388
rect 4376 116444 4440 116448
rect 4376 116388 4380 116444
rect 4380 116388 4436 116444
rect 4436 116388 4440 116444
rect 4376 116384 4440 116388
rect 4456 116444 4520 116448
rect 4456 116388 4460 116444
rect 4460 116388 4516 116444
rect 4516 116388 4520 116444
rect 4456 116384 4520 116388
rect 34936 116444 35000 116448
rect 34936 116388 34940 116444
rect 34940 116388 34996 116444
rect 34996 116388 35000 116444
rect 34936 116384 35000 116388
rect 35016 116444 35080 116448
rect 35016 116388 35020 116444
rect 35020 116388 35076 116444
rect 35076 116388 35080 116444
rect 35016 116384 35080 116388
rect 35096 116444 35160 116448
rect 35096 116388 35100 116444
rect 35100 116388 35156 116444
rect 35156 116388 35160 116444
rect 35096 116384 35160 116388
rect 35176 116444 35240 116448
rect 35176 116388 35180 116444
rect 35180 116388 35236 116444
rect 35236 116388 35240 116444
rect 35176 116384 35240 116388
rect 19576 115900 19640 115904
rect 19576 115844 19580 115900
rect 19580 115844 19636 115900
rect 19636 115844 19640 115900
rect 19576 115840 19640 115844
rect 19656 115900 19720 115904
rect 19656 115844 19660 115900
rect 19660 115844 19716 115900
rect 19716 115844 19720 115900
rect 19656 115840 19720 115844
rect 19736 115900 19800 115904
rect 19736 115844 19740 115900
rect 19740 115844 19796 115900
rect 19796 115844 19800 115900
rect 19736 115840 19800 115844
rect 19816 115900 19880 115904
rect 19816 115844 19820 115900
rect 19820 115844 19876 115900
rect 19876 115844 19880 115900
rect 19816 115840 19880 115844
rect 4216 115356 4280 115360
rect 4216 115300 4220 115356
rect 4220 115300 4276 115356
rect 4276 115300 4280 115356
rect 4216 115296 4280 115300
rect 4296 115356 4360 115360
rect 4296 115300 4300 115356
rect 4300 115300 4356 115356
rect 4356 115300 4360 115356
rect 4296 115296 4360 115300
rect 4376 115356 4440 115360
rect 4376 115300 4380 115356
rect 4380 115300 4436 115356
rect 4436 115300 4440 115356
rect 4376 115296 4440 115300
rect 4456 115356 4520 115360
rect 4456 115300 4460 115356
rect 4460 115300 4516 115356
rect 4516 115300 4520 115356
rect 4456 115296 4520 115300
rect 34936 115356 35000 115360
rect 34936 115300 34940 115356
rect 34940 115300 34996 115356
rect 34996 115300 35000 115356
rect 34936 115296 35000 115300
rect 35016 115356 35080 115360
rect 35016 115300 35020 115356
rect 35020 115300 35076 115356
rect 35076 115300 35080 115356
rect 35016 115296 35080 115300
rect 35096 115356 35160 115360
rect 35096 115300 35100 115356
rect 35100 115300 35156 115356
rect 35156 115300 35160 115356
rect 35096 115296 35160 115300
rect 35176 115356 35240 115360
rect 35176 115300 35180 115356
rect 35180 115300 35236 115356
rect 35236 115300 35240 115356
rect 35176 115296 35240 115300
rect 19576 114812 19640 114816
rect 19576 114756 19580 114812
rect 19580 114756 19636 114812
rect 19636 114756 19640 114812
rect 19576 114752 19640 114756
rect 19656 114812 19720 114816
rect 19656 114756 19660 114812
rect 19660 114756 19716 114812
rect 19716 114756 19720 114812
rect 19656 114752 19720 114756
rect 19736 114812 19800 114816
rect 19736 114756 19740 114812
rect 19740 114756 19796 114812
rect 19796 114756 19800 114812
rect 19736 114752 19800 114756
rect 19816 114812 19880 114816
rect 19816 114756 19820 114812
rect 19820 114756 19876 114812
rect 19876 114756 19880 114812
rect 19816 114752 19880 114756
rect 4216 114268 4280 114272
rect 4216 114212 4220 114268
rect 4220 114212 4276 114268
rect 4276 114212 4280 114268
rect 4216 114208 4280 114212
rect 4296 114268 4360 114272
rect 4296 114212 4300 114268
rect 4300 114212 4356 114268
rect 4356 114212 4360 114268
rect 4296 114208 4360 114212
rect 4376 114268 4440 114272
rect 4376 114212 4380 114268
rect 4380 114212 4436 114268
rect 4436 114212 4440 114268
rect 4376 114208 4440 114212
rect 4456 114268 4520 114272
rect 4456 114212 4460 114268
rect 4460 114212 4516 114268
rect 4516 114212 4520 114268
rect 4456 114208 4520 114212
rect 34936 114268 35000 114272
rect 34936 114212 34940 114268
rect 34940 114212 34996 114268
rect 34996 114212 35000 114268
rect 34936 114208 35000 114212
rect 35016 114268 35080 114272
rect 35016 114212 35020 114268
rect 35020 114212 35076 114268
rect 35076 114212 35080 114268
rect 35016 114208 35080 114212
rect 35096 114268 35160 114272
rect 35096 114212 35100 114268
rect 35100 114212 35156 114268
rect 35156 114212 35160 114268
rect 35096 114208 35160 114212
rect 35176 114268 35240 114272
rect 35176 114212 35180 114268
rect 35180 114212 35236 114268
rect 35236 114212 35240 114268
rect 35176 114208 35240 114212
rect 19576 113724 19640 113728
rect 19576 113668 19580 113724
rect 19580 113668 19636 113724
rect 19636 113668 19640 113724
rect 19576 113664 19640 113668
rect 19656 113724 19720 113728
rect 19656 113668 19660 113724
rect 19660 113668 19716 113724
rect 19716 113668 19720 113724
rect 19656 113664 19720 113668
rect 19736 113724 19800 113728
rect 19736 113668 19740 113724
rect 19740 113668 19796 113724
rect 19796 113668 19800 113724
rect 19736 113664 19800 113668
rect 19816 113724 19880 113728
rect 19816 113668 19820 113724
rect 19820 113668 19876 113724
rect 19876 113668 19880 113724
rect 19816 113664 19880 113668
rect 4216 113180 4280 113184
rect 4216 113124 4220 113180
rect 4220 113124 4276 113180
rect 4276 113124 4280 113180
rect 4216 113120 4280 113124
rect 4296 113180 4360 113184
rect 4296 113124 4300 113180
rect 4300 113124 4356 113180
rect 4356 113124 4360 113180
rect 4296 113120 4360 113124
rect 4376 113180 4440 113184
rect 4376 113124 4380 113180
rect 4380 113124 4436 113180
rect 4436 113124 4440 113180
rect 4376 113120 4440 113124
rect 4456 113180 4520 113184
rect 4456 113124 4460 113180
rect 4460 113124 4516 113180
rect 4516 113124 4520 113180
rect 4456 113120 4520 113124
rect 34936 113180 35000 113184
rect 34936 113124 34940 113180
rect 34940 113124 34996 113180
rect 34996 113124 35000 113180
rect 34936 113120 35000 113124
rect 35016 113180 35080 113184
rect 35016 113124 35020 113180
rect 35020 113124 35076 113180
rect 35076 113124 35080 113180
rect 35016 113120 35080 113124
rect 35096 113180 35160 113184
rect 35096 113124 35100 113180
rect 35100 113124 35156 113180
rect 35156 113124 35160 113180
rect 35096 113120 35160 113124
rect 35176 113180 35240 113184
rect 35176 113124 35180 113180
rect 35180 113124 35236 113180
rect 35236 113124 35240 113180
rect 35176 113120 35240 113124
rect 19576 112636 19640 112640
rect 19576 112580 19580 112636
rect 19580 112580 19636 112636
rect 19636 112580 19640 112636
rect 19576 112576 19640 112580
rect 19656 112636 19720 112640
rect 19656 112580 19660 112636
rect 19660 112580 19716 112636
rect 19716 112580 19720 112636
rect 19656 112576 19720 112580
rect 19736 112636 19800 112640
rect 19736 112580 19740 112636
rect 19740 112580 19796 112636
rect 19796 112580 19800 112636
rect 19736 112576 19800 112580
rect 19816 112636 19880 112640
rect 19816 112580 19820 112636
rect 19820 112580 19876 112636
rect 19876 112580 19880 112636
rect 19816 112576 19880 112580
rect 4216 112092 4280 112096
rect 4216 112036 4220 112092
rect 4220 112036 4276 112092
rect 4276 112036 4280 112092
rect 4216 112032 4280 112036
rect 4296 112092 4360 112096
rect 4296 112036 4300 112092
rect 4300 112036 4356 112092
rect 4356 112036 4360 112092
rect 4296 112032 4360 112036
rect 4376 112092 4440 112096
rect 4376 112036 4380 112092
rect 4380 112036 4436 112092
rect 4436 112036 4440 112092
rect 4376 112032 4440 112036
rect 4456 112092 4520 112096
rect 4456 112036 4460 112092
rect 4460 112036 4516 112092
rect 4516 112036 4520 112092
rect 4456 112032 4520 112036
rect 34936 112092 35000 112096
rect 34936 112036 34940 112092
rect 34940 112036 34996 112092
rect 34996 112036 35000 112092
rect 34936 112032 35000 112036
rect 35016 112092 35080 112096
rect 35016 112036 35020 112092
rect 35020 112036 35076 112092
rect 35076 112036 35080 112092
rect 35016 112032 35080 112036
rect 35096 112092 35160 112096
rect 35096 112036 35100 112092
rect 35100 112036 35156 112092
rect 35156 112036 35160 112092
rect 35096 112032 35160 112036
rect 35176 112092 35240 112096
rect 35176 112036 35180 112092
rect 35180 112036 35236 112092
rect 35236 112036 35240 112092
rect 35176 112032 35240 112036
rect 19576 111548 19640 111552
rect 19576 111492 19580 111548
rect 19580 111492 19636 111548
rect 19636 111492 19640 111548
rect 19576 111488 19640 111492
rect 19656 111548 19720 111552
rect 19656 111492 19660 111548
rect 19660 111492 19716 111548
rect 19716 111492 19720 111548
rect 19656 111488 19720 111492
rect 19736 111548 19800 111552
rect 19736 111492 19740 111548
rect 19740 111492 19796 111548
rect 19796 111492 19800 111548
rect 19736 111488 19800 111492
rect 19816 111548 19880 111552
rect 19816 111492 19820 111548
rect 19820 111492 19876 111548
rect 19876 111492 19880 111548
rect 19816 111488 19880 111492
rect 4216 111004 4280 111008
rect 4216 110948 4220 111004
rect 4220 110948 4276 111004
rect 4276 110948 4280 111004
rect 4216 110944 4280 110948
rect 4296 111004 4360 111008
rect 4296 110948 4300 111004
rect 4300 110948 4356 111004
rect 4356 110948 4360 111004
rect 4296 110944 4360 110948
rect 4376 111004 4440 111008
rect 4376 110948 4380 111004
rect 4380 110948 4436 111004
rect 4436 110948 4440 111004
rect 4376 110944 4440 110948
rect 4456 111004 4520 111008
rect 4456 110948 4460 111004
rect 4460 110948 4516 111004
rect 4516 110948 4520 111004
rect 4456 110944 4520 110948
rect 34936 111004 35000 111008
rect 34936 110948 34940 111004
rect 34940 110948 34996 111004
rect 34996 110948 35000 111004
rect 34936 110944 35000 110948
rect 35016 111004 35080 111008
rect 35016 110948 35020 111004
rect 35020 110948 35076 111004
rect 35076 110948 35080 111004
rect 35016 110944 35080 110948
rect 35096 111004 35160 111008
rect 35096 110948 35100 111004
rect 35100 110948 35156 111004
rect 35156 110948 35160 111004
rect 35096 110944 35160 110948
rect 35176 111004 35240 111008
rect 35176 110948 35180 111004
rect 35180 110948 35236 111004
rect 35236 110948 35240 111004
rect 35176 110944 35240 110948
rect 19576 110460 19640 110464
rect 19576 110404 19580 110460
rect 19580 110404 19636 110460
rect 19636 110404 19640 110460
rect 19576 110400 19640 110404
rect 19656 110460 19720 110464
rect 19656 110404 19660 110460
rect 19660 110404 19716 110460
rect 19716 110404 19720 110460
rect 19656 110400 19720 110404
rect 19736 110460 19800 110464
rect 19736 110404 19740 110460
rect 19740 110404 19796 110460
rect 19796 110404 19800 110460
rect 19736 110400 19800 110404
rect 19816 110460 19880 110464
rect 19816 110404 19820 110460
rect 19820 110404 19876 110460
rect 19876 110404 19880 110460
rect 19816 110400 19880 110404
rect 4216 109916 4280 109920
rect 4216 109860 4220 109916
rect 4220 109860 4276 109916
rect 4276 109860 4280 109916
rect 4216 109856 4280 109860
rect 4296 109916 4360 109920
rect 4296 109860 4300 109916
rect 4300 109860 4356 109916
rect 4356 109860 4360 109916
rect 4296 109856 4360 109860
rect 4376 109916 4440 109920
rect 4376 109860 4380 109916
rect 4380 109860 4436 109916
rect 4436 109860 4440 109916
rect 4376 109856 4440 109860
rect 4456 109916 4520 109920
rect 4456 109860 4460 109916
rect 4460 109860 4516 109916
rect 4516 109860 4520 109916
rect 4456 109856 4520 109860
rect 34936 109916 35000 109920
rect 34936 109860 34940 109916
rect 34940 109860 34996 109916
rect 34996 109860 35000 109916
rect 34936 109856 35000 109860
rect 35016 109916 35080 109920
rect 35016 109860 35020 109916
rect 35020 109860 35076 109916
rect 35076 109860 35080 109916
rect 35016 109856 35080 109860
rect 35096 109916 35160 109920
rect 35096 109860 35100 109916
rect 35100 109860 35156 109916
rect 35156 109860 35160 109916
rect 35096 109856 35160 109860
rect 35176 109916 35240 109920
rect 35176 109860 35180 109916
rect 35180 109860 35236 109916
rect 35236 109860 35240 109916
rect 35176 109856 35240 109860
rect 19576 109372 19640 109376
rect 19576 109316 19580 109372
rect 19580 109316 19636 109372
rect 19636 109316 19640 109372
rect 19576 109312 19640 109316
rect 19656 109372 19720 109376
rect 19656 109316 19660 109372
rect 19660 109316 19716 109372
rect 19716 109316 19720 109372
rect 19656 109312 19720 109316
rect 19736 109372 19800 109376
rect 19736 109316 19740 109372
rect 19740 109316 19796 109372
rect 19796 109316 19800 109372
rect 19736 109312 19800 109316
rect 19816 109372 19880 109376
rect 19816 109316 19820 109372
rect 19820 109316 19876 109372
rect 19876 109316 19880 109372
rect 19816 109312 19880 109316
rect 4216 108828 4280 108832
rect 4216 108772 4220 108828
rect 4220 108772 4276 108828
rect 4276 108772 4280 108828
rect 4216 108768 4280 108772
rect 4296 108828 4360 108832
rect 4296 108772 4300 108828
rect 4300 108772 4356 108828
rect 4356 108772 4360 108828
rect 4296 108768 4360 108772
rect 4376 108828 4440 108832
rect 4376 108772 4380 108828
rect 4380 108772 4436 108828
rect 4436 108772 4440 108828
rect 4376 108768 4440 108772
rect 4456 108828 4520 108832
rect 4456 108772 4460 108828
rect 4460 108772 4516 108828
rect 4516 108772 4520 108828
rect 4456 108768 4520 108772
rect 34936 108828 35000 108832
rect 34936 108772 34940 108828
rect 34940 108772 34996 108828
rect 34996 108772 35000 108828
rect 34936 108768 35000 108772
rect 35016 108828 35080 108832
rect 35016 108772 35020 108828
rect 35020 108772 35076 108828
rect 35076 108772 35080 108828
rect 35016 108768 35080 108772
rect 35096 108828 35160 108832
rect 35096 108772 35100 108828
rect 35100 108772 35156 108828
rect 35156 108772 35160 108828
rect 35096 108768 35160 108772
rect 35176 108828 35240 108832
rect 35176 108772 35180 108828
rect 35180 108772 35236 108828
rect 35236 108772 35240 108828
rect 35176 108768 35240 108772
rect 19576 108284 19640 108288
rect 19576 108228 19580 108284
rect 19580 108228 19636 108284
rect 19636 108228 19640 108284
rect 19576 108224 19640 108228
rect 19656 108284 19720 108288
rect 19656 108228 19660 108284
rect 19660 108228 19716 108284
rect 19716 108228 19720 108284
rect 19656 108224 19720 108228
rect 19736 108284 19800 108288
rect 19736 108228 19740 108284
rect 19740 108228 19796 108284
rect 19796 108228 19800 108284
rect 19736 108224 19800 108228
rect 19816 108284 19880 108288
rect 19816 108228 19820 108284
rect 19820 108228 19876 108284
rect 19876 108228 19880 108284
rect 19816 108224 19880 108228
rect 4216 107740 4280 107744
rect 4216 107684 4220 107740
rect 4220 107684 4276 107740
rect 4276 107684 4280 107740
rect 4216 107680 4280 107684
rect 4296 107740 4360 107744
rect 4296 107684 4300 107740
rect 4300 107684 4356 107740
rect 4356 107684 4360 107740
rect 4296 107680 4360 107684
rect 4376 107740 4440 107744
rect 4376 107684 4380 107740
rect 4380 107684 4436 107740
rect 4436 107684 4440 107740
rect 4376 107680 4440 107684
rect 4456 107740 4520 107744
rect 4456 107684 4460 107740
rect 4460 107684 4516 107740
rect 4516 107684 4520 107740
rect 4456 107680 4520 107684
rect 34936 107740 35000 107744
rect 34936 107684 34940 107740
rect 34940 107684 34996 107740
rect 34996 107684 35000 107740
rect 34936 107680 35000 107684
rect 35016 107740 35080 107744
rect 35016 107684 35020 107740
rect 35020 107684 35076 107740
rect 35076 107684 35080 107740
rect 35016 107680 35080 107684
rect 35096 107740 35160 107744
rect 35096 107684 35100 107740
rect 35100 107684 35156 107740
rect 35156 107684 35160 107740
rect 35096 107680 35160 107684
rect 35176 107740 35240 107744
rect 35176 107684 35180 107740
rect 35180 107684 35236 107740
rect 35236 107684 35240 107740
rect 35176 107680 35240 107684
rect 19576 107196 19640 107200
rect 19576 107140 19580 107196
rect 19580 107140 19636 107196
rect 19636 107140 19640 107196
rect 19576 107136 19640 107140
rect 19656 107196 19720 107200
rect 19656 107140 19660 107196
rect 19660 107140 19716 107196
rect 19716 107140 19720 107196
rect 19656 107136 19720 107140
rect 19736 107196 19800 107200
rect 19736 107140 19740 107196
rect 19740 107140 19796 107196
rect 19796 107140 19800 107196
rect 19736 107136 19800 107140
rect 19816 107196 19880 107200
rect 19816 107140 19820 107196
rect 19820 107140 19876 107196
rect 19876 107140 19880 107196
rect 19816 107136 19880 107140
rect 4216 106652 4280 106656
rect 4216 106596 4220 106652
rect 4220 106596 4276 106652
rect 4276 106596 4280 106652
rect 4216 106592 4280 106596
rect 4296 106652 4360 106656
rect 4296 106596 4300 106652
rect 4300 106596 4356 106652
rect 4356 106596 4360 106652
rect 4296 106592 4360 106596
rect 4376 106652 4440 106656
rect 4376 106596 4380 106652
rect 4380 106596 4436 106652
rect 4436 106596 4440 106652
rect 4376 106592 4440 106596
rect 4456 106652 4520 106656
rect 4456 106596 4460 106652
rect 4460 106596 4516 106652
rect 4516 106596 4520 106652
rect 4456 106592 4520 106596
rect 34936 106652 35000 106656
rect 34936 106596 34940 106652
rect 34940 106596 34996 106652
rect 34996 106596 35000 106652
rect 34936 106592 35000 106596
rect 35016 106652 35080 106656
rect 35016 106596 35020 106652
rect 35020 106596 35076 106652
rect 35076 106596 35080 106652
rect 35016 106592 35080 106596
rect 35096 106652 35160 106656
rect 35096 106596 35100 106652
rect 35100 106596 35156 106652
rect 35156 106596 35160 106652
rect 35096 106592 35160 106596
rect 35176 106652 35240 106656
rect 35176 106596 35180 106652
rect 35180 106596 35236 106652
rect 35236 106596 35240 106652
rect 35176 106592 35240 106596
rect 19576 106108 19640 106112
rect 19576 106052 19580 106108
rect 19580 106052 19636 106108
rect 19636 106052 19640 106108
rect 19576 106048 19640 106052
rect 19656 106108 19720 106112
rect 19656 106052 19660 106108
rect 19660 106052 19716 106108
rect 19716 106052 19720 106108
rect 19656 106048 19720 106052
rect 19736 106108 19800 106112
rect 19736 106052 19740 106108
rect 19740 106052 19796 106108
rect 19796 106052 19800 106108
rect 19736 106048 19800 106052
rect 19816 106108 19880 106112
rect 19816 106052 19820 106108
rect 19820 106052 19876 106108
rect 19876 106052 19880 106108
rect 19816 106048 19880 106052
rect 4216 105564 4280 105568
rect 4216 105508 4220 105564
rect 4220 105508 4276 105564
rect 4276 105508 4280 105564
rect 4216 105504 4280 105508
rect 4296 105564 4360 105568
rect 4296 105508 4300 105564
rect 4300 105508 4356 105564
rect 4356 105508 4360 105564
rect 4296 105504 4360 105508
rect 4376 105564 4440 105568
rect 4376 105508 4380 105564
rect 4380 105508 4436 105564
rect 4436 105508 4440 105564
rect 4376 105504 4440 105508
rect 4456 105564 4520 105568
rect 4456 105508 4460 105564
rect 4460 105508 4516 105564
rect 4516 105508 4520 105564
rect 4456 105504 4520 105508
rect 34936 105564 35000 105568
rect 34936 105508 34940 105564
rect 34940 105508 34996 105564
rect 34996 105508 35000 105564
rect 34936 105504 35000 105508
rect 35016 105564 35080 105568
rect 35016 105508 35020 105564
rect 35020 105508 35076 105564
rect 35076 105508 35080 105564
rect 35016 105504 35080 105508
rect 35096 105564 35160 105568
rect 35096 105508 35100 105564
rect 35100 105508 35156 105564
rect 35156 105508 35160 105564
rect 35096 105504 35160 105508
rect 35176 105564 35240 105568
rect 35176 105508 35180 105564
rect 35180 105508 35236 105564
rect 35236 105508 35240 105564
rect 35176 105504 35240 105508
rect 19576 105020 19640 105024
rect 19576 104964 19580 105020
rect 19580 104964 19636 105020
rect 19636 104964 19640 105020
rect 19576 104960 19640 104964
rect 19656 105020 19720 105024
rect 19656 104964 19660 105020
rect 19660 104964 19716 105020
rect 19716 104964 19720 105020
rect 19656 104960 19720 104964
rect 19736 105020 19800 105024
rect 19736 104964 19740 105020
rect 19740 104964 19796 105020
rect 19796 104964 19800 105020
rect 19736 104960 19800 104964
rect 19816 105020 19880 105024
rect 19816 104964 19820 105020
rect 19820 104964 19876 105020
rect 19876 104964 19880 105020
rect 19816 104960 19880 104964
rect 4216 104476 4280 104480
rect 4216 104420 4220 104476
rect 4220 104420 4276 104476
rect 4276 104420 4280 104476
rect 4216 104416 4280 104420
rect 4296 104476 4360 104480
rect 4296 104420 4300 104476
rect 4300 104420 4356 104476
rect 4356 104420 4360 104476
rect 4296 104416 4360 104420
rect 4376 104476 4440 104480
rect 4376 104420 4380 104476
rect 4380 104420 4436 104476
rect 4436 104420 4440 104476
rect 4376 104416 4440 104420
rect 4456 104476 4520 104480
rect 4456 104420 4460 104476
rect 4460 104420 4516 104476
rect 4516 104420 4520 104476
rect 4456 104416 4520 104420
rect 34936 104476 35000 104480
rect 34936 104420 34940 104476
rect 34940 104420 34996 104476
rect 34996 104420 35000 104476
rect 34936 104416 35000 104420
rect 35016 104476 35080 104480
rect 35016 104420 35020 104476
rect 35020 104420 35076 104476
rect 35076 104420 35080 104476
rect 35016 104416 35080 104420
rect 35096 104476 35160 104480
rect 35096 104420 35100 104476
rect 35100 104420 35156 104476
rect 35156 104420 35160 104476
rect 35096 104416 35160 104420
rect 35176 104476 35240 104480
rect 35176 104420 35180 104476
rect 35180 104420 35236 104476
rect 35236 104420 35240 104476
rect 35176 104416 35240 104420
rect 19576 103932 19640 103936
rect 19576 103876 19580 103932
rect 19580 103876 19636 103932
rect 19636 103876 19640 103932
rect 19576 103872 19640 103876
rect 19656 103932 19720 103936
rect 19656 103876 19660 103932
rect 19660 103876 19716 103932
rect 19716 103876 19720 103932
rect 19656 103872 19720 103876
rect 19736 103932 19800 103936
rect 19736 103876 19740 103932
rect 19740 103876 19796 103932
rect 19796 103876 19800 103932
rect 19736 103872 19800 103876
rect 19816 103932 19880 103936
rect 19816 103876 19820 103932
rect 19820 103876 19876 103932
rect 19876 103876 19880 103932
rect 19816 103872 19880 103876
rect 4216 103388 4280 103392
rect 4216 103332 4220 103388
rect 4220 103332 4276 103388
rect 4276 103332 4280 103388
rect 4216 103328 4280 103332
rect 4296 103388 4360 103392
rect 4296 103332 4300 103388
rect 4300 103332 4356 103388
rect 4356 103332 4360 103388
rect 4296 103328 4360 103332
rect 4376 103388 4440 103392
rect 4376 103332 4380 103388
rect 4380 103332 4436 103388
rect 4436 103332 4440 103388
rect 4376 103328 4440 103332
rect 4456 103388 4520 103392
rect 4456 103332 4460 103388
rect 4460 103332 4516 103388
rect 4516 103332 4520 103388
rect 4456 103328 4520 103332
rect 34936 103388 35000 103392
rect 34936 103332 34940 103388
rect 34940 103332 34996 103388
rect 34996 103332 35000 103388
rect 34936 103328 35000 103332
rect 35016 103388 35080 103392
rect 35016 103332 35020 103388
rect 35020 103332 35076 103388
rect 35076 103332 35080 103388
rect 35016 103328 35080 103332
rect 35096 103388 35160 103392
rect 35096 103332 35100 103388
rect 35100 103332 35156 103388
rect 35156 103332 35160 103388
rect 35096 103328 35160 103332
rect 35176 103388 35240 103392
rect 35176 103332 35180 103388
rect 35180 103332 35236 103388
rect 35236 103332 35240 103388
rect 35176 103328 35240 103332
rect 19576 102844 19640 102848
rect 19576 102788 19580 102844
rect 19580 102788 19636 102844
rect 19636 102788 19640 102844
rect 19576 102784 19640 102788
rect 19656 102844 19720 102848
rect 19656 102788 19660 102844
rect 19660 102788 19716 102844
rect 19716 102788 19720 102844
rect 19656 102784 19720 102788
rect 19736 102844 19800 102848
rect 19736 102788 19740 102844
rect 19740 102788 19796 102844
rect 19796 102788 19800 102844
rect 19736 102784 19800 102788
rect 19816 102844 19880 102848
rect 19816 102788 19820 102844
rect 19820 102788 19876 102844
rect 19876 102788 19880 102844
rect 19816 102784 19880 102788
rect 4216 102300 4280 102304
rect 4216 102244 4220 102300
rect 4220 102244 4276 102300
rect 4276 102244 4280 102300
rect 4216 102240 4280 102244
rect 4296 102300 4360 102304
rect 4296 102244 4300 102300
rect 4300 102244 4356 102300
rect 4356 102244 4360 102300
rect 4296 102240 4360 102244
rect 4376 102300 4440 102304
rect 4376 102244 4380 102300
rect 4380 102244 4436 102300
rect 4436 102244 4440 102300
rect 4376 102240 4440 102244
rect 4456 102300 4520 102304
rect 4456 102244 4460 102300
rect 4460 102244 4516 102300
rect 4516 102244 4520 102300
rect 4456 102240 4520 102244
rect 34936 102300 35000 102304
rect 34936 102244 34940 102300
rect 34940 102244 34996 102300
rect 34996 102244 35000 102300
rect 34936 102240 35000 102244
rect 35016 102300 35080 102304
rect 35016 102244 35020 102300
rect 35020 102244 35076 102300
rect 35076 102244 35080 102300
rect 35016 102240 35080 102244
rect 35096 102300 35160 102304
rect 35096 102244 35100 102300
rect 35100 102244 35156 102300
rect 35156 102244 35160 102300
rect 35096 102240 35160 102244
rect 35176 102300 35240 102304
rect 35176 102244 35180 102300
rect 35180 102244 35236 102300
rect 35236 102244 35240 102300
rect 35176 102240 35240 102244
rect 19576 101756 19640 101760
rect 19576 101700 19580 101756
rect 19580 101700 19636 101756
rect 19636 101700 19640 101756
rect 19576 101696 19640 101700
rect 19656 101756 19720 101760
rect 19656 101700 19660 101756
rect 19660 101700 19716 101756
rect 19716 101700 19720 101756
rect 19656 101696 19720 101700
rect 19736 101756 19800 101760
rect 19736 101700 19740 101756
rect 19740 101700 19796 101756
rect 19796 101700 19800 101756
rect 19736 101696 19800 101700
rect 19816 101756 19880 101760
rect 19816 101700 19820 101756
rect 19820 101700 19876 101756
rect 19876 101700 19880 101756
rect 19816 101696 19880 101700
rect 4216 101212 4280 101216
rect 4216 101156 4220 101212
rect 4220 101156 4276 101212
rect 4276 101156 4280 101212
rect 4216 101152 4280 101156
rect 4296 101212 4360 101216
rect 4296 101156 4300 101212
rect 4300 101156 4356 101212
rect 4356 101156 4360 101212
rect 4296 101152 4360 101156
rect 4376 101212 4440 101216
rect 4376 101156 4380 101212
rect 4380 101156 4436 101212
rect 4436 101156 4440 101212
rect 4376 101152 4440 101156
rect 4456 101212 4520 101216
rect 4456 101156 4460 101212
rect 4460 101156 4516 101212
rect 4516 101156 4520 101212
rect 4456 101152 4520 101156
rect 34936 101212 35000 101216
rect 34936 101156 34940 101212
rect 34940 101156 34996 101212
rect 34996 101156 35000 101212
rect 34936 101152 35000 101156
rect 35016 101212 35080 101216
rect 35016 101156 35020 101212
rect 35020 101156 35076 101212
rect 35076 101156 35080 101212
rect 35016 101152 35080 101156
rect 35096 101212 35160 101216
rect 35096 101156 35100 101212
rect 35100 101156 35156 101212
rect 35156 101156 35160 101212
rect 35096 101152 35160 101156
rect 35176 101212 35240 101216
rect 35176 101156 35180 101212
rect 35180 101156 35236 101212
rect 35236 101156 35240 101212
rect 35176 101152 35240 101156
rect 19576 100668 19640 100672
rect 19576 100612 19580 100668
rect 19580 100612 19636 100668
rect 19636 100612 19640 100668
rect 19576 100608 19640 100612
rect 19656 100668 19720 100672
rect 19656 100612 19660 100668
rect 19660 100612 19716 100668
rect 19716 100612 19720 100668
rect 19656 100608 19720 100612
rect 19736 100668 19800 100672
rect 19736 100612 19740 100668
rect 19740 100612 19796 100668
rect 19796 100612 19800 100668
rect 19736 100608 19800 100612
rect 19816 100668 19880 100672
rect 19816 100612 19820 100668
rect 19820 100612 19876 100668
rect 19876 100612 19880 100668
rect 19816 100608 19880 100612
rect 4216 100124 4280 100128
rect 4216 100068 4220 100124
rect 4220 100068 4276 100124
rect 4276 100068 4280 100124
rect 4216 100064 4280 100068
rect 4296 100124 4360 100128
rect 4296 100068 4300 100124
rect 4300 100068 4356 100124
rect 4356 100068 4360 100124
rect 4296 100064 4360 100068
rect 4376 100124 4440 100128
rect 4376 100068 4380 100124
rect 4380 100068 4436 100124
rect 4436 100068 4440 100124
rect 4376 100064 4440 100068
rect 4456 100124 4520 100128
rect 4456 100068 4460 100124
rect 4460 100068 4516 100124
rect 4516 100068 4520 100124
rect 4456 100064 4520 100068
rect 34936 100124 35000 100128
rect 34936 100068 34940 100124
rect 34940 100068 34996 100124
rect 34996 100068 35000 100124
rect 34936 100064 35000 100068
rect 35016 100124 35080 100128
rect 35016 100068 35020 100124
rect 35020 100068 35076 100124
rect 35076 100068 35080 100124
rect 35016 100064 35080 100068
rect 35096 100124 35160 100128
rect 35096 100068 35100 100124
rect 35100 100068 35156 100124
rect 35156 100068 35160 100124
rect 35096 100064 35160 100068
rect 35176 100124 35240 100128
rect 35176 100068 35180 100124
rect 35180 100068 35236 100124
rect 35236 100068 35240 100124
rect 35176 100064 35240 100068
rect 19576 99580 19640 99584
rect 19576 99524 19580 99580
rect 19580 99524 19636 99580
rect 19636 99524 19640 99580
rect 19576 99520 19640 99524
rect 19656 99580 19720 99584
rect 19656 99524 19660 99580
rect 19660 99524 19716 99580
rect 19716 99524 19720 99580
rect 19656 99520 19720 99524
rect 19736 99580 19800 99584
rect 19736 99524 19740 99580
rect 19740 99524 19796 99580
rect 19796 99524 19800 99580
rect 19736 99520 19800 99524
rect 19816 99580 19880 99584
rect 19816 99524 19820 99580
rect 19820 99524 19876 99580
rect 19876 99524 19880 99580
rect 19816 99520 19880 99524
rect 4216 99036 4280 99040
rect 4216 98980 4220 99036
rect 4220 98980 4276 99036
rect 4276 98980 4280 99036
rect 4216 98976 4280 98980
rect 4296 99036 4360 99040
rect 4296 98980 4300 99036
rect 4300 98980 4356 99036
rect 4356 98980 4360 99036
rect 4296 98976 4360 98980
rect 4376 99036 4440 99040
rect 4376 98980 4380 99036
rect 4380 98980 4436 99036
rect 4436 98980 4440 99036
rect 4376 98976 4440 98980
rect 4456 99036 4520 99040
rect 4456 98980 4460 99036
rect 4460 98980 4516 99036
rect 4516 98980 4520 99036
rect 4456 98976 4520 98980
rect 34936 99036 35000 99040
rect 34936 98980 34940 99036
rect 34940 98980 34996 99036
rect 34996 98980 35000 99036
rect 34936 98976 35000 98980
rect 35016 99036 35080 99040
rect 35016 98980 35020 99036
rect 35020 98980 35076 99036
rect 35076 98980 35080 99036
rect 35016 98976 35080 98980
rect 35096 99036 35160 99040
rect 35096 98980 35100 99036
rect 35100 98980 35156 99036
rect 35156 98980 35160 99036
rect 35096 98976 35160 98980
rect 35176 99036 35240 99040
rect 35176 98980 35180 99036
rect 35180 98980 35236 99036
rect 35236 98980 35240 99036
rect 35176 98976 35240 98980
rect 19576 98492 19640 98496
rect 19576 98436 19580 98492
rect 19580 98436 19636 98492
rect 19636 98436 19640 98492
rect 19576 98432 19640 98436
rect 19656 98492 19720 98496
rect 19656 98436 19660 98492
rect 19660 98436 19716 98492
rect 19716 98436 19720 98492
rect 19656 98432 19720 98436
rect 19736 98492 19800 98496
rect 19736 98436 19740 98492
rect 19740 98436 19796 98492
rect 19796 98436 19800 98492
rect 19736 98432 19800 98436
rect 19816 98492 19880 98496
rect 19816 98436 19820 98492
rect 19820 98436 19876 98492
rect 19876 98436 19880 98492
rect 19816 98432 19880 98436
rect 4216 97948 4280 97952
rect 4216 97892 4220 97948
rect 4220 97892 4276 97948
rect 4276 97892 4280 97948
rect 4216 97888 4280 97892
rect 4296 97948 4360 97952
rect 4296 97892 4300 97948
rect 4300 97892 4356 97948
rect 4356 97892 4360 97948
rect 4296 97888 4360 97892
rect 4376 97948 4440 97952
rect 4376 97892 4380 97948
rect 4380 97892 4436 97948
rect 4436 97892 4440 97948
rect 4376 97888 4440 97892
rect 4456 97948 4520 97952
rect 4456 97892 4460 97948
rect 4460 97892 4516 97948
rect 4516 97892 4520 97948
rect 4456 97888 4520 97892
rect 34936 97948 35000 97952
rect 34936 97892 34940 97948
rect 34940 97892 34996 97948
rect 34996 97892 35000 97948
rect 34936 97888 35000 97892
rect 35016 97948 35080 97952
rect 35016 97892 35020 97948
rect 35020 97892 35076 97948
rect 35076 97892 35080 97948
rect 35016 97888 35080 97892
rect 35096 97948 35160 97952
rect 35096 97892 35100 97948
rect 35100 97892 35156 97948
rect 35156 97892 35160 97948
rect 35096 97888 35160 97892
rect 35176 97948 35240 97952
rect 35176 97892 35180 97948
rect 35180 97892 35236 97948
rect 35236 97892 35240 97948
rect 35176 97888 35240 97892
rect 19576 97404 19640 97408
rect 19576 97348 19580 97404
rect 19580 97348 19636 97404
rect 19636 97348 19640 97404
rect 19576 97344 19640 97348
rect 19656 97404 19720 97408
rect 19656 97348 19660 97404
rect 19660 97348 19716 97404
rect 19716 97348 19720 97404
rect 19656 97344 19720 97348
rect 19736 97404 19800 97408
rect 19736 97348 19740 97404
rect 19740 97348 19796 97404
rect 19796 97348 19800 97404
rect 19736 97344 19800 97348
rect 19816 97404 19880 97408
rect 19816 97348 19820 97404
rect 19820 97348 19876 97404
rect 19876 97348 19880 97404
rect 19816 97344 19880 97348
rect 4216 96860 4280 96864
rect 4216 96804 4220 96860
rect 4220 96804 4276 96860
rect 4276 96804 4280 96860
rect 4216 96800 4280 96804
rect 4296 96860 4360 96864
rect 4296 96804 4300 96860
rect 4300 96804 4356 96860
rect 4356 96804 4360 96860
rect 4296 96800 4360 96804
rect 4376 96860 4440 96864
rect 4376 96804 4380 96860
rect 4380 96804 4436 96860
rect 4436 96804 4440 96860
rect 4376 96800 4440 96804
rect 4456 96860 4520 96864
rect 4456 96804 4460 96860
rect 4460 96804 4516 96860
rect 4516 96804 4520 96860
rect 4456 96800 4520 96804
rect 34936 96860 35000 96864
rect 34936 96804 34940 96860
rect 34940 96804 34996 96860
rect 34996 96804 35000 96860
rect 34936 96800 35000 96804
rect 35016 96860 35080 96864
rect 35016 96804 35020 96860
rect 35020 96804 35076 96860
rect 35076 96804 35080 96860
rect 35016 96800 35080 96804
rect 35096 96860 35160 96864
rect 35096 96804 35100 96860
rect 35100 96804 35156 96860
rect 35156 96804 35160 96860
rect 35096 96800 35160 96804
rect 35176 96860 35240 96864
rect 35176 96804 35180 96860
rect 35180 96804 35236 96860
rect 35236 96804 35240 96860
rect 35176 96800 35240 96804
rect 19576 96316 19640 96320
rect 19576 96260 19580 96316
rect 19580 96260 19636 96316
rect 19636 96260 19640 96316
rect 19576 96256 19640 96260
rect 19656 96316 19720 96320
rect 19656 96260 19660 96316
rect 19660 96260 19716 96316
rect 19716 96260 19720 96316
rect 19656 96256 19720 96260
rect 19736 96316 19800 96320
rect 19736 96260 19740 96316
rect 19740 96260 19796 96316
rect 19796 96260 19800 96316
rect 19736 96256 19800 96260
rect 19816 96316 19880 96320
rect 19816 96260 19820 96316
rect 19820 96260 19876 96316
rect 19876 96260 19880 96316
rect 19816 96256 19880 96260
rect 4216 95772 4280 95776
rect 4216 95716 4220 95772
rect 4220 95716 4276 95772
rect 4276 95716 4280 95772
rect 4216 95712 4280 95716
rect 4296 95772 4360 95776
rect 4296 95716 4300 95772
rect 4300 95716 4356 95772
rect 4356 95716 4360 95772
rect 4296 95712 4360 95716
rect 4376 95772 4440 95776
rect 4376 95716 4380 95772
rect 4380 95716 4436 95772
rect 4436 95716 4440 95772
rect 4376 95712 4440 95716
rect 4456 95772 4520 95776
rect 4456 95716 4460 95772
rect 4460 95716 4516 95772
rect 4516 95716 4520 95772
rect 4456 95712 4520 95716
rect 34936 95772 35000 95776
rect 34936 95716 34940 95772
rect 34940 95716 34996 95772
rect 34996 95716 35000 95772
rect 34936 95712 35000 95716
rect 35016 95772 35080 95776
rect 35016 95716 35020 95772
rect 35020 95716 35076 95772
rect 35076 95716 35080 95772
rect 35016 95712 35080 95716
rect 35096 95772 35160 95776
rect 35096 95716 35100 95772
rect 35100 95716 35156 95772
rect 35156 95716 35160 95772
rect 35096 95712 35160 95716
rect 35176 95772 35240 95776
rect 35176 95716 35180 95772
rect 35180 95716 35236 95772
rect 35236 95716 35240 95772
rect 35176 95712 35240 95716
rect 19576 95228 19640 95232
rect 19576 95172 19580 95228
rect 19580 95172 19636 95228
rect 19636 95172 19640 95228
rect 19576 95168 19640 95172
rect 19656 95228 19720 95232
rect 19656 95172 19660 95228
rect 19660 95172 19716 95228
rect 19716 95172 19720 95228
rect 19656 95168 19720 95172
rect 19736 95228 19800 95232
rect 19736 95172 19740 95228
rect 19740 95172 19796 95228
rect 19796 95172 19800 95228
rect 19736 95168 19800 95172
rect 19816 95228 19880 95232
rect 19816 95172 19820 95228
rect 19820 95172 19876 95228
rect 19876 95172 19880 95228
rect 19816 95168 19880 95172
rect 4216 94684 4280 94688
rect 4216 94628 4220 94684
rect 4220 94628 4276 94684
rect 4276 94628 4280 94684
rect 4216 94624 4280 94628
rect 4296 94684 4360 94688
rect 4296 94628 4300 94684
rect 4300 94628 4356 94684
rect 4356 94628 4360 94684
rect 4296 94624 4360 94628
rect 4376 94684 4440 94688
rect 4376 94628 4380 94684
rect 4380 94628 4436 94684
rect 4436 94628 4440 94684
rect 4376 94624 4440 94628
rect 4456 94684 4520 94688
rect 4456 94628 4460 94684
rect 4460 94628 4516 94684
rect 4516 94628 4520 94684
rect 4456 94624 4520 94628
rect 34936 94684 35000 94688
rect 34936 94628 34940 94684
rect 34940 94628 34996 94684
rect 34996 94628 35000 94684
rect 34936 94624 35000 94628
rect 35016 94684 35080 94688
rect 35016 94628 35020 94684
rect 35020 94628 35076 94684
rect 35076 94628 35080 94684
rect 35016 94624 35080 94628
rect 35096 94684 35160 94688
rect 35096 94628 35100 94684
rect 35100 94628 35156 94684
rect 35156 94628 35160 94684
rect 35096 94624 35160 94628
rect 35176 94684 35240 94688
rect 35176 94628 35180 94684
rect 35180 94628 35236 94684
rect 35236 94628 35240 94684
rect 35176 94624 35240 94628
rect 19576 94140 19640 94144
rect 19576 94084 19580 94140
rect 19580 94084 19636 94140
rect 19636 94084 19640 94140
rect 19576 94080 19640 94084
rect 19656 94140 19720 94144
rect 19656 94084 19660 94140
rect 19660 94084 19716 94140
rect 19716 94084 19720 94140
rect 19656 94080 19720 94084
rect 19736 94140 19800 94144
rect 19736 94084 19740 94140
rect 19740 94084 19796 94140
rect 19796 94084 19800 94140
rect 19736 94080 19800 94084
rect 19816 94140 19880 94144
rect 19816 94084 19820 94140
rect 19820 94084 19876 94140
rect 19876 94084 19880 94140
rect 19816 94080 19880 94084
rect 4216 93596 4280 93600
rect 4216 93540 4220 93596
rect 4220 93540 4276 93596
rect 4276 93540 4280 93596
rect 4216 93536 4280 93540
rect 4296 93596 4360 93600
rect 4296 93540 4300 93596
rect 4300 93540 4356 93596
rect 4356 93540 4360 93596
rect 4296 93536 4360 93540
rect 4376 93596 4440 93600
rect 4376 93540 4380 93596
rect 4380 93540 4436 93596
rect 4436 93540 4440 93596
rect 4376 93536 4440 93540
rect 4456 93596 4520 93600
rect 4456 93540 4460 93596
rect 4460 93540 4516 93596
rect 4516 93540 4520 93596
rect 4456 93536 4520 93540
rect 34936 93596 35000 93600
rect 34936 93540 34940 93596
rect 34940 93540 34996 93596
rect 34996 93540 35000 93596
rect 34936 93536 35000 93540
rect 35016 93596 35080 93600
rect 35016 93540 35020 93596
rect 35020 93540 35076 93596
rect 35076 93540 35080 93596
rect 35016 93536 35080 93540
rect 35096 93596 35160 93600
rect 35096 93540 35100 93596
rect 35100 93540 35156 93596
rect 35156 93540 35160 93596
rect 35096 93536 35160 93540
rect 35176 93596 35240 93600
rect 35176 93540 35180 93596
rect 35180 93540 35236 93596
rect 35236 93540 35240 93596
rect 35176 93536 35240 93540
rect 19576 93052 19640 93056
rect 19576 92996 19580 93052
rect 19580 92996 19636 93052
rect 19636 92996 19640 93052
rect 19576 92992 19640 92996
rect 19656 93052 19720 93056
rect 19656 92996 19660 93052
rect 19660 92996 19716 93052
rect 19716 92996 19720 93052
rect 19656 92992 19720 92996
rect 19736 93052 19800 93056
rect 19736 92996 19740 93052
rect 19740 92996 19796 93052
rect 19796 92996 19800 93052
rect 19736 92992 19800 92996
rect 19816 93052 19880 93056
rect 19816 92996 19820 93052
rect 19820 92996 19876 93052
rect 19876 92996 19880 93052
rect 19816 92992 19880 92996
rect 4216 92508 4280 92512
rect 4216 92452 4220 92508
rect 4220 92452 4276 92508
rect 4276 92452 4280 92508
rect 4216 92448 4280 92452
rect 4296 92508 4360 92512
rect 4296 92452 4300 92508
rect 4300 92452 4356 92508
rect 4356 92452 4360 92508
rect 4296 92448 4360 92452
rect 4376 92508 4440 92512
rect 4376 92452 4380 92508
rect 4380 92452 4436 92508
rect 4436 92452 4440 92508
rect 4376 92448 4440 92452
rect 4456 92508 4520 92512
rect 4456 92452 4460 92508
rect 4460 92452 4516 92508
rect 4516 92452 4520 92508
rect 4456 92448 4520 92452
rect 34936 92508 35000 92512
rect 34936 92452 34940 92508
rect 34940 92452 34996 92508
rect 34996 92452 35000 92508
rect 34936 92448 35000 92452
rect 35016 92508 35080 92512
rect 35016 92452 35020 92508
rect 35020 92452 35076 92508
rect 35076 92452 35080 92508
rect 35016 92448 35080 92452
rect 35096 92508 35160 92512
rect 35096 92452 35100 92508
rect 35100 92452 35156 92508
rect 35156 92452 35160 92508
rect 35096 92448 35160 92452
rect 35176 92508 35240 92512
rect 35176 92452 35180 92508
rect 35180 92452 35236 92508
rect 35236 92452 35240 92508
rect 35176 92448 35240 92452
rect 19576 91964 19640 91968
rect 19576 91908 19580 91964
rect 19580 91908 19636 91964
rect 19636 91908 19640 91964
rect 19576 91904 19640 91908
rect 19656 91964 19720 91968
rect 19656 91908 19660 91964
rect 19660 91908 19716 91964
rect 19716 91908 19720 91964
rect 19656 91904 19720 91908
rect 19736 91964 19800 91968
rect 19736 91908 19740 91964
rect 19740 91908 19796 91964
rect 19796 91908 19800 91964
rect 19736 91904 19800 91908
rect 19816 91964 19880 91968
rect 19816 91908 19820 91964
rect 19820 91908 19876 91964
rect 19876 91908 19880 91964
rect 19816 91904 19880 91908
rect 4216 91420 4280 91424
rect 4216 91364 4220 91420
rect 4220 91364 4276 91420
rect 4276 91364 4280 91420
rect 4216 91360 4280 91364
rect 4296 91420 4360 91424
rect 4296 91364 4300 91420
rect 4300 91364 4356 91420
rect 4356 91364 4360 91420
rect 4296 91360 4360 91364
rect 4376 91420 4440 91424
rect 4376 91364 4380 91420
rect 4380 91364 4436 91420
rect 4436 91364 4440 91420
rect 4376 91360 4440 91364
rect 4456 91420 4520 91424
rect 4456 91364 4460 91420
rect 4460 91364 4516 91420
rect 4516 91364 4520 91420
rect 4456 91360 4520 91364
rect 34936 91420 35000 91424
rect 34936 91364 34940 91420
rect 34940 91364 34996 91420
rect 34996 91364 35000 91420
rect 34936 91360 35000 91364
rect 35016 91420 35080 91424
rect 35016 91364 35020 91420
rect 35020 91364 35076 91420
rect 35076 91364 35080 91420
rect 35016 91360 35080 91364
rect 35096 91420 35160 91424
rect 35096 91364 35100 91420
rect 35100 91364 35156 91420
rect 35156 91364 35160 91420
rect 35096 91360 35160 91364
rect 35176 91420 35240 91424
rect 35176 91364 35180 91420
rect 35180 91364 35236 91420
rect 35236 91364 35240 91420
rect 35176 91360 35240 91364
rect 19576 90876 19640 90880
rect 19576 90820 19580 90876
rect 19580 90820 19636 90876
rect 19636 90820 19640 90876
rect 19576 90816 19640 90820
rect 19656 90876 19720 90880
rect 19656 90820 19660 90876
rect 19660 90820 19716 90876
rect 19716 90820 19720 90876
rect 19656 90816 19720 90820
rect 19736 90876 19800 90880
rect 19736 90820 19740 90876
rect 19740 90820 19796 90876
rect 19796 90820 19800 90876
rect 19736 90816 19800 90820
rect 19816 90876 19880 90880
rect 19816 90820 19820 90876
rect 19820 90820 19876 90876
rect 19876 90820 19880 90876
rect 19816 90816 19880 90820
rect 4216 90332 4280 90336
rect 4216 90276 4220 90332
rect 4220 90276 4276 90332
rect 4276 90276 4280 90332
rect 4216 90272 4280 90276
rect 4296 90332 4360 90336
rect 4296 90276 4300 90332
rect 4300 90276 4356 90332
rect 4356 90276 4360 90332
rect 4296 90272 4360 90276
rect 4376 90332 4440 90336
rect 4376 90276 4380 90332
rect 4380 90276 4436 90332
rect 4436 90276 4440 90332
rect 4376 90272 4440 90276
rect 4456 90332 4520 90336
rect 4456 90276 4460 90332
rect 4460 90276 4516 90332
rect 4516 90276 4520 90332
rect 4456 90272 4520 90276
rect 34936 90332 35000 90336
rect 34936 90276 34940 90332
rect 34940 90276 34996 90332
rect 34996 90276 35000 90332
rect 34936 90272 35000 90276
rect 35016 90332 35080 90336
rect 35016 90276 35020 90332
rect 35020 90276 35076 90332
rect 35076 90276 35080 90332
rect 35016 90272 35080 90276
rect 35096 90332 35160 90336
rect 35096 90276 35100 90332
rect 35100 90276 35156 90332
rect 35156 90276 35160 90332
rect 35096 90272 35160 90276
rect 35176 90332 35240 90336
rect 35176 90276 35180 90332
rect 35180 90276 35236 90332
rect 35236 90276 35240 90332
rect 35176 90272 35240 90276
rect 19576 89788 19640 89792
rect 19576 89732 19580 89788
rect 19580 89732 19636 89788
rect 19636 89732 19640 89788
rect 19576 89728 19640 89732
rect 19656 89788 19720 89792
rect 19656 89732 19660 89788
rect 19660 89732 19716 89788
rect 19716 89732 19720 89788
rect 19656 89728 19720 89732
rect 19736 89788 19800 89792
rect 19736 89732 19740 89788
rect 19740 89732 19796 89788
rect 19796 89732 19800 89788
rect 19736 89728 19800 89732
rect 19816 89788 19880 89792
rect 19816 89732 19820 89788
rect 19820 89732 19876 89788
rect 19876 89732 19880 89788
rect 19816 89728 19880 89732
rect 4216 89244 4280 89248
rect 4216 89188 4220 89244
rect 4220 89188 4276 89244
rect 4276 89188 4280 89244
rect 4216 89184 4280 89188
rect 4296 89244 4360 89248
rect 4296 89188 4300 89244
rect 4300 89188 4356 89244
rect 4356 89188 4360 89244
rect 4296 89184 4360 89188
rect 4376 89244 4440 89248
rect 4376 89188 4380 89244
rect 4380 89188 4436 89244
rect 4436 89188 4440 89244
rect 4376 89184 4440 89188
rect 4456 89244 4520 89248
rect 4456 89188 4460 89244
rect 4460 89188 4516 89244
rect 4516 89188 4520 89244
rect 4456 89184 4520 89188
rect 34936 89244 35000 89248
rect 34936 89188 34940 89244
rect 34940 89188 34996 89244
rect 34996 89188 35000 89244
rect 34936 89184 35000 89188
rect 35016 89244 35080 89248
rect 35016 89188 35020 89244
rect 35020 89188 35076 89244
rect 35076 89188 35080 89244
rect 35016 89184 35080 89188
rect 35096 89244 35160 89248
rect 35096 89188 35100 89244
rect 35100 89188 35156 89244
rect 35156 89188 35160 89244
rect 35096 89184 35160 89188
rect 35176 89244 35240 89248
rect 35176 89188 35180 89244
rect 35180 89188 35236 89244
rect 35236 89188 35240 89244
rect 35176 89184 35240 89188
rect 19576 88700 19640 88704
rect 19576 88644 19580 88700
rect 19580 88644 19636 88700
rect 19636 88644 19640 88700
rect 19576 88640 19640 88644
rect 19656 88700 19720 88704
rect 19656 88644 19660 88700
rect 19660 88644 19716 88700
rect 19716 88644 19720 88700
rect 19656 88640 19720 88644
rect 19736 88700 19800 88704
rect 19736 88644 19740 88700
rect 19740 88644 19796 88700
rect 19796 88644 19800 88700
rect 19736 88640 19800 88644
rect 19816 88700 19880 88704
rect 19816 88644 19820 88700
rect 19820 88644 19876 88700
rect 19876 88644 19880 88700
rect 19816 88640 19880 88644
rect 4216 88156 4280 88160
rect 4216 88100 4220 88156
rect 4220 88100 4276 88156
rect 4276 88100 4280 88156
rect 4216 88096 4280 88100
rect 4296 88156 4360 88160
rect 4296 88100 4300 88156
rect 4300 88100 4356 88156
rect 4356 88100 4360 88156
rect 4296 88096 4360 88100
rect 4376 88156 4440 88160
rect 4376 88100 4380 88156
rect 4380 88100 4436 88156
rect 4436 88100 4440 88156
rect 4376 88096 4440 88100
rect 4456 88156 4520 88160
rect 4456 88100 4460 88156
rect 4460 88100 4516 88156
rect 4516 88100 4520 88156
rect 4456 88096 4520 88100
rect 34936 88156 35000 88160
rect 34936 88100 34940 88156
rect 34940 88100 34996 88156
rect 34996 88100 35000 88156
rect 34936 88096 35000 88100
rect 35016 88156 35080 88160
rect 35016 88100 35020 88156
rect 35020 88100 35076 88156
rect 35076 88100 35080 88156
rect 35016 88096 35080 88100
rect 35096 88156 35160 88160
rect 35096 88100 35100 88156
rect 35100 88100 35156 88156
rect 35156 88100 35160 88156
rect 35096 88096 35160 88100
rect 35176 88156 35240 88160
rect 35176 88100 35180 88156
rect 35180 88100 35236 88156
rect 35236 88100 35240 88156
rect 35176 88096 35240 88100
rect 19576 87612 19640 87616
rect 19576 87556 19580 87612
rect 19580 87556 19636 87612
rect 19636 87556 19640 87612
rect 19576 87552 19640 87556
rect 19656 87612 19720 87616
rect 19656 87556 19660 87612
rect 19660 87556 19716 87612
rect 19716 87556 19720 87612
rect 19656 87552 19720 87556
rect 19736 87612 19800 87616
rect 19736 87556 19740 87612
rect 19740 87556 19796 87612
rect 19796 87556 19800 87612
rect 19736 87552 19800 87556
rect 19816 87612 19880 87616
rect 19816 87556 19820 87612
rect 19820 87556 19876 87612
rect 19876 87556 19880 87612
rect 19816 87552 19880 87556
rect 4216 87068 4280 87072
rect 4216 87012 4220 87068
rect 4220 87012 4276 87068
rect 4276 87012 4280 87068
rect 4216 87008 4280 87012
rect 4296 87068 4360 87072
rect 4296 87012 4300 87068
rect 4300 87012 4356 87068
rect 4356 87012 4360 87068
rect 4296 87008 4360 87012
rect 4376 87068 4440 87072
rect 4376 87012 4380 87068
rect 4380 87012 4436 87068
rect 4436 87012 4440 87068
rect 4376 87008 4440 87012
rect 4456 87068 4520 87072
rect 4456 87012 4460 87068
rect 4460 87012 4516 87068
rect 4516 87012 4520 87068
rect 4456 87008 4520 87012
rect 34936 87068 35000 87072
rect 34936 87012 34940 87068
rect 34940 87012 34996 87068
rect 34996 87012 35000 87068
rect 34936 87008 35000 87012
rect 35016 87068 35080 87072
rect 35016 87012 35020 87068
rect 35020 87012 35076 87068
rect 35076 87012 35080 87068
rect 35016 87008 35080 87012
rect 35096 87068 35160 87072
rect 35096 87012 35100 87068
rect 35100 87012 35156 87068
rect 35156 87012 35160 87068
rect 35096 87008 35160 87012
rect 35176 87068 35240 87072
rect 35176 87012 35180 87068
rect 35180 87012 35236 87068
rect 35236 87012 35240 87068
rect 35176 87008 35240 87012
rect 19576 86524 19640 86528
rect 19576 86468 19580 86524
rect 19580 86468 19636 86524
rect 19636 86468 19640 86524
rect 19576 86464 19640 86468
rect 19656 86524 19720 86528
rect 19656 86468 19660 86524
rect 19660 86468 19716 86524
rect 19716 86468 19720 86524
rect 19656 86464 19720 86468
rect 19736 86524 19800 86528
rect 19736 86468 19740 86524
rect 19740 86468 19796 86524
rect 19796 86468 19800 86524
rect 19736 86464 19800 86468
rect 19816 86524 19880 86528
rect 19816 86468 19820 86524
rect 19820 86468 19876 86524
rect 19876 86468 19880 86524
rect 19816 86464 19880 86468
rect 4216 85980 4280 85984
rect 4216 85924 4220 85980
rect 4220 85924 4276 85980
rect 4276 85924 4280 85980
rect 4216 85920 4280 85924
rect 4296 85980 4360 85984
rect 4296 85924 4300 85980
rect 4300 85924 4356 85980
rect 4356 85924 4360 85980
rect 4296 85920 4360 85924
rect 4376 85980 4440 85984
rect 4376 85924 4380 85980
rect 4380 85924 4436 85980
rect 4436 85924 4440 85980
rect 4376 85920 4440 85924
rect 4456 85980 4520 85984
rect 4456 85924 4460 85980
rect 4460 85924 4516 85980
rect 4516 85924 4520 85980
rect 4456 85920 4520 85924
rect 34936 85980 35000 85984
rect 34936 85924 34940 85980
rect 34940 85924 34996 85980
rect 34996 85924 35000 85980
rect 34936 85920 35000 85924
rect 35016 85980 35080 85984
rect 35016 85924 35020 85980
rect 35020 85924 35076 85980
rect 35076 85924 35080 85980
rect 35016 85920 35080 85924
rect 35096 85980 35160 85984
rect 35096 85924 35100 85980
rect 35100 85924 35156 85980
rect 35156 85924 35160 85980
rect 35096 85920 35160 85924
rect 35176 85980 35240 85984
rect 35176 85924 35180 85980
rect 35180 85924 35236 85980
rect 35236 85924 35240 85980
rect 35176 85920 35240 85924
rect 19576 85436 19640 85440
rect 19576 85380 19580 85436
rect 19580 85380 19636 85436
rect 19636 85380 19640 85436
rect 19576 85376 19640 85380
rect 19656 85436 19720 85440
rect 19656 85380 19660 85436
rect 19660 85380 19716 85436
rect 19716 85380 19720 85436
rect 19656 85376 19720 85380
rect 19736 85436 19800 85440
rect 19736 85380 19740 85436
rect 19740 85380 19796 85436
rect 19796 85380 19800 85436
rect 19736 85376 19800 85380
rect 19816 85436 19880 85440
rect 19816 85380 19820 85436
rect 19820 85380 19876 85436
rect 19876 85380 19880 85436
rect 19816 85376 19880 85380
rect 4216 84892 4280 84896
rect 4216 84836 4220 84892
rect 4220 84836 4276 84892
rect 4276 84836 4280 84892
rect 4216 84832 4280 84836
rect 4296 84892 4360 84896
rect 4296 84836 4300 84892
rect 4300 84836 4356 84892
rect 4356 84836 4360 84892
rect 4296 84832 4360 84836
rect 4376 84892 4440 84896
rect 4376 84836 4380 84892
rect 4380 84836 4436 84892
rect 4436 84836 4440 84892
rect 4376 84832 4440 84836
rect 4456 84892 4520 84896
rect 4456 84836 4460 84892
rect 4460 84836 4516 84892
rect 4516 84836 4520 84892
rect 4456 84832 4520 84836
rect 34936 84892 35000 84896
rect 34936 84836 34940 84892
rect 34940 84836 34996 84892
rect 34996 84836 35000 84892
rect 34936 84832 35000 84836
rect 35016 84892 35080 84896
rect 35016 84836 35020 84892
rect 35020 84836 35076 84892
rect 35076 84836 35080 84892
rect 35016 84832 35080 84836
rect 35096 84892 35160 84896
rect 35096 84836 35100 84892
rect 35100 84836 35156 84892
rect 35156 84836 35160 84892
rect 35096 84832 35160 84836
rect 35176 84892 35240 84896
rect 35176 84836 35180 84892
rect 35180 84836 35236 84892
rect 35236 84836 35240 84892
rect 35176 84832 35240 84836
rect 19576 84348 19640 84352
rect 19576 84292 19580 84348
rect 19580 84292 19636 84348
rect 19636 84292 19640 84348
rect 19576 84288 19640 84292
rect 19656 84348 19720 84352
rect 19656 84292 19660 84348
rect 19660 84292 19716 84348
rect 19716 84292 19720 84348
rect 19656 84288 19720 84292
rect 19736 84348 19800 84352
rect 19736 84292 19740 84348
rect 19740 84292 19796 84348
rect 19796 84292 19800 84348
rect 19736 84288 19800 84292
rect 19816 84348 19880 84352
rect 19816 84292 19820 84348
rect 19820 84292 19876 84348
rect 19876 84292 19880 84348
rect 19816 84288 19880 84292
rect 4216 83804 4280 83808
rect 4216 83748 4220 83804
rect 4220 83748 4276 83804
rect 4276 83748 4280 83804
rect 4216 83744 4280 83748
rect 4296 83804 4360 83808
rect 4296 83748 4300 83804
rect 4300 83748 4356 83804
rect 4356 83748 4360 83804
rect 4296 83744 4360 83748
rect 4376 83804 4440 83808
rect 4376 83748 4380 83804
rect 4380 83748 4436 83804
rect 4436 83748 4440 83804
rect 4376 83744 4440 83748
rect 4456 83804 4520 83808
rect 4456 83748 4460 83804
rect 4460 83748 4516 83804
rect 4516 83748 4520 83804
rect 4456 83744 4520 83748
rect 34936 83804 35000 83808
rect 34936 83748 34940 83804
rect 34940 83748 34996 83804
rect 34996 83748 35000 83804
rect 34936 83744 35000 83748
rect 35016 83804 35080 83808
rect 35016 83748 35020 83804
rect 35020 83748 35076 83804
rect 35076 83748 35080 83804
rect 35016 83744 35080 83748
rect 35096 83804 35160 83808
rect 35096 83748 35100 83804
rect 35100 83748 35156 83804
rect 35156 83748 35160 83804
rect 35096 83744 35160 83748
rect 35176 83804 35240 83808
rect 35176 83748 35180 83804
rect 35180 83748 35236 83804
rect 35236 83748 35240 83804
rect 35176 83744 35240 83748
rect 19576 83260 19640 83264
rect 19576 83204 19580 83260
rect 19580 83204 19636 83260
rect 19636 83204 19640 83260
rect 19576 83200 19640 83204
rect 19656 83260 19720 83264
rect 19656 83204 19660 83260
rect 19660 83204 19716 83260
rect 19716 83204 19720 83260
rect 19656 83200 19720 83204
rect 19736 83260 19800 83264
rect 19736 83204 19740 83260
rect 19740 83204 19796 83260
rect 19796 83204 19800 83260
rect 19736 83200 19800 83204
rect 19816 83260 19880 83264
rect 19816 83204 19820 83260
rect 19820 83204 19876 83260
rect 19876 83204 19880 83260
rect 19816 83200 19880 83204
rect 4216 82716 4280 82720
rect 4216 82660 4220 82716
rect 4220 82660 4276 82716
rect 4276 82660 4280 82716
rect 4216 82656 4280 82660
rect 4296 82716 4360 82720
rect 4296 82660 4300 82716
rect 4300 82660 4356 82716
rect 4356 82660 4360 82716
rect 4296 82656 4360 82660
rect 4376 82716 4440 82720
rect 4376 82660 4380 82716
rect 4380 82660 4436 82716
rect 4436 82660 4440 82716
rect 4376 82656 4440 82660
rect 4456 82716 4520 82720
rect 4456 82660 4460 82716
rect 4460 82660 4516 82716
rect 4516 82660 4520 82716
rect 4456 82656 4520 82660
rect 34936 82716 35000 82720
rect 34936 82660 34940 82716
rect 34940 82660 34996 82716
rect 34996 82660 35000 82716
rect 34936 82656 35000 82660
rect 35016 82716 35080 82720
rect 35016 82660 35020 82716
rect 35020 82660 35076 82716
rect 35076 82660 35080 82716
rect 35016 82656 35080 82660
rect 35096 82716 35160 82720
rect 35096 82660 35100 82716
rect 35100 82660 35156 82716
rect 35156 82660 35160 82716
rect 35096 82656 35160 82660
rect 35176 82716 35240 82720
rect 35176 82660 35180 82716
rect 35180 82660 35236 82716
rect 35236 82660 35240 82716
rect 35176 82656 35240 82660
rect 19576 82172 19640 82176
rect 19576 82116 19580 82172
rect 19580 82116 19636 82172
rect 19636 82116 19640 82172
rect 19576 82112 19640 82116
rect 19656 82172 19720 82176
rect 19656 82116 19660 82172
rect 19660 82116 19716 82172
rect 19716 82116 19720 82172
rect 19656 82112 19720 82116
rect 19736 82172 19800 82176
rect 19736 82116 19740 82172
rect 19740 82116 19796 82172
rect 19796 82116 19800 82172
rect 19736 82112 19800 82116
rect 19816 82172 19880 82176
rect 19816 82116 19820 82172
rect 19820 82116 19876 82172
rect 19876 82116 19880 82172
rect 19816 82112 19880 82116
rect 4216 81628 4280 81632
rect 4216 81572 4220 81628
rect 4220 81572 4276 81628
rect 4276 81572 4280 81628
rect 4216 81568 4280 81572
rect 4296 81628 4360 81632
rect 4296 81572 4300 81628
rect 4300 81572 4356 81628
rect 4356 81572 4360 81628
rect 4296 81568 4360 81572
rect 4376 81628 4440 81632
rect 4376 81572 4380 81628
rect 4380 81572 4436 81628
rect 4436 81572 4440 81628
rect 4376 81568 4440 81572
rect 4456 81628 4520 81632
rect 4456 81572 4460 81628
rect 4460 81572 4516 81628
rect 4516 81572 4520 81628
rect 4456 81568 4520 81572
rect 34936 81628 35000 81632
rect 34936 81572 34940 81628
rect 34940 81572 34996 81628
rect 34996 81572 35000 81628
rect 34936 81568 35000 81572
rect 35016 81628 35080 81632
rect 35016 81572 35020 81628
rect 35020 81572 35076 81628
rect 35076 81572 35080 81628
rect 35016 81568 35080 81572
rect 35096 81628 35160 81632
rect 35096 81572 35100 81628
rect 35100 81572 35156 81628
rect 35156 81572 35160 81628
rect 35096 81568 35160 81572
rect 35176 81628 35240 81632
rect 35176 81572 35180 81628
rect 35180 81572 35236 81628
rect 35236 81572 35240 81628
rect 35176 81568 35240 81572
rect 19576 81084 19640 81088
rect 19576 81028 19580 81084
rect 19580 81028 19636 81084
rect 19636 81028 19640 81084
rect 19576 81024 19640 81028
rect 19656 81084 19720 81088
rect 19656 81028 19660 81084
rect 19660 81028 19716 81084
rect 19716 81028 19720 81084
rect 19656 81024 19720 81028
rect 19736 81084 19800 81088
rect 19736 81028 19740 81084
rect 19740 81028 19796 81084
rect 19796 81028 19800 81084
rect 19736 81024 19800 81028
rect 19816 81084 19880 81088
rect 19816 81028 19820 81084
rect 19820 81028 19876 81084
rect 19876 81028 19880 81084
rect 19816 81024 19880 81028
rect 4216 80540 4280 80544
rect 4216 80484 4220 80540
rect 4220 80484 4276 80540
rect 4276 80484 4280 80540
rect 4216 80480 4280 80484
rect 4296 80540 4360 80544
rect 4296 80484 4300 80540
rect 4300 80484 4356 80540
rect 4356 80484 4360 80540
rect 4296 80480 4360 80484
rect 4376 80540 4440 80544
rect 4376 80484 4380 80540
rect 4380 80484 4436 80540
rect 4436 80484 4440 80540
rect 4376 80480 4440 80484
rect 4456 80540 4520 80544
rect 4456 80484 4460 80540
rect 4460 80484 4516 80540
rect 4516 80484 4520 80540
rect 4456 80480 4520 80484
rect 19576 79996 19640 80000
rect 19576 79940 19580 79996
rect 19580 79940 19636 79996
rect 19636 79940 19640 79996
rect 19576 79936 19640 79940
rect 19656 79996 19720 80000
rect 19656 79940 19660 79996
rect 19660 79940 19716 79996
rect 19716 79940 19720 79996
rect 19656 79936 19720 79940
rect 19736 79996 19800 80000
rect 19736 79940 19740 79996
rect 19740 79940 19796 79996
rect 19796 79940 19800 79996
rect 19736 79936 19800 79940
rect 19816 79996 19880 80000
rect 19816 79940 19820 79996
rect 19820 79940 19876 79996
rect 19876 79940 19880 79996
rect 19816 79936 19880 79940
rect 4216 79452 4280 79456
rect 4216 79396 4220 79452
rect 4220 79396 4276 79452
rect 4276 79396 4280 79452
rect 4216 79392 4280 79396
rect 4296 79452 4360 79456
rect 4296 79396 4300 79452
rect 4300 79396 4356 79452
rect 4356 79396 4360 79452
rect 4296 79392 4360 79396
rect 4376 79452 4440 79456
rect 4376 79396 4380 79452
rect 4380 79396 4436 79452
rect 4436 79396 4440 79452
rect 4376 79392 4440 79396
rect 4456 79452 4520 79456
rect 4456 79396 4460 79452
rect 4460 79396 4516 79452
rect 4516 79396 4520 79452
rect 4456 79392 4520 79396
rect 34936 80540 35000 80544
rect 34936 80484 34940 80540
rect 34940 80484 34996 80540
rect 34996 80484 35000 80540
rect 34936 80480 35000 80484
rect 35016 80540 35080 80544
rect 35016 80484 35020 80540
rect 35020 80484 35076 80540
rect 35076 80484 35080 80540
rect 35016 80480 35080 80484
rect 35096 80540 35160 80544
rect 35096 80484 35100 80540
rect 35100 80484 35156 80540
rect 35156 80484 35160 80540
rect 35096 80480 35160 80484
rect 35176 80540 35240 80544
rect 35176 80484 35180 80540
rect 35180 80484 35236 80540
rect 35236 80484 35240 80540
rect 35176 80480 35240 80484
rect 19576 78908 19640 78912
rect 19576 78852 19580 78908
rect 19580 78852 19636 78908
rect 19636 78852 19640 78908
rect 19576 78848 19640 78852
rect 19656 78908 19720 78912
rect 19656 78852 19660 78908
rect 19660 78852 19716 78908
rect 19716 78852 19720 78908
rect 19656 78848 19720 78852
rect 19736 78908 19800 78912
rect 19736 78852 19740 78908
rect 19740 78852 19796 78908
rect 19796 78852 19800 78908
rect 19736 78848 19800 78852
rect 19816 78908 19880 78912
rect 19816 78852 19820 78908
rect 19820 78852 19876 78908
rect 19876 78852 19880 78908
rect 19816 78848 19880 78852
rect 34936 79452 35000 79456
rect 34936 79396 34940 79452
rect 34940 79396 34996 79452
rect 34996 79396 35000 79452
rect 34936 79392 35000 79396
rect 35016 79452 35080 79456
rect 35016 79396 35020 79452
rect 35020 79396 35076 79452
rect 35076 79396 35080 79452
rect 35016 79392 35080 79396
rect 35096 79452 35160 79456
rect 35096 79396 35100 79452
rect 35100 79396 35156 79452
rect 35156 79396 35160 79452
rect 35096 79392 35160 79396
rect 35176 79452 35240 79456
rect 35176 79396 35180 79452
rect 35180 79396 35236 79452
rect 35236 79396 35240 79452
rect 35176 79392 35240 79396
rect 4216 78364 4280 78368
rect 4216 78308 4220 78364
rect 4220 78308 4276 78364
rect 4276 78308 4280 78364
rect 4216 78304 4280 78308
rect 4296 78364 4360 78368
rect 4296 78308 4300 78364
rect 4300 78308 4356 78364
rect 4356 78308 4360 78364
rect 4296 78304 4360 78308
rect 4376 78364 4440 78368
rect 4376 78308 4380 78364
rect 4380 78308 4436 78364
rect 4436 78308 4440 78364
rect 4376 78304 4440 78308
rect 4456 78364 4520 78368
rect 4456 78308 4460 78364
rect 4460 78308 4516 78364
rect 4516 78308 4520 78364
rect 4456 78304 4520 78308
rect 34936 78364 35000 78368
rect 34936 78308 34940 78364
rect 34940 78308 34996 78364
rect 34996 78308 35000 78364
rect 34936 78304 35000 78308
rect 35016 78364 35080 78368
rect 35016 78308 35020 78364
rect 35020 78308 35076 78364
rect 35076 78308 35080 78364
rect 35016 78304 35080 78308
rect 35096 78364 35160 78368
rect 35096 78308 35100 78364
rect 35100 78308 35156 78364
rect 35156 78308 35160 78364
rect 35096 78304 35160 78308
rect 35176 78364 35240 78368
rect 35176 78308 35180 78364
rect 35180 78308 35236 78364
rect 35236 78308 35240 78364
rect 35176 78304 35240 78308
rect 19576 77820 19640 77824
rect 19576 77764 19580 77820
rect 19580 77764 19636 77820
rect 19636 77764 19640 77820
rect 19576 77760 19640 77764
rect 19656 77820 19720 77824
rect 19656 77764 19660 77820
rect 19660 77764 19716 77820
rect 19716 77764 19720 77820
rect 19656 77760 19720 77764
rect 19736 77820 19800 77824
rect 19736 77764 19740 77820
rect 19740 77764 19796 77820
rect 19796 77764 19800 77820
rect 19736 77760 19800 77764
rect 19816 77820 19880 77824
rect 19816 77764 19820 77820
rect 19820 77764 19876 77820
rect 19876 77764 19880 77820
rect 19816 77760 19880 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 34936 77276 35000 77280
rect 34936 77220 34940 77276
rect 34940 77220 34996 77276
rect 34996 77220 35000 77276
rect 34936 77216 35000 77220
rect 35016 77276 35080 77280
rect 35016 77220 35020 77276
rect 35020 77220 35076 77276
rect 35076 77220 35080 77276
rect 35016 77216 35080 77220
rect 35096 77276 35160 77280
rect 35096 77220 35100 77276
rect 35100 77220 35156 77276
rect 35156 77220 35160 77276
rect 35096 77216 35160 77220
rect 35176 77276 35240 77280
rect 35176 77220 35180 77276
rect 35180 77220 35236 77276
rect 35236 77220 35240 77276
rect 35176 77216 35240 77220
rect 19576 76732 19640 76736
rect 19576 76676 19580 76732
rect 19580 76676 19636 76732
rect 19636 76676 19640 76732
rect 19576 76672 19640 76676
rect 19656 76732 19720 76736
rect 19656 76676 19660 76732
rect 19660 76676 19716 76732
rect 19716 76676 19720 76732
rect 19656 76672 19720 76676
rect 19736 76732 19800 76736
rect 19736 76676 19740 76732
rect 19740 76676 19796 76732
rect 19796 76676 19800 76732
rect 19736 76672 19800 76676
rect 19816 76732 19880 76736
rect 19816 76676 19820 76732
rect 19820 76676 19876 76732
rect 19876 76676 19880 76732
rect 19816 76672 19880 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 34936 76188 35000 76192
rect 34936 76132 34940 76188
rect 34940 76132 34996 76188
rect 34996 76132 35000 76188
rect 34936 76128 35000 76132
rect 35016 76188 35080 76192
rect 35016 76132 35020 76188
rect 35020 76132 35076 76188
rect 35076 76132 35080 76188
rect 35016 76128 35080 76132
rect 35096 76188 35160 76192
rect 35096 76132 35100 76188
rect 35100 76132 35156 76188
rect 35156 76132 35160 76188
rect 35096 76128 35160 76132
rect 35176 76188 35240 76192
rect 35176 76132 35180 76188
rect 35180 76132 35236 76188
rect 35236 76132 35240 76188
rect 35176 76128 35240 76132
rect 19576 75644 19640 75648
rect 19576 75588 19580 75644
rect 19580 75588 19636 75644
rect 19636 75588 19640 75644
rect 19576 75584 19640 75588
rect 19656 75644 19720 75648
rect 19656 75588 19660 75644
rect 19660 75588 19716 75644
rect 19716 75588 19720 75644
rect 19656 75584 19720 75588
rect 19736 75644 19800 75648
rect 19736 75588 19740 75644
rect 19740 75588 19796 75644
rect 19796 75588 19800 75644
rect 19736 75584 19800 75588
rect 19816 75644 19880 75648
rect 19816 75588 19820 75644
rect 19820 75588 19876 75644
rect 19876 75588 19880 75644
rect 19816 75584 19880 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 34936 75100 35000 75104
rect 34936 75044 34940 75100
rect 34940 75044 34996 75100
rect 34996 75044 35000 75100
rect 34936 75040 35000 75044
rect 35016 75100 35080 75104
rect 35016 75044 35020 75100
rect 35020 75044 35076 75100
rect 35076 75044 35080 75100
rect 35016 75040 35080 75044
rect 35096 75100 35160 75104
rect 35096 75044 35100 75100
rect 35100 75044 35156 75100
rect 35156 75044 35160 75100
rect 35096 75040 35160 75044
rect 35176 75100 35240 75104
rect 35176 75044 35180 75100
rect 35180 75044 35236 75100
rect 35236 75044 35240 75100
rect 35176 75040 35240 75044
rect 19576 74556 19640 74560
rect 19576 74500 19580 74556
rect 19580 74500 19636 74556
rect 19636 74500 19640 74556
rect 19576 74496 19640 74500
rect 19656 74556 19720 74560
rect 19656 74500 19660 74556
rect 19660 74500 19716 74556
rect 19716 74500 19720 74556
rect 19656 74496 19720 74500
rect 19736 74556 19800 74560
rect 19736 74500 19740 74556
rect 19740 74500 19796 74556
rect 19796 74500 19800 74556
rect 19736 74496 19800 74500
rect 19816 74556 19880 74560
rect 19816 74500 19820 74556
rect 19820 74500 19876 74556
rect 19876 74500 19880 74556
rect 19816 74496 19880 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 34936 74012 35000 74016
rect 34936 73956 34940 74012
rect 34940 73956 34996 74012
rect 34996 73956 35000 74012
rect 34936 73952 35000 73956
rect 35016 74012 35080 74016
rect 35016 73956 35020 74012
rect 35020 73956 35076 74012
rect 35076 73956 35080 74012
rect 35016 73952 35080 73956
rect 35096 74012 35160 74016
rect 35096 73956 35100 74012
rect 35100 73956 35156 74012
rect 35156 73956 35160 74012
rect 35096 73952 35160 73956
rect 35176 74012 35240 74016
rect 35176 73956 35180 74012
rect 35180 73956 35236 74012
rect 35236 73956 35240 74012
rect 35176 73952 35240 73956
rect 19576 73468 19640 73472
rect 19576 73412 19580 73468
rect 19580 73412 19636 73468
rect 19636 73412 19640 73468
rect 19576 73408 19640 73412
rect 19656 73468 19720 73472
rect 19656 73412 19660 73468
rect 19660 73412 19716 73468
rect 19716 73412 19720 73468
rect 19656 73408 19720 73412
rect 19736 73468 19800 73472
rect 19736 73412 19740 73468
rect 19740 73412 19796 73468
rect 19796 73412 19800 73468
rect 19736 73408 19800 73412
rect 19816 73468 19880 73472
rect 19816 73412 19820 73468
rect 19820 73412 19876 73468
rect 19876 73412 19880 73468
rect 19816 73408 19880 73412
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 34936 72924 35000 72928
rect 34936 72868 34940 72924
rect 34940 72868 34996 72924
rect 34996 72868 35000 72924
rect 34936 72864 35000 72868
rect 35016 72924 35080 72928
rect 35016 72868 35020 72924
rect 35020 72868 35076 72924
rect 35076 72868 35080 72924
rect 35016 72864 35080 72868
rect 35096 72924 35160 72928
rect 35096 72868 35100 72924
rect 35100 72868 35156 72924
rect 35156 72868 35160 72924
rect 35096 72864 35160 72868
rect 35176 72924 35240 72928
rect 35176 72868 35180 72924
rect 35180 72868 35236 72924
rect 35236 72868 35240 72924
rect 35176 72864 35240 72868
rect 19576 72380 19640 72384
rect 19576 72324 19580 72380
rect 19580 72324 19636 72380
rect 19636 72324 19640 72380
rect 19576 72320 19640 72324
rect 19656 72380 19720 72384
rect 19656 72324 19660 72380
rect 19660 72324 19716 72380
rect 19716 72324 19720 72380
rect 19656 72320 19720 72324
rect 19736 72380 19800 72384
rect 19736 72324 19740 72380
rect 19740 72324 19796 72380
rect 19796 72324 19800 72380
rect 19736 72320 19800 72324
rect 19816 72380 19880 72384
rect 19816 72324 19820 72380
rect 19820 72324 19876 72380
rect 19876 72324 19880 72380
rect 19816 72320 19880 72324
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 34936 71836 35000 71840
rect 34936 71780 34940 71836
rect 34940 71780 34996 71836
rect 34996 71780 35000 71836
rect 34936 71776 35000 71780
rect 35016 71836 35080 71840
rect 35016 71780 35020 71836
rect 35020 71780 35076 71836
rect 35076 71780 35080 71836
rect 35016 71776 35080 71780
rect 35096 71836 35160 71840
rect 35096 71780 35100 71836
rect 35100 71780 35156 71836
rect 35156 71780 35160 71836
rect 35096 71776 35160 71780
rect 35176 71836 35240 71840
rect 35176 71780 35180 71836
rect 35180 71780 35236 71836
rect 35236 71780 35240 71836
rect 35176 71776 35240 71780
rect 19576 71292 19640 71296
rect 19576 71236 19580 71292
rect 19580 71236 19636 71292
rect 19636 71236 19640 71292
rect 19576 71232 19640 71236
rect 19656 71292 19720 71296
rect 19656 71236 19660 71292
rect 19660 71236 19716 71292
rect 19716 71236 19720 71292
rect 19656 71232 19720 71236
rect 19736 71292 19800 71296
rect 19736 71236 19740 71292
rect 19740 71236 19796 71292
rect 19796 71236 19800 71292
rect 19736 71232 19800 71236
rect 19816 71292 19880 71296
rect 19816 71236 19820 71292
rect 19820 71236 19876 71292
rect 19876 71236 19880 71292
rect 19816 71232 19880 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 34936 70748 35000 70752
rect 34936 70692 34940 70748
rect 34940 70692 34996 70748
rect 34996 70692 35000 70748
rect 34936 70688 35000 70692
rect 35016 70748 35080 70752
rect 35016 70692 35020 70748
rect 35020 70692 35076 70748
rect 35076 70692 35080 70748
rect 35016 70688 35080 70692
rect 35096 70748 35160 70752
rect 35096 70692 35100 70748
rect 35100 70692 35156 70748
rect 35156 70692 35160 70748
rect 35096 70688 35160 70692
rect 35176 70748 35240 70752
rect 35176 70692 35180 70748
rect 35180 70692 35236 70748
rect 35236 70692 35240 70748
rect 35176 70688 35240 70692
rect 19576 70204 19640 70208
rect 19576 70148 19580 70204
rect 19580 70148 19636 70204
rect 19636 70148 19640 70204
rect 19576 70144 19640 70148
rect 19656 70204 19720 70208
rect 19656 70148 19660 70204
rect 19660 70148 19716 70204
rect 19716 70148 19720 70204
rect 19656 70144 19720 70148
rect 19736 70204 19800 70208
rect 19736 70148 19740 70204
rect 19740 70148 19796 70204
rect 19796 70148 19800 70204
rect 19736 70144 19800 70148
rect 19816 70204 19880 70208
rect 19816 70148 19820 70204
rect 19820 70148 19876 70204
rect 19876 70148 19880 70204
rect 19816 70144 19880 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 34936 69660 35000 69664
rect 34936 69604 34940 69660
rect 34940 69604 34996 69660
rect 34996 69604 35000 69660
rect 34936 69600 35000 69604
rect 35016 69660 35080 69664
rect 35016 69604 35020 69660
rect 35020 69604 35076 69660
rect 35076 69604 35080 69660
rect 35016 69600 35080 69604
rect 35096 69660 35160 69664
rect 35096 69604 35100 69660
rect 35100 69604 35156 69660
rect 35156 69604 35160 69660
rect 35096 69600 35160 69604
rect 35176 69660 35240 69664
rect 35176 69604 35180 69660
rect 35180 69604 35236 69660
rect 35236 69604 35240 69660
rect 35176 69600 35240 69604
rect 19576 69116 19640 69120
rect 19576 69060 19580 69116
rect 19580 69060 19636 69116
rect 19636 69060 19640 69116
rect 19576 69056 19640 69060
rect 19656 69116 19720 69120
rect 19656 69060 19660 69116
rect 19660 69060 19716 69116
rect 19716 69060 19720 69116
rect 19656 69056 19720 69060
rect 19736 69116 19800 69120
rect 19736 69060 19740 69116
rect 19740 69060 19796 69116
rect 19796 69060 19800 69116
rect 19736 69056 19800 69060
rect 19816 69116 19880 69120
rect 19816 69060 19820 69116
rect 19820 69060 19876 69116
rect 19876 69060 19880 69116
rect 19816 69056 19880 69060
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 34936 68572 35000 68576
rect 34936 68516 34940 68572
rect 34940 68516 34996 68572
rect 34996 68516 35000 68572
rect 34936 68512 35000 68516
rect 35016 68572 35080 68576
rect 35016 68516 35020 68572
rect 35020 68516 35076 68572
rect 35076 68516 35080 68572
rect 35016 68512 35080 68516
rect 35096 68572 35160 68576
rect 35096 68516 35100 68572
rect 35100 68516 35156 68572
rect 35156 68516 35160 68572
rect 35096 68512 35160 68516
rect 35176 68572 35240 68576
rect 35176 68516 35180 68572
rect 35180 68516 35236 68572
rect 35236 68516 35240 68572
rect 35176 68512 35240 68516
rect 19576 68028 19640 68032
rect 19576 67972 19580 68028
rect 19580 67972 19636 68028
rect 19636 67972 19640 68028
rect 19576 67968 19640 67972
rect 19656 68028 19720 68032
rect 19656 67972 19660 68028
rect 19660 67972 19716 68028
rect 19716 67972 19720 68028
rect 19656 67968 19720 67972
rect 19736 68028 19800 68032
rect 19736 67972 19740 68028
rect 19740 67972 19796 68028
rect 19796 67972 19800 68028
rect 19736 67968 19800 67972
rect 19816 68028 19880 68032
rect 19816 67972 19820 68028
rect 19820 67972 19876 68028
rect 19876 67972 19880 68028
rect 19816 67968 19880 67972
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 34936 67484 35000 67488
rect 34936 67428 34940 67484
rect 34940 67428 34996 67484
rect 34996 67428 35000 67484
rect 34936 67424 35000 67428
rect 35016 67484 35080 67488
rect 35016 67428 35020 67484
rect 35020 67428 35076 67484
rect 35076 67428 35080 67484
rect 35016 67424 35080 67428
rect 35096 67484 35160 67488
rect 35096 67428 35100 67484
rect 35100 67428 35156 67484
rect 35156 67428 35160 67484
rect 35096 67424 35160 67428
rect 35176 67484 35240 67488
rect 35176 67428 35180 67484
rect 35180 67428 35236 67484
rect 35236 67428 35240 67484
rect 35176 67424 35240 67428
rect 19576 66940 19640 66944
rect 19576 66884 19580 66940
rect 19580 66884 19636 66940
rect 19636 66884 19640 66940
rect 19576 66880 19640 66884
rect 19656 66940 19720 66944
rect 19656 66884 19660 66940
rect 19660 66884 19716 66940
rect 19716 66884 19720 66940
rect 19656 66880 19720 66884
rect 19736 66940 19800 66944
rect 19736 66884 19740 66940
rect 19740 66884 19796 66940
rect 19796 66884 19800 66940
rect 19736 66880 19800 66884
rect 19816 66940 19880 66944
rect 19816 66884 19820 66940
rect 19820 66884 19876 66940
rect 19876 66884 19880 66940
rect 19816 66880 19880 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 34936 66396 35000 66400
rect 34936 66340 34940 66396
rect 34940 66340 34996 66396
rect 34996 66340 35000 66396
rect 34936 66336 35000 66340
rect 35016 66396 35080 66400
rect 35016 66340 35020 66396
rect 35020 66340 35076 66396
rect 35076 66340 35080 66396
rect 35016 66336 35080 66340
rect 35096 66396 35160 66400
rect 35096 66340 35100 66396
rect 35100 66340 35156 66396
rect 35156 66340 35160 66396
rect 35096 66336 35160 66340
rect 35176 66396 35240 66400
rect 35176 66340 35180 66396
rect 35180 66340 35236 66396
rect 35236 66340 35240 66396
rect 35176 66336 35240 66340
rect 19576 65852 19640 65856
rect 19576 65796 19580 65852
rect 19580 65796 19636 65852
rect 19636 65796 19640 65852
rect 19576 65792 19640 65796
rect 19656 65852 19720 65856
rect 19656 65796 19660 65852
rect 19660 65796 19716 65852
rect 19716 65796 19720 65852
rect 19656 65792 19720 65796
rect 19736 65852 19800 65856
rect 19736 65796 19740 65852
rect 19740 65796 19796 65852
rect 19796 65796 19800 65852
rect 19736 65792 19800 65796
rect 19816 65852 19880 65856
rect 19816 65796 19820 65852
rect 19820 65796 19876 65852
rect 19876 65796 19880 65852
rect 19816 65792 19880 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 34936 65308 35000 65312
rect 34936 65252 34940 65308
rect 34940 65252 34996 65308
rect 34996 65252 35000 65308
rect 34936 65248 35000 65252
rect 35016 65308 35080 65312
rect 35016 65252 35020 65308
rect 35020 65252 35076 65308
rect 35076 65252 35080 65308
rect 35016 65248 35080 65252
rect 35096 65308 35160 65312
rect 35096 65252 35100 65308
rect 35100 65252 35156 65308
rect 35156 65252 35160 65308
rect 35096 65248 35160 65252
rect 35176 65308 35240 65312
rect 35176 65252 35180 65308
rect 35180 65252 35236 65308
rect 35236 65252 35240 65308
rect 35176 65248 35240 65252
rect 19576 64764 19640 64768
rect 19576 64708 19580 64764
rect 19580 64708 19636 64764
rect 19636 64708 19640 64764
rect 19576 64704 19640 64708
rect 19656 64764 19720 64768
rect 19656 64708 19660 64764
rect 19660 64708 19716 64764
rect 19716 64708 19720 64764
rect 19656 64704 19720 64708
rect 19736 64764 19800 64768
rect 19736 64708 19740 64764
rect 19740 64708 19796 64764
rect 19796 64708 19800 64764
rect 19736 64704 19800 64708
rect 19816 64764 19880 64768
rect 19816 64708 19820 64764
rect 19820 64708 19876 64764
rect 19876 64708 19880 64764
rect 19816 64704 19880 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 34936 64220 35000 64224
rect 34936 64164 34940 64220
rect 34940 64164 34996 64220
rect 34996 64164 35000 64220
rect 34936 64160 35000 64164
rect 35016 64220 35080 64224
rect 35016 64164 35020 64220
rect 35020 64164 35076 64220
rect 35076 64164 35080 64220
rect 35016 64160 35080 64164
rect 35096 64220 35160 64224
rect 35096 64164 35100 64220
rect 35100 64164 35156 64220
rect 35156 64164 35160 64220
rect 35096 64160 35160 64164
rect 35176 64220 35240 64224
rect 35176 64164 35180 64220
rect 35180 64164 35236 64220
rect 35236 64164 35240 64220
rect 35176 64160 35240 64164
rect 19576 63676 19640 63680
rect 19576 63620 19580 63676
rect 19580 63620 19636 63676
rect 19636 63620 19640 63676
rect 19576 63616 19640 63620
rect 19656 63676 19720 63680
rect 19656 63620 19660 63676
rect 19660 63620 19716 63676
rect 19716 63620 19720 63676
rect 19656 63616 19720 63620
rect 19736 63676 19800 63680
rect 19736 63620 19740 63676
rect 19740 63620 19796 63676
rect 19796 63620 19800 63676
rect 19736 63616 19800 63620
rect 19816 63676 19880 63680
rect 19816 63620 19820 63676
rect 19820 63620 19876 63676
rect 19876 63620 19880 63676
rect 19816 63616 19880 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 34936 63132 35000 63136
rect 34936 63076 34940 63132
rect 34940 63076 34996 63132
rect 34996 63076 35000 63132
rect 34936 63072 35000 63076
rect 35016 63132 35080 63136
rect 35016 63076 35020 63132
rect 35020 63076 35076 63132
rect 35076 63076 35080 63132
rect 35016 63072 35080 63076
rect 35096 63132 35160 63136
rect 35096 63076 35100 63132
rect 35100 63076 35156 63132
rect 35156 63076 35160 63132
rect 35096 63072 35160 63076
rect 35176 63132 35240 63136
rect 35176 63076 35180 63132
rect 35180 63076 35236 63132
rect 35236 63076 35240 63132
rect 35176 63072 35240 63076
rect 19576 62588 19640 62592
rect 19576 62532 19580 62588
rect 19580 62532 19636 62588
rect 19636 62532 19640 62588
rect 19576 62528 19640 62532
rect 19656 62588 19720 62592
rect 19656 62532 19660 62588
rect 19660 62532 19716 62588
rect 19716 62532 19720 62588
rect 19656 62528 19720 62532
rect 19736 62588 19800 62592
rect 19736 62532 19740 62588
rect 19740 62532 19796 62588
rect 19796 62532 19800 62588
rect 19736 62528 19800 62532
rect 19816 62588 19880 62592
rect 19816 62532 19820 62588
rect 19820 62532 19876 62588
rect 19876 62532 19880 62588
rect 19816 62528 19880 62532
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 34936 62044 35000 62048
rect 34936 61988 34940 62044
rect 34940 61988 34996 62044
rect 34996 61988 35000 62044
rect 34936 61984 35000 61988
rect 35016 62044 35080 62048
rect 35016 61988 35020 62044
rect 35020 61988 35076 62044
rect 35076 61988 35080 62044
rect 35016 61984 35080 61988
rect 35096 62044 35160 62048
rect 35096 61988 35100 62044
rect 35100 61988 35156 62044
rect 35156 61988 35160 62044
rect 35096 61984 35160 61988
rect 35176 62044 35240 62048
rect 35176 61988 35180 62044
rect 35180 61988 35236 62044
rect 35236 61988 35240 62044
rect 35176 61984 35240 61988
rect 19576 61500 19640 61504
rect 19576 61444 19580 61500
rect 19580 61444 19636 61500
rect 19636 61444 19640 61500
rect 19576 61440 19640 61444
rect 19656 61500 19720 61504
rect 19656 61444 19660 61500
rect 19660 61444 19716 61500
rect 19716 61444 19720 61500
rect 19656 61440 19720 61444
rect 19736 61500 19800 61504
rect 19736 61444 19740 61500
rect 19740 61444 19796 61500
rect 19796 61444 19800 61500
rect 19736 61440 19800 61444
rect 19816 61500 19880 61504
rect 19816 61444 19820 61500
rect 19820 61444 19876 61500
rect 19876 61444 19880 61500
rect 19816 61440 19880 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 34936 60956 35000 60960
rect 34936 60900 34940 60956
rect 34940 60900 34996 60956
rect 34996 60900 35000 60956
rect 34936 60896 35000 60900
rect 35016 60956 35080 60960
rect 35016 60900 35020 60956
rect 35020 60900 35076 60956
rect 35076 60900 35080 60956
rect 35016 60896 35080 60900
rect 35096 60956 35160 60960
rect 35096 60900 35100 60956
rect 35100 60900 35156 60956
rect 35156 60900 35160 60956
rect 35096 60896 35160 60900
rect 35176 60956 35240 60960
rect 35176 60900 35180 60956
rect 35180 60900 35236 60956
rect 35236 60900 35240 60956
rect 35176 60896 35240 60900
rect 19576 60412 19640 60416
rect 19576 60356 19580 60412
rect 19580 60356 19636 60412
rect 19636 60356 19640 60412
rect 19576 60352 19640 60356
rect 19656 60412 19720 60416
rect 19656 60356 19660 60412
rect 19660 60356 19716 60412
rect 19716 60356 19720 60412
rect 19656 60352 19720 60356
rect 19736 60412 19800 60416
rect 19736 60356 19740 60412
rect 19740 60356 19796 60412
rect 19796 60356 19800 60412
rect 19736 60352 19800 60356
rect 19816 60412 19880 60416
rect 19816 60356 19820 60412
rect 19820 60356 19876 60412
rect 19876 60356 19880 60412
rect 19816 60352 19880 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 34936 59868 35000 59872
rect 34936 59812 34940 59868
rect 34940 59812 34996 59868
rect 34996 59812 35000 59868
rect 34936 59808 35000 59812
rect 35016 59868 35080 59872
rect 35016 59812 35020 59868
rect 35020 59812 35076 59868
rect 35076 59812 35080 59868
rect 35016 59808 35080 59812
rect 35096 59868 35160 59872
rect 35096 59812 35100 59868
rect 35100 59812 35156 59868
rect 35156 59812 35160 59868
rect 35096 59808 35160 59812
rect 35176 59868 35240 59872
rect 35176 59812 35180 59868
rect 35180 59812 35236 59868
rect 35236 59812 35240 59868
rect 35176 59808 35240 59812
rect 19576 59324 19640 59328
rect 19576 59268 19580 59324
rect 19580 59268 19636 59324
rect 19636 59268 19640 59324
rect 19576 59264 19640 59268
rect 19656 59324 19720 59328
rect 19656 59268 19660 59324
rect 19660 59268 19716 59324
rect 19716 59268 19720 59324
rect 19656 59264 19720 59268
rect 19736 59324 19800 59328
rect 19736 59268 19740 59324
rect 19740 59268 19796 59324
rect 19796 59268 19800 59324
rect 19736 59264 19800 59268
rect 19816 59324 19880 59328
rect 19816 59268 19820 59324
rect 19820 59268 19876 59324
rect 19876 59268 19880 59324
rect 19816 59264 19880 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 34936 58780 35000 58784
rect 34936 58724 34940 58780
rect 34940 58724 34996 58780
rect 34996 58724 35000 58780
rect 34936 58720 35000 58724
rect 35016 58780 35080 58784
rect 35016 58724 35020 58780
rect 35020 58724 35076 58780
rect 35076 58724 35080 58780
rect 35016 58720 35080 58724
rect 35096 58780 35160 58784
rect 35096 58724 35100 58780
rect 35100 58724 35156 58780
rect 35156 58724 35160 58780
rect 35096 58720 35160 58724
rect 35176 58780 35240 58784
rect 35176 58724 35180 58780
rect 35180 58724 35236 58780
rect 35236 58724 35240 58780
rect 35176 58720 35240 58724
rect 19576 58236 19640 58240
rect 19576 58180 19580 58236
rect 19580 58180 19636 58236
rect 19636 58180 19640 58236
rect 19576 58176 19640 58180
rect 19656 58236 19720 58240
rect 19656 58180 19660 58236
rect 19660 58180 19716 58236
rect 19716 58180 19720 58236
rect 19656 58176 19720 58180
rect 19736 58236 19800 58240
rect 19736 58180 19740 58236
rect 19740 58180 19796 58236
rect 19796 58180 19800 58236
rect 19736 58176 19800 58180
rect 19816 58236 19880 58240
rect 19816 58180 19820 58236
rect 19820 58180 19876 58236
rect 19876 58180 19880 58236
rect 19816 58176 19880 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 117536 4528 117552
rect 4208 117472 4216 117536
rect 4280 117472 4296 117536
rect 4360 117472 4376 117536
rect 4440 117472 4456 117536
rect 4520 117472 4528 117536
rect 4208 116448 4528 117472
rect 4208 116384 4216 116448
rect 4280 116384 4296 116448
rect 4360 116384 4376 116448
rect 4440 116384 4456 116448
rect 4520 116384 4528 116448
rect 4208 115360 4528 116384
rect 4208 115296 4216 115360
rect 4280 115296 4296 115360
rect 4360 115296 4376 115360
rect 4440 115296 4456 115360
rect 4520 115296 4528 115360
rect 4208 114272 4528 115296
rect 4208 114208 4216 114272
rect 4280 114208 4296 114272
rect 4360 114208 4376 114272
rect 4440 114208 4456 114272
rect 4520 114208 4528 114272
rect 4208 113184 4528 114208
rect 4208 113120 4216 113184
rect 4280 113120 4296 113184
rect 4360 113120 4376 113184
rect 4440 113120 4456 113184
rect 4520 113120 4528 113184
rect 4208 112096 4528 113120
rect 4208 112032 4216 112096
rect 4280 112032 4296 112096
rect 4360 112032 4376 112096
rect 4440 112032 4456 112096
rect 4520 112032 4528 112096
rect 4208 111008 4528 112032
rect 4208 110944 4216 111008
rect 4280 110944 4296 111008
rect 4360 110944 4376 111008
rect 4440 110944 4456 111008
rect 4520 110944 4528 111008
rect 4208 109920 4528 110944
rect 4208 109856 4216 109920
rect 4280 109856 4296 109920
rect 4360 109856 4376 109920
rect 4440 109856 4456 109920
rect 4520 109856 4528 109920
rect 4208 108832 4528 109856
rect 4208 108768 4216 108832
rect 4280 108768 4296 108832
rect 4360 108768 4376 108832
rect 4440 108768 4456 108832
rect 4520 108768 4528 108832
rect 4208 107744 4528 108768
rect 4208 107680 4216 107744
rect 4280 107680 4296 107744
rect 4360 107680 4376 107744
rect 4440 107680 4456 107744
rect 4520 107680 4528 107744
rect 4208 106656 4528 107680
rect 4208 106592 4216 106656
rect 4280 106592 4296 106656
rect 4360 106592 4376 106656
rect 4440 106592 4456 106656
rect 4520 106592 4528 106656
rect 4208 105568 4528 106592
rect 4208 105504 4216 105568
rect 4280 105504 4296 105568
rect 4360 105504 4376 105568
rect 4440 105504 4456 105568
rect 4520 105504 4528 105568
rect 4208 104480 4528 105504
rect 4208 104416 4216 104480
rect 4280 104416 4296 104480
rect 4360 104416 4376 104480
rect 4440 104416 4456 104480
rect 4520 104416 4528 104480
rect 4208 103392 4528 104416
rect 4208 103328 4216 103392
rect 4280 103328 4296 103392
rect 4360 103328 4376 103392
rect 4440 103328 4456 103392
rect 4520 103328 4528 103392
rect 4208 102304 4528 103328
rect 4208 102240 4216 102304
rect 4280 102240 4296 102304
rect 4360 102240 4376 102304
rect 4440 102240 4456 102304
rect 4520 102240 4528 102304
rect 4208 101216 4528 102240
rect 4208 101152 4216 101216
rect 4280 101152 4296 101216
rect 4360 101152 4376 101216
rect 4440 101152 4456 101216
rect 4520 101152 4528 101216
rect 4208 100128 4528 101152
rect 4208 100064 4216 100128
rect 4280 100064 4296 100128
rect 4360 100064 4376 100128
rect 4440 100064 4456 100128
rect 4520 100064 4528 100128
rect 4208 99040 4528 100064
rect 4208 98976 4216 99040
rect 4280 98976 4296 99040
rect 4360 98976 4376 99040
rect 4440 98976 4456 99040
rect 4520 98976 4528 99040
rect 4208 97952 4528 98976
rect 4208 97888 4216 97952
rect 4280 97888 4296 97952
rect 4360 97888 4376 97952
rect 4440 97888 4456 97952
rect 4520 97888 4528 97952
rect 4208 96864 4528 97888
rect 4208 96800 4216 96864
rect 4280 96800 4296 96864
rect 4360 96800 4376 96864
rect 4440 96800 4456 96864
rect 4520 96800 4528 96864
rect 4208 95776 4528 96800
rect 4208 95712 4216 95776
rect 4280 95712 4296 95776
rect 4360 95712 4376 95776
rect 4440 95712 4456 95776
rect 4520 95712 4528 95776
rect 4208 94688 4528 95712
rect 4208 94624 4216 94688
rect 4280 94624 4296 94688
rect 4360 94624 4376 94688
rect 4440 94624 4456 94688
rect 4520 94624 4528 94688
rect 4208 93600 4528 94624
rect 4208 93536 4216 93600
rect 4280 93536 4296 93600
rect 4360 93536 4376 93600
rect 4440 93536 4456 93600
rect 4520 93536 4528 93600
rect 4208 92512 4528 93536
rect 4208 92448 4216 92512
rect 4280 92448 4296 92512
rect 4360 92448 4376 92512
rect 4440 92448 4456 92512
rect 4520 92448 4528 92512
rect 4208 91424 4528 92448
rect 4208 91360 4216 91424
rect 4280 91360 4296 91424
rect 4360 91360 4376 91424
rect 4440 91360 4456 91424
rect 4520 91360 4528 91424
rect 4208 90336 4528 91360
rect 4208 90272 4216 90336
rect 4280 90272 4296 90336
rect 4360 90272 4376 90336
rect 4440 90272 4456 90336
rect 4520 90272 4528 90336
rect 4208 89248 4528 90272
rect 4208 89184 4216 89248
rect 4280 89184 4296 89248
rect 4360 89184 4376 89248
rect 4440 89184 4456 89248
rect 4520 89184 4528 89248
rect 4208 88160 4528 89184
rect 4208 88096 4216 88160
rect 4280 88096 4296 88160
rect 4360 88096 4376 88160
rect 4440 88096 4456 88160
rect 4520 88096 4528 88160
rect 4208 87072 4528 88096
rect 4208 87008 4216 87072
rect 4280 87008 4296 87072
rect 4360 87008 4376 87072
rect 4440 87008 4456 87072
rect 4520 87008 4528 87072
rect 4208 85984 4528 87008
rect 4208 85920 4216 85984
rect 4280 85920 4296 85984
rect 4360 85920 4376 85984
rect 4440 85920 4456 85984
rect 4520 85920 4528 85984
rect 4208 84896 4528 85920
rect 4208 84832 4216 84896
rect 4280 84832 4296 84896
rect 4360 84832 4376 84896
rect 4440 84832 4456 84896
rect 4520 84832 4528 84896
rect 4208 83808 4528 84832
rect 4208 83744 4216 83808
rect 4280 83744 4296 83808
rect 4360 83744 4376 83808
rect 4440 83744 4456 83808
rect 4520 83744 4528 83808
rect 4208 82720 4528 83744
rect 4208 82656 4216 82720
rect 4280 82656 4296 82720
rect 4360 82656 4376 82720
rect 4440 82656 4456 82720
rect 4520 82656 4528 82720
rect 4208 81632 4528 82656
rect 4208 81568 4216 81632
rect 4280 81568 4296 81632
rect 4360 81568 4376 81632
rect 4440 81568 4456 81632
rect 4520 81568 4528 81632
rect 4208 80544 4528 81568
rect 4208 80480 4216 80544
rect 4280 80480 4296 80544
rect 4360 80480 4376 80544
rect 4440 80480 4456 80544
rect 4520 80480 4528 80544
rect 4208 79456 4528 80480
rect 4208 79392 4216 79456
rect 4280 79392 4296 79456
rect 4360 79392 4376 79456
rect 4440 79392 4456 79456
rect 4520 79392 4528 79456
rect 4208 78368 4528 79392
rect 4208 78304 4216 78368
rect 4280 78304 4296 78368
rect 4360 78304 4376 78368
rect 4440 78304 4456 78368
rect 4520 78304 4528 78368
rect 4208 77280 4528 78304
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66400 4528 67424
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 116992 19888 117552
rect 19568 116928 19576 116992
rect 19640 116928 19656 116992
rect 19720 116928 19736 116992
rect 19800 116928 19816 116992
rect 19880 116928 19888 116992
rect 19568 115904 19888 116928
rect 19568 115840 19576 115904
rect 19640 115840 19656 115904
rect 19720 115840 19736 115904
rect 19800 115840 19816 115904
rect 19880 115840 19888 115904
rect 19568 114816 19888 115840
rect 19568 114752 19576 114816
rect 19640 114752 19656 114816
rect 19720 114752 19736 114816
rect 19800 114752 19816 114816
rect 19880 114752 19888 114816
rect 19568 113728 19888 114752
rect 19568 113664 19576 113728
rect 19640 113664 19656 113728
rect 19720 113664 19736 113728
rect 19800 113664 19816 113728
rect 19880 113664 19888 113728
rect 19568 112640 19888 113664
rect 19568 112576 19576 112640
rect 19640 112576 19656 112640
rect 19720 112576 19736 112640
rect 19800 112576 19816 112640
rect 19880 112576 19888 112640
rect 19568 111552 19888 112576
rect 19568 111488 19576 111552
rect 19640 111488 19656 111552
rect 19720 111488 19736 111552
rect 19800 111488 19816 111552
rect 19880 111488 19888 111552
rect 19568 110464 19888 111488
rect 19568 110400 19576 110464
rect 19640 110400 19656 110464
rect 19720 110400 19736 110464
rect 19800 110400 19816 110464
rect 19880 110400 19888 110464
rect 19568 109376 19888 110400
rect 19568 109312 19576 109376
rect 19640 109312 19656 109376
rect 19720 109312 19736 109376
rect 19800 109312 19816 109376
rect 19880 109312 19888 109376
rect 19568 108288 19888 109312
rect 19568 108224 19576 108288
rect 19640 108224 19656 108288
rect 19720 108224 19736 108288
rect 19800 108224 19816 108288
rect 19880 108224 19888 108288
rect 19568 107200 19888 108224
rect 19568 107136 19576 107200
rect 19640 107136 19656 107200
rect 19720 107136 19736 107200
rect 19800 107136 19816 107200
rect 19880 107136 19888 107200
rect 19568 106112 19888 107136
rect 19568 106048 19576 106112
rect 19640 106048 19656 106112
rect 19720 106048 19736 106112
rect 19800 106048 19816 106112
rect 19880 106048 19888 106112
rect 19568 105024 19888 106048
rect 19568 104960 19576 105024
rect 19640 104960 19656 105024
rect 19720 104960 19736 105024
rect 19800 104960 19816 105024
rect 19880 104960 19888 105024
rect 19568 103936 19888 104960
rect 19568 103872 19576 103936
rect 19640 103872 19656 103936
rect 19720 103872 19736 103936
rect 19800 103872 19816 103936
rect 19880 103872 19888 103936
rect 19568 102848 19888 103872
rect 19568 102784 19576 102848
rect 19640 102784 19656 102848
rect 19720 102784 19736 102848
rect 19800 102784 19816 102848
rect 19880 102784 19888 102848
rect 19568 101760 19888 102784
rect 19568 101696 19576 101760
rect 19640 101696 19656 101760
rect 19720 101696 19736 101760
rect 19800 101696 19816 101760
rect 19880 101696 19888 101760
rect 19568 100672 19888 101696
rect 19568 100608 19576 100672
rect 19640 100608 19656 100672
rect 19720 100608 19736 100672
rect 19800 100608 19816 100672
rect 19880 100608 19888 100672
rect 19568 99584 19888 100608
rect 19568 99520 19576 99584
rect 19640 99520 19656 99584
rect 19720 99520 19736 99584
rect 19800 99520 19816 99584
rect 19880 99520 19888 99584
rect 19568 98496 19888 99520
rect 19568 98432 19576 98496
rect 19640 98432 19656 98496
rect 19720 98432 19736 98496
rect 19800 98432 19816 98496
rect 19880 98432 19888 98496
rect 19568 97408 19888 98432
rect 19568 97344 19576 97408
rect 19640 97344 19656 97408
rect 19720 97344 19736 97408
rect 19800 97344 19816 97408
rect 19880 97344 19888 97408
rect 19568 96320 19888 97344
rect 19568 96256 19576 96320
rect 19640 96256 19656 96320
rect 19720 96256 19736 96320
rect 19800 96256 19816 96320
rect 19880 96256 19888 96320
rect 19568 95232 19888 96256
rect 19568 95168 19576 95232
rect 19640 95168 19656 95232
rect 19720 95168 19736 95232
rect 19800 95168 19816 95232
rect 19880 95168 19888 95232
rect 19568 94144 19888 95168
rect 19568 94080 19576 94144
rect 19640 94080 19656 94144
rect 19720 94080 19736 94144
rect 19800 94080 19816 94144
rect 19880 94080 19888 94144
rect 19568 93056 19888 94080
rect 19568 92992 19576 93056
rect 19640 92992 19656 93056
rect 19720 92992 19736 93056
rect 19800 92992 19816 93056
rect 19880 92992 19888 93056
rect 19568 91968 19888 92992
rect 19568 91904 19576 91968
rect 19640 91904 19656 91968
rect 19720 91904 19736 91968
rect 19800 91904 19816 91968
rect 19880 91904 19888 91968
rect 19568 90880 19888 91904
rect 19568 90816 19576 90880
rect 19640 90816 19656 90880
rect 19720 90816 19736 90880
rect 19800 90816 19816 90880
rect 19880 90816 19888 90880
rect 19568 89792 19888 90816
rect 19568 89728 19576 89792
rect 19640 89728 19656 89792
rect 19720 89728 19736 89792
rect 19800 89728 19816 89792
rect 19880 89728 19888 89792
rect 19568 88704 19888 89728
rect 19568 88640 19576 88704
rect 19640 88640 19656 88704
rect 19720 88640 19736 88704
rect 19800 88640 19816 88704
rect 19880 88640 19888 88704
rect 19568 87616 19888 88640
rect 19568 87552 19576 87616
rect 19640 87552 19656 87616
rect 19720 87552 19736 87616
rect 19800 87552 19816 87616
rect 19880 87552 19888 87616
rect 19568 86528 19888 87552
rect 19568 86464 19576 86528
rect 19640 86464 19656 86528
rect 19720 86464 19736 86528
rect 19800 86464 19816 86528
rect 19880 86464 19888 86528
rect 19568 85440 19888 86464
rect 19568 85376 19576 85440
rect 19640 85376 19656 85440
rect 19720 85376 19736 85440
rect 19800 85376 19816 85440
rect 19880 85376 19888 85440
rect 19568 84352 19888 85376
rect 19568 84288 19576 84352
rect 19640 84288 19656 84352
rect 19720 84288 19736 84352
rect 19800 84288 19816 84352
rect 19880 84288 19888 84352
rect 19568 83264 19888 84288
rect 19568 83200 19576 83264
rect 19640 83200 19656 83264
rect 19720 83200 19736 83264
rect 19800 83200 19816 83264
rect 19880 83200 19888 83264
rect 19568 82176 19888 83200
rect 19568 82112 19576 82176
rect 19640 82112 19656 82176
rect 19720 82112 19736 82176
rect 19800 82112 19816 82176
rect 19880 82112 19888 82176
rect 19568 81088 19888 82112
rect 19568 81024 19576 81088
rect 19640 81024 19656 81088
rect 19720 81024 19736 81088
rect 19800 81024 19816 81088
rect 19880 81024 19888 81088
rect 19568 80000 19888 81024
rect 19568 79936 19576 80000
rect 19640 79936 19656 80000
rect 19720 79936 19736 80000
rect 19800 79936 19816 80000
rect 19880 79936 19888 80000
rect 19568 78912 19888 79936
rect 19568 78848 19576 78912
rect 19640 78848 19656 78912
rect 19720 78848 19736 78912
rect 19800 78848 19816 78912
rect 19880 78848 19888 78912
rect 19568 77824 19888 78848
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 76736 19888 77760
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 75648 19888 76672
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 74560 19888 75584
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 73472 19888 74496
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 72384 19888 73408
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 71296 19888 72320
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 70208 19888 71232
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 69120 19888 70144
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 68032 19888 69056
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 66944 19888 67968
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 65856 19888 66880
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 64768 19888 65792
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 63680 19888 64704
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 62592 19888 63616
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 61504 19888 62528
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 60416 19888 61440
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 59328 19888 60352
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 58240 19888 59264
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 57152 19888 58176
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 117536 35248 117552
rect 34928 117472 34936 117536
rect 35000 117472 35016 117536
rect 35080 117472 35096 117536
rect 35160 117472 35176 117536
rect 35240 117472 35248 117536
rect 34928 116448 35248 117472
rect 34928 116384 34936 116448
rect 35000 116384 35016 116448
rect 35080 116384 35096 116448
rect 35160 116384 35176 116448
rect 35240 116384 35248 116448
rect 34928 115360 35248 116384
rect 34928 115296 34936 115360
rect 35000 115296 35016 115360
rect 35080 115296 35096 115360
rect 35160 115296 35176 115360
rect 35240 115296 35248 115360
rect 34928 114272 35248 115296
rect 34928 114208 34936 114272
rect 35000 114208 35016 114272
rect 35080 114208 35096 114272
rect 35160 114208 35176 114272
rect 35240 114208 35248 114272
rect 34928 113184 35248 114208
rect 34928 113120 34936 113184
rect 35000 113120 35016 113184
rect 35080 113120 35096 113184
rect 35160 113120 35176 113184
rect 35240 113120 35248 113184
rect 34928 112096 35248 113120
rect 34928 112032 34936 112096
rect 35000 112032 35016 112096
rect 35080 112032 35096 112096
rect 35160 112032 35176 112096
rect 35240 112032 35248 112096
rect 34928 111008 35248 112032
rect 34928 110944 34936 111008
rect 35000 110944 35016 111008
rect 35080 110944 35096 111008
rect 35160 110944 35176 111008
rect 35240 110944 35248 111008
rect 34928 109920 35248 110944
rect 34928 109856 34936 109920
rect 35000 109856 35016 109920
rect 35080 109856 35096 109920
rect 35160 109856 35176 109920
rect 35240 109856 35248 109920
rect 34928 108832 35248 109856
rect 34928 108768 34936 108832
rect 35000 108768 35016 108832
rect 35080 108768 35096 108832
rect 35160 108768 35176 108832
rect 35240 108768 35248 108832
rect 34928 107744 35248 108768
rect 34928 107680 34936 107744
rect 35000 107680 35016 107744
rect 35080 107680 35096 107744
rect 35160 107680 35176 107744
rect 35240 107680 35248 107744
rect 34928 106656 35248 107680
rect 34928 106592 34936 106656
rect 35000 106592 35016 106656
rect 35080 106592 35096 106656
rect 35160 106592 35176 106656
rect 35240 106592 35248 106656
rect 34928 105568 35248 106592
rect 34928 105504 34936 105568
rect 35000 105504 35016 105568
rect 35080 105504 35096 105568
rect 35160 105504 35176 105568
rect 35240 105504 35248 105568
rect 34928 104480 35248 105504
rect 34928 104416 34936 104480
rect 35000 104416 35016 104480
rect 35080 104416 35096 104480
rect 35160 104416 35176 104480
rect 35240 104416 35248 104480
rect 34928 103392 35248 104416
rect 34928 103328 34936 103392
rect 35000 103328 35016 103392
rect 35080 103328 35096 103392
rect 35160 103328 35176 103392
rect 35240 103328 35248 103392
rect 34928 102304 35248 103328
rect 34928 102240 34936 102304
rect 35000 102240 35016 102304
rect 35080 102240 35096 102304
rect 35160 102240 35176 102304
rect 35240 102240 35248 102304
rect 34928 101216 35248 102240
rect 34928 101152 34936 101216
rect 35000 101152 35016 101216
rect 35080 101152 35096 101216
rect 35160 101152 35176 101216
rect 35240 101152 35248 101216
rect 34928 100128 35248 101152
rect 34928 100064 34936 100128
rect 35000 100064 35016 100128
rect 35080 100064 35096 100128
rect 35160 100064 35176 100128
rect 35240 100064 35248 100128
rect 34928 99040 35248 100064
rect 34928 98976 34936 99040
rect 35000 98976 35016 99040
rect 35080 98976 35096 99040
rect 35160 98976 35176 99040
rect 35240 98976 35248 99040
rect 34928 97952 35248 98976
rect 34928 97888 34936 97952
rect 35000 97888 35016 97952
rect 35080 97888 35096 97952
rect 35160 97888 35176 97952
rect 35240 97888 35248 97952
rect 34928 96864 35248 97888
rect 34928 96800 34936 96864
rect 35000 96800 35016 96864
rect 35080 96800 35096 96864
rect 35160 96800 35176 96864
rect 35240 96800 35248 96864
rect 34928 95776 35248 96800
rect 34928 95712 34936 95776
rect 35000 95712 35016 95776
rect 35080 95712 35096 95776
rect 35160 95712 35176 95776
rect 35240 95712 35248 95776
rect 34928 94688 35248 95712
rect 34928 94624 34936 94688
rect 35000 94624 35016 94688
rect 35080 94624 35096 94688
rect 35160 94624 35176 94688
rect 35240 94624 35248 94688
rect 34928 93600 35248 94624
rect 34928 93536 34936 93600
rect 35000 93536 35016 93600
rect 35080 93536 35096 93600
rect 35160 93536 35176 93600
rect 35240 93536 35248 93600
rect 34928 92512 35248 93536
rect 34928 92448 34936 92512
rect 35000 92448 35016 92512
rect 35080 92448 35096 92512
rect 35160 92448 35176 92512
rect 35240 92448 35248 92512
rect 34928 91424 35248 92448
rect 34928 91360 34936 91424
rect 35000 91360 35016 91424
rect 35080 91360 35096 91424
rect 35160 91360 35176 91424
rect 35240 91360 35248 91424
rect 34928 90336 35248 91360
rect 34928 90272 34936 90336
rect 35000 90272 35016 90336
rect 35080 90272 35096 90336
rect 35160 90272 35176 90336
rect 35240 90272 35248 90336
rect 34928 89248 35248 90272
rect 34928 89184 34936 89248
rect 35000 89184 35016 89248
rect 35080 89184 35096 89248
rect 35160 89184 35176 89248
rect 35240 89184 35248 89248
rect 34928 88160 35248 89184
rect 34928 88096 34936 88160
rect 35000 88096 35016 88160
rect 35080 88096 35096 88160
rect 35160 88096 35176 88160
rect 35240 88096 35248 88160
rect 34928 87072 35248 88096
rect 34928 87008 34936 87072
rect 35000 87008 35016 87072
rect 35080 87008 35096 87072
rect 35160 87008 35176 87072
rect 35240 87008 35248 87072
rect 34928 85984 35248 87008
rect 34928 85920 34936 85984
rect 35000 85920 35016 85984
rect 35080 85920 35096 85984
rect 35160 85920 35176 85984
rect 35240 85920 35248 85984
rect 34928 84896 35248 85920
rect 34928 84832 34936 84896
rect 35000 84832 35016 84896
rect 35080 84832 35096 84896
rect 35160 84832 35176 84896
rect 35240 84832 35248 84896
rect 34928 83808 35248 84832
rect 34928 83744 34936 83808
rect 35000 83744 35016 83808
rect 35080 83744 35096 83808
rect 35160 83744 35176 83808
rect 35240 83744 35248 83808
rect 34928 82720 35248 83744
rect 34928 82656 34936 82720
rect 35000 82656 35016 82720
rect 35080 82656 35096 82720
rect 35160 82656 35176 82720
rect 35240 82656 35248 82720
rect 34928 81632 35248 82656
rect 34928 81568 34936 81632
rect 35000 81568 35016 81632
rect 35080 81568 35096 81632
rect 35160 81568 35176 81632
rect 35240 81568 35248 81632
rect 34928 80544 35248 81568
rect 34928 80480 34936 80544
rect 35000 80480 35016 80544
rect 35080 80480 35096 80544
rect 35160 80480 35176 80544
rect 35240 80480 35248 80544
rect 34928 79456 35248 80480
rect 34928 79392 34936 79456
rect 35000 79392 35016 79456
rect 35080 79392 35096 79456
rect 35160 79392 35176 79456
rect 35240 79392 35248 79456
rect 34928 78368 35248 79392
rect 34928 78304 34936 78368
rect 35000 78304 35016 78368
rect 35080 78304 35096 78368
rect 35160 78304 35176 78368
rect 35240 78304 35248 78368
rect 34928 77280 35248 78304
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 76192 35248 77216
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 75104 35248 76128
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 74016 35248 75040
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 72928 35248 73952
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 71840 35248 72864
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 70752 35248 71776
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 69664 35248 70688
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 68576 35248 69600
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 67488 35248 68512
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 66400 35248 67424
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 65312 35248 66336
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 64224 35248 65248
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 63136 35248 64160
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 62048 35248 63072
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 60960 35248 61984
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 59872 35248 60896
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 58784 35248 59808
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 57696 35248 58720
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input475 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input331 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623621585
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2116 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12
timestamp 1623621585
transform 1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input509 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2852 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input476
timestamp 1623621585
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_25
timestamp 1623621585
transform 1 0 3404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1623621585
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1623621585
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input520 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 4232 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input487
timestamp 1623621585
transform 1 0 4232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1623621585
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1623621585
transform 1 0 4600 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1623621585
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1623621585
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1623621585
transform 1 0 5520 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output739
timestamp 1623621585
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output728
timestamp 1623621585
transform 1 0 4968 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output631
timestamp 1623621585
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_54
timestamp 1623621585
transform 1 0 6072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1623621585
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  input534
timestamp 1623621585
transform 1 0 6440 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1623621585
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1623621585
transform 1 0 7544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_64
timestamp 1623621585
transform 1 0 6992 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1623621585
transform 1 0 7452 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input535
timestamp 1623621585
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input501
timestamp 1623621585
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1623621585
transform 1 0 8004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1623621585
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input504
timestamp 1623621585
transform 1 0 8372 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input503 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 8372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1623621585
transform 1 0 8648 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1623621585
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1623621585
transform 1 0 9108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88
timestamp 1623621585
transform 1 0 9200 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output743
timestamp 1623621585
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1623621585
transform 1 0 9016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1623621585
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1623621585
transform 1 0 9844 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input537
timestamp 1623621585
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input505
timestamp 1623621585
transform 1 0 9936 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1623621585
transform 1 0 10488 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1623621585
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1623621585
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input477
timestamp 1623621585
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input506
timestamp 1623621585
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input507
timestamp 1623621585
transform 1 0 11776 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input538
timestamp 1623621585
transform 1 0 10856 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1623621585
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1623621585
transform 1 0 11868 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_110
timestamp 1623621585
transform 1 0 11224 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_122
timestamp 1623621585
transform 1 0 12328 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1623621585
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1623621585
transform 1 0 14260 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input478
timestamp 1623621585
transform 1 0 13524 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input510
timestamp 1623621585
transform 1 0 12880 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1623621585
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1623621585
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134
timestamp 1623621585
transform 1 0 13432 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1623621585
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1623621585
transform 1 0 14352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1623621585
transform 1 0 15088 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1623621585
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output718
timestamp 1623621585
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input479
timestamp 1623621585
transform 1 0 14904 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1623621585
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1623621585
transform 1 0 15456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1623621585
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input513
timestamp 1623621585
transform 1 0 15548 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input480
timestamp 1623621585
transform 1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_166
timestamp 1623621585
transform 1 0 16376 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0820_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17296 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1623621585
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input482
timestamp 1623621585
transform 1 0 16560 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input515
timestamp 1623621585
transform 1 0 17572 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1623621585
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185
timestamp 1623621585
transform 1 0 18124 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1623621585
transform 1 0 16468 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1623621585
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1623621585
transform 1 0 18124 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_193
timestamp 1623621585
transform 1 0 18860 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input517
timestamp 1623621585
transform 1 0 18860 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input516
timestamp 1623621585
transform 1 0 18492 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_201
timestamp 1623621585
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1623621585
transform 1 0 19412 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1623621585
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1623621585
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1623621585
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output725
timestamp 1623621585
transform 1 0 19964 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input518
timestamp 1623621585
transform 1 0 20240 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1623621585
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_213
timestamp 1623621585
transform 1 0 20700 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp 1623621585
transform 1 0 20332 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_212
timestamp 1623621585
transform 1 0 20608 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input519
timestamp 1623621585
transform 1 0 20792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_226
timestamp 1623621585
transform 1 0 21896 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1623621585
transform 1 0 21160 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_220
timestamp 1623621585
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output727
timestamp 1623621585
transform 1 0 21528 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input521
timestamp 1623621585
transform 1 0 21528 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1623621585
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0823_
timestamp 1623621585
transform 1 0 23368 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1623621585
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input523
timestamp 1623621585
transform 1 0 23460 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output729
timestamp 1623621585
transform 1 0 22264 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_233
timestamp 1623621585
transform 1 0 22540 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_241
timestamp 1623621585
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1623621585
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_234
timestamp 1623621585
transform 1 0 22632 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_251
timestamp 1623621585
transform 1 0 24196 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output726
timestamp 1623621585
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1623621585
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1623621585
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1623621585
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output732
timestamp 1623621585
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1623621585
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1623621585
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_266
timestamp 1623621585
transform 1 0 25576 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input524
timestamp 1623621585
transform 1 0 25576 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0822_
timestamp 1623621585
transform 1 0 26128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1623621585
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input527 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 26864 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output734
timestamp 1623621585
transform 1 0 27324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1623621585
transform 1 0 26128 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1623621585
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1623621585
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1623621585
transform 1 0 26956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1623621585
transform 1 0 27692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input528
timestamp 1623621585
transform 1 0 28244 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input529
timestamp 1623621585
transform 1 0 29164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input530
timestamp 1623621585
transform 1 0 29256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output735
timestamp 1623621585
transform 1 0 28060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_301
timestamp 1623621585
transform 1 0 28796 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_309
timestamp 1623621585
transform 1 0 29532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_297
timestamp 1623621585
transform 1 0 28428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_305
timestamp 1623621585
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1623621585
transform 1 0 29624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_315
timestamp 1623621585
transform 1 0 30084 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_317
timestamp 1623621585
transform 1 0 30268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1623621585
transform 1 0 29992 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1623621585
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_326
timestamp 1623621585
transform 1 0 31096 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_321
timestamp 1623621585
transform 1 0 30636 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1623621585
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output696
timestamp 1623621585
transform 1 0 30728 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input532
timestamp 1623621585
transform 1 0 30912 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_330
timestamp 1623621585
transform 1 0 31464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output669
timestamp 1623621585
transform 1 0 31464 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_342
timestamp 1623621585
transform 1 0 32568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_334
timestamp 1623621585
transform 1 0 31832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_339
timestamp 1623621585
transform 1 0 32292 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_334
timestamp 1623621585
transform 1 0 31832 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1623621585
transform 1 0 32200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1623621585
transform 1 0 31924 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1623621585
transform 1 0 33304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1623621585
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_347
timestamp 1623621585
transform 1 0 33028 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1623621585
transform 1 0 32936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1623621585
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1623621585
transform 1 0 33672 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1623621585
transform 1 0 33580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_358
timestamp 1623621585
transform 1 0 34040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_357
timestamp 1623621585
transform 1 0 33948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1623621585
transform 1 0 34408 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_370
timestamp 1623621585
transform 1 0 35144 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_366
timestamp 1623621585
transform 1 0 34776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_365
timestamp 1623621585
transform 1 0 34684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input40
timestamp 1623621585
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1623621585
transform 1 0 35236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1623621585
transform 1 0 35328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_372
timestamp 1623621585
transform 1 0 35328 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1623621585
transform 1 0 36248 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_378
timestamp 1623621585
transform 1 0 35880 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_376
timestamp 1623621585
transform 1 0 35696 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input41
timestamp 1623621585
transform 1 0 35696 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1623621585
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_390
timestamp 1623621585
transform 1 0 36984 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_391
timestamp 1623621585
transform 1 0 37076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_384
timestamp 1623621585
transform 1 0 36432 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1623621585
transform 1 0 37076 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input69
timestamp 1623621585
transform 1 0 36524 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_395
timestamp 1623621585
transform 1 0 37444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623621585
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623621585
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1623621585
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1623621585
transform 1 0 37720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1623621585
transform 1 0 37812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_397
timestamp 1623621585
transform 1 0 37628 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1623621585
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1623621585
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623621585
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input342
timestamp 1623621585
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input353
timestamp 1623621585
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1623621585
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1623621585
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_19
timestamp 1623621585
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input546
timestamp 1623621585
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output717
timestamp 1623621585
transform 1 0 3956 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1623621585
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_35
timestamp 1623621585
transform 1 0 4324 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1623621585
transform 1 0 4876 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1623621585
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input498
timestamp 1623621585
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input531
timestamp 1623621585
transform 1 0 5612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output742
timestamp 1623621585
transform 1 0 6808 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1623621585
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1623621585
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1623621585
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1623621585
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input502
timestamp 1623621585
transform 1 0 7544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input536
timestamp 1623621585
transform 1 0 8556 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1623621585
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1623621585
transform 1 0 7820 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output744
timestamp 1623621585
transform 1 0 9292 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output745
timestamp 1623621585
transform 1 0 10028 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1623621585
transform 1 0 8924 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_93
timestamp 1623621585
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1623621585
transform 1 0 10396 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1623621585
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input539
timestamp 1623621585
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input540
timestamp 1623621585
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_105
timestamp 1623621585
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_110
timestamp 1623621585
transform 1 0 11224 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1623621585
transform 1 0 11684 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_123
timestamp 1623621585
transform 1 0 12420 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input511
timestamp 1623621585
transform 1 0 13800 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output748
timestamp 1623621585
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_131
timestamp 1623621585
transform 1 0 13156 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_137
timestamp 1623621585
transform 1 0 13708 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1623621585
transform 1 0 14352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input481
timestamp 1623621585
transform 1 0 15456 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input514
timestamp 1623621585
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output719
timestamp 1623621585
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_152
timestamp 1623621585
transform 1 0 15088 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1623621585
transform 1 0 15732 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1623621585
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output722
timestamp 1623621585
transform 1 0 17296 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output723
timestamp 1623621585
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1623621585
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1623621585
transform 1 0 16928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1623621585
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input484 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output724
timestamp 1623621585
transform 1 0 18768 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_188
timestamp 1623621585
transform 1 0 18400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_196
timestamp 1623621585
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_203
timestamp 1623621585
transform 1 0 19780 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0918_
timestamp 1623621585
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0930_
timestamp 1623621585
transform 1 0 20976 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1623621585
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_212
timestamp 1623621585
transform 1 0 20608 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_219
timestamp 1623621585
transform 1 0 21252 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_227
timestamp 1623621585
transform 1 0 21988 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_229
timestamp 1623621585
transform 1 0 22172 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output730
timestamp 1623621585
transform 1 0 22816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output731
timestamp 1623621585
transform 1 0 23736 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_235
timestamp 1623621585
transform 1 0 22724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_240
timestamp 1623621585
transform 1 0 23184 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_250
timestamp 1623621585
transform 1 0 24104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input491
timestamp 1623621585
transform 1 0 24472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output733
timestamp 1623621585
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_257
timestamp 1623621585
transform 1 0 24748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_267
timestamp 1623621585
transform 1 0 25668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1623621585
transform 1 0 27324 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input526
timestamp 1623621585
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_275
timestamp 1623621585
transform 1 0 26404 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_283
timestamp 1623621585
transform 1 0 27140 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_286
timestamp 1623621585
transform 1 0 27416 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _0826_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 29532 0 -1 3808
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  output736
timestamp 1623621585
transform 1 0 28060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output737
timestamp 1623621585
transform 1 0 28796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_292
timestamp 1623621585
transform 1 0 27968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_297
timestamp 1623621585
transform 1 0 28428 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_305
timestamp 1623621585
transform 1 0 29164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output738
timestamp 1623621585
transform 1 0 30912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_320
timestamp 1623621585
transform 1 0 30544 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_328
timestamp 1623621585
transform 1 0 31280 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1623621585
transform 1 0 32568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1623621585
transform 1 0 33304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output694
timestamp 1623621585
transform 1 0 31832 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_338
timestamp 1623621585
transform 1 0 32200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_343
timestamp 1623621585
transform 1 0 32660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_349
timestamp 1623621585
transform 1 0 33212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_354
timestamp 1623621585
transform 1 0 33672 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1623621585
transform 1 0 34040 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input49
timestamp 1623621585
transform 1 0 34776 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_362
timestamp 1623621585
transform 1 0 34408 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_370
timestamp 1623621585
transform 1 0 35144 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1623621585
transform 1 0 35696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1623621585
transform 1 0 37076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_380
timestamp 1623621585
transform 1 0 36064 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_388
timestamp 1623621585
transform 1 0 36800 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1623621585
transform 1 0 37444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623621585
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1623621585
transform 1 0 37812 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_400
timestamp 1623621585
transform 1 0 37904 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1623621585
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623621585
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output632
timestamp 1623621585
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output716
timestamp 1623621585
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1623621585
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_11
timestamp 1623621585
transform 1 0 2116 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp 1623621585
transform 1 0 2852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1623621585
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input508
timestamp 1623621585
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input541
timestamp 1623621585
transform 1 0 4876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1623621585
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1623621585
transform 1 0 3864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_37
timestamp 1623621585
transform 1 0 4508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input542
timestamp 1623621585
transform 1 0 5520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input543
timestamp 1623621585
transform 1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1623621585
transform 1 0 5152 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1623621585
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_58
timestamp 1623621585
transform 1 0 6440 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input544
timestamp 1623621585
transform 1 0 7084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_64
timestamp 1623621585
transform 1 0 6992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 7360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_80
timestamp 1623621585
transform 1 0 8464 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 9844 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1623621585
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_87
timestamp 1623621585
transform 1 0 9108 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1623621585
transform 1 0 10488 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output746
timestamp 1623621585
transform 1 0 10856 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output747
timestamp 1623621585
transform 1 0 11592 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1623621585
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_118
timestamp 1623621585
transform 1 0 11960 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1623621585
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_130
timestamp 1623621585
transform 1 0 13064 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_142
timestamp 1623621585
transform 1 0 14168 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_144
timestamp 1623621585
transform 1 0 14352 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output720
timestamp 1623621585
transform 1 0 14904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output721
timestamp 1623621585
transform 1 0 15824 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_154
timestamp 1623621585
transform 1 0 15272 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_164
timestamp 1623621585
transform 1 0 16192 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input483
timestamp 1623621585
transform 1 0 17848 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_176
timestamp 1623621585
transform 1 0 17296 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_185
timestamp 1623621585
transform 1 0 18124 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1623621585
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input485
timestamp 1623621585
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_197
timestamp 1623621585
transform 1 0 19228 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_201
timestamp 1623621585
transform 1 0 19596 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_208
timestamp 1623621585
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0920_
timestamp 1623621585
transform 1 0 21988 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input486
timestamp 1623621585
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input488
timestamp 1623621585
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1623621585
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1623621585
transform 1 0 21252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_223
timestamp 1623621585
transform 1 0 21620 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0921_
timestamp 1623621585
transform 1 0 22632 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0934_
timestamp 1623621585
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input490
timestamp 1623621585
transform 1 0 23920 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_230
timestamp 1623621585
transform 1 0 22264 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 1623621585
transform 1 0 22908 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1623621585
transform 1 0 23552 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1623621585
transform 1 0 24748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input492
timestamp 1623621585
transform 1 0 25208 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input493
timestamp 1623621585
transform 1 0 25852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_251
timestamp 1623621585
transform 1 0 24196 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1623621585
transform 1 0 24840 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_265
timestamp 1623621585
transform 1 0 25484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0825_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0940_
timestamp 1623621585
transform 1 0 26588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input495
timestamp 1623621585
transform 1 0 27876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1623621585
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1623621585
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_280
timestamp 1623621585
transform 1 0 26864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_287
timestamp 1623621585
transform 1 0 27508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input496
timestamp 1623621585
transform 1 0 28520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input497
timestamp 1623621585
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_294
timestamp 1623621585
transform 1 0 28152 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_301
timestamp 1623621585
transform 1 0 28796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_305
timestamp 1623621585
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_309
timestamp 1623621585
transform 1 0 29532 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1623621585
transform 1 0 29992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output740
timestamp 1623621585
transform 1 0 30728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output741
timestamp 1623621585
transform 1 0 31556 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_313
timestamp 1623621585
transform 1 0 29900 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_315
timestamp 1623621585
transform 1 0 30084 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_321
timestamp 1623621585
transform 1 0 30636 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_326
timestamp 1623621585
transform 1 0 31096 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_330
timestamp 1623621585
transform 1 0 31464 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1623621585
transform 1 0 32292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output685
timestamp 1623621585
transform 1 0 33028 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_335
timestamp 1623621585
transform 1 0 31924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_342
timestamp 1623621585
transform 1 0 32568 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_346
timestamp 1623621585
transform 1 0 32936 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_351
timestamp 1623621585
transform 1 0 33396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1623621585
transform 1 0 35236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1623621585
transform 1 0 34500 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output654
timestamp 1623621585
transform 1 0 33764 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_359
timestamp 1623621585
transform 1 0 34132 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1623621585
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_372
timestamp 1623621585
transform 1 0 35328 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1623621585
transform 1 0 35696 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1623621585
transform 1 0 37076 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1623621585
transform 1 0 36340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_379
timestamp 1623621585
transform 1 0 35972 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1623621585
transform 1 0 36708 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1623621585
transform 1 0 37444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623621585
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1623621585
transform 1 0 37812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1623621585
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 2484 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623621585
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output633
timestamp 1623621585
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1623621585
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1623621585
transform 1 0 2116 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_18
timestamp 1623621585
transform 1 0 2760 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0898_
timestamp 1623621585
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_25
timestamp 1623621585
transform 1 0 3404 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_37
timestamp 1623621585
transform 1 0 4508 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1623621585
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_49
timestamp 1623621585
transform 1 0 5612 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_58
timestamp 1623621585
transform 1 0 6440 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1623621585
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_82
timestamp 1623621585
transform 1 0 8648 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_94
timestamp 1623621585
transform 1 0 9752 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1623621585
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_106
timestamp 1623621585
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1623621585
transform 1 0 11684 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1623621585
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_139
timestamp 1623621585
transform 1 0 13892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input512
timestamp 1623621585
transform 1 0 14628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_150
timestamp 1623621585
transform 1 0 14904 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_162
timestamp 1623621585
transform 1 0 16008 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1623621585
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_170
timestamp 1623621585
transform 1 0 16744 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_172
timestamp 1623621585
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1623621585
transform 1 0 18032 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1623621585
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_208
timestamp 1623621585
transform 1 0 20240 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1623621585
transform 1 0 22080 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_220
timestamp 1623621585
transform 1 0 21344 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_229
timestamp 1623621585
transform 1 0 22172 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input489
timestamp 1623621585
transform 1 0 22540 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input522
timestamp 1623621585
transform 1 0 23184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1623621585
transform 1 0 22816 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_243
timestamp 1623621585
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input525
timestamp 1623621585
transform 1 0 25208 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_255
timestamp 1623621585
transform 1 0 24564 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_261
timestamp 1623621585
transform 1 0 25116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1623621585
transform 1 0 25484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1623621585
transform 1 0 27324 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input494
timestamp 1623621585
transform 1 0 26588 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_280
timestamp 1623621585
transform 1 0 26864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_284
timestamp 1623621585
transform 1 0 27232 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_286
timestamp 1623621585
transform 1 0 27416 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_298
timestamp 1623621585
transform 1 0 28520 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_310
timestamp 1623621585
transform 1 0 29624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1623621585
transform 1 0 30728 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input499
timestamp 1623621585
transform 1 0 30084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input500
timestamp 1623621585
transform 1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_314
timestamp 1623621585
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_318
timestamp 1623621585
transform 1 0 30360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_325
timestamp 1623621585
transform 1 0 31004 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_332
timestamp 1623621585
transform 1 0 31648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1623621585
transform 1 0 32568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output688
timestamp 1623621585
transform 1 0 33396 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_340
timestamp 1623621585
transform 1 0 32384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_343
timestamp 1623621585
transform 1 0 32660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1623621585
transform 1 0 35604 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output646
timestamp 1623621585
transform 1 0 34868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output662
timestamp 1623621585
transform 1 0 34132 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_355
timestamp 1623621585
transform 1 0 33764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_363
timestamp 1623621585
transform 1 0 34500 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_371
timestamp 1623621585
transform 1 0 35236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1623621585
transform 1 0 37076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1623621585
transform 1 0 36340 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_379
timestamp 1623621585
transform 1 0 35972 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_387
timestamp 1623621585
transform 1 0 36708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1623621585
transform 1 0 37444 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623621585
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1623621585
transform 1 0 37812 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_400
timestamp 1623621585
transform 1 0 37904 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1623621585
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623621585
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input356
timestamp 1623621585
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input357
timestamp 1623621585
transform 1 0 2760 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input359
timestamp 1623621585
transform 1 0 2024 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1623621585
transform 1 0 1656 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1623621585
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_17
timestamp 1623621585
transform 1 0 2668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1623621585
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_21
timestamp 1623621585
transform 1 0 3036 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1623621585
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1623621585
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_54
timestamp 1623621585
transform 1 0 6072 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1623621585
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1623621585
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1623621585
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_87
timestamp 1623621585
transform 1 0 9108 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_99
timestamp 1623621585
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_111
timestamp 1623621585
transform 1 0 11316 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1623621585
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1623621585
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1623621585
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1623621585
transform 1 0 14352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1623621585
transform 1 0 15456 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_168
timestamp 1623621585
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_180
timestamp 1623621585
transform 1 0 17664 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1623621585
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_192
timestamp 1623621585
transform 1 0 18768 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_201
timestamp 1623621585
transform 1 0 19596 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_213
timestamp 1623621585
transform 1 0 20700 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1623621585
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1623621585
transform 1 0 22908 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_249
timestamp 1623621585
transform 1 0 24012 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1623621585
transform 1 0 24748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_258
timestamp 1623621585
transform 1 0 24840 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_270
timestamp 1623621585
transform 1 0 25944 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_282
timestamp 1623621585
transform 1 0 27048 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_294
timestamp 1623621585
transform 1 0 28152 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_306
timestamp 1623621585
transform 1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1623621585
transform 1 0 29992 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input533
timestamp 1623621585
transform 1 0 31280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_315
timestamp 1623621585
transform 1 0 30084 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_327
timestamp 1623621585
transform 1 0 31188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_331
timestamp 1623621585
transform 1 0 31556 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1623621585
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1623621585
transform 1 0 35236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output675
timestamp 1623621585
transform 1 0 34500 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output700
timestamp 1623621585
transform 1 0 33764 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_359
timestamp 1623621585
transform 1 0 34132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1623621585
transform 1 0 34868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_372
timestamp 1623621585
transform 1 0 35328 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1623621585
transform 1 0 37076 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1623621585
transform 1 0 36340 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_380
timestamp 1623621585
transform 1 0 36064 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_387
timestamp 1623621585
transform 1 0 36708 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1623621585
transform 1 0 37444 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623621585
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1623621585
transform 1 0 37812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1623621585
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_6
timestamp 1623621585
transform 1 0 1656 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input360
timestamp 1623621585
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input358
timestamp 1623621585
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623621585
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623621585
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_18
timestamp 1623621585
transform 1 0 2760 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_14
timestamp 1623621585
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input545
timestamp 1623621585
transform 1 0 2668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_6
timestamp 1623621585
transform 1 0 1656 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_20
timestamp 1623621585
transform 1 0 2944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1623621585
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1623621585
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_26
timestamp 1623621585
transform 1 0 3496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1623621585
transform 1 0 3864 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1623621585
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1623621585
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1623621585
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1623621585
transform 1 0 6440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_42
timestamp 1623621585
transform 1 0 4968 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_54
timestamp 1623621585
transform 1 0 6072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1623621585
transform 1 0 7544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_82
timestamp 1623621585
transform 1 0 8648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_66
timestamp 1623621585
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1623621585
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1623621585
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_94
timestamp 1623621585
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_87
timestamp 1623621585
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_99
timestamp 1623621585
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1623621585
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp 1623621585
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1623621585
transform 1 0 11684 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_111
timestamp 1623621585
transform 1 0 11316 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1623621585
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1623621585
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1623621585
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1623621585
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1623621585
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_144
timestamp 1623621585
transform 1 0 14352 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1623621585
transform 1 0 14996 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1623621585
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_156
timestamp 1623621585
transform 1 0 15456 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1623621585
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_172
timestamp 1623621585
transform 1 0 16928 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1623621585
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_168
timestamp 1623621585
transform 1 0 16560 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_180
timestamp 1623621585
transform 1 0 17664 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1623621585
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1623621585
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1623621585
transform 1 0 20240 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_192
timestamp 1623621585
transform 1 0 18768 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_201
timestamp 1623621585
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1623621585
transform 1 0 22080 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_220
timestamp 1623621585
transform 1 0 21344 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1623621585
transform 1 0 22172 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_213
timestamp 1623621585
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1623621585
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_241
timestamp 1623621585
transform 1 0 23276 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1623621585
transform 1 0 22908 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1623621585
transform 1 0 24012 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1623621585
transform 1 0 24748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1623621585
transform 1 0 24380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1623621585
transform 1 0 25484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_258
timestamp 1623621585
transform 1 0 24840 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_270
timestamp 1623621585
transform 1 0 25944 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1623621585
transform 1 0 27324 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1623621585
transform 1 0 26588 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_286
timestamp 1623621585
transform 1 0 27416 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_282
timestamp 1623621585
transform 1 0 27048 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_298
timestamp 1623621585
transform 1 0 28520 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_310
timestamp 1623621585
transform 1 0 29624 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_294
timestamp 1623621585
transform 1 0 28152 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_306
timestamp 1623621585
transform 1 0 29256 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1623621585
transform 1 0 29992 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_322
timestamp 1623621585
transform 1 0 30728 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_315
timestamp 1623621585
transform 1 0 30084 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_327
timestamp 1623621585
transform 1 0 31188 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1623621585
transform 1 0 32568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_334
timestamp 1623621585
transform 1 0 31832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_343
timestamp 1623621585
transform 1 0 32660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_339
timestamp 1623621585
transform 1 0 32292 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_351
timestamp 1623621585
transform 1 0 33396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1623621585
transform 1 0 35236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output671
timestamp 1623621585
transform 1 0 35236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_355
timestamp 1623621585
transform 1 0 33764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_367
timestamp 1623621585
transform 1 0 34868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_375
timestamp 1623621585
transform 1 0 35604 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_363
timestamp 1623621585
transform 1 0 34500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_372
timestamp 1623621585
transform 1 0 35328 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1623621585
transform 1 0 37076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1623621585
transform 1 0 37076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output652
timestamp 1623621585
transform 1 0 35972 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output655
timestamp 1623621585
transform 1 0 36340 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_383
timestamp 1623621585
transform 1 0 36340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1623621585
transform 1 0 37444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_380
timestamp 1623621585
transform 1 0 36064 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1623621585
transform 1 0 36708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_395
timestamp 1623621585
transform 1 0 37444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623621585
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623621585
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1623621585
transform 1 0 37812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1623621585
transform 1 0 37812 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_400
timestamp 1623621585
transform 1 0 37904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1623621585
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1623621585
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623621585
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input361
timestamp 1623621585
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_6
timestamp 1623621585
transform 1 0 1656 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_18
timestamp 1623621585
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1623621585
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1623621585
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1623621585
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_54
timestamp 1623621585
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_58
timestamp 1623621585
transform 1 0 6440 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_70
timestamp 1623621585
transform 1 0 7544 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_82
timestamp 1623621585
transform 1 0 8648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_94
timestamp 1623621585
transform 1 0 9752 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1623621585
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_106
timestamp 1623621585
transform 1 0 10856 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_115
timestamp 1623621585
transform 1 0 11684 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_127
timestamp 1623621585
transform 1 0 12788 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_139
timestamp 1623621585
transform 1 0 13892 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_151
timestamp 1623621585
transform 1 0 14996 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_163
timestamp 1623621585
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1623621585
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_172
timestamp 1623621585
transform 1 0 16928 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1623621585
transform 1 0 18032 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1623621585
transform 1 0 19136 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1623621585
transform 1 0 20240 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1623621585
transform 1 0 22080 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_220
timestamp 1623621585
transform 1 0 21344 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_229
timestamp 1623621585
transform 1 0 22172 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_241
timestamp 1623621585
transform 1 0 23276 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1623621585
transform 1 0 24380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1623621585
transform 1 0 25484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1623621585
transform 1 0 27324 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_277
timestamp 1623621585
transform 1 0 26588 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_286
timestamp 1623621585
transform 1 0 27416 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_298
timestamp 1623621585
transform 1 0 28520 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_310
timestamp 1623621585
transform 1 0 29624 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_322
timestamp 1623621585
transform 1 0 30728 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1623621585
transform 1 0 32568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_334
timestamp 1623621585
transform 1 0 31832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_343
timestamp 1623621585
transform 1 0 32660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_355
timestamp 1623621585
transform 1 0 33764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_367
timestamp 1623621585
transform 1 0 34868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1623621585
transform 1 0 37076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_379
timestamp 1623621585
transform 1 0 35972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1623621585
transform 1 0 37444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623621585
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1623621585
transform 1 0 37812 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_400
timestamp 1623621585
transform 1 0 37904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1623621585
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623621585
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1623621585
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1623621585
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1623621585
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1623621585
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1623621585
transform 1 0 3864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1623621585
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_54
timestamp 1623621585
transform 1 0 6072 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1623621585
transform 1 0 7176 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1623621585
transform 1 0 8280 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1623621585
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_87
timestamp 1623621585
transform 1 0 9108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1623621585
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_111
timestamp 1623621585
transform 1 0 11316 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1623621585
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1623621585
transform 1 0 14260 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1623621585
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1623621585
transform 1 0 14352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1623621585
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  _0782_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 16836 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1623621585
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_176
timestamp 1623621585
transform 1 0 17296 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1623621585
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_188
timestamp 1623621585
transform 1 0 18400 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_201
timestamp 1623621585
transform 1 0 19596 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_213
timestamp 1623621585
transform 1 0 20700 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1623621585
transform 1 0 21804 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1623621585
transform 1 0 22908 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1623621585
transform 1 0 24012 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1623621585
transform 1 0 24748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_258
timestamp 1623621585
transform 1 0 24840 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_270
timestamp 1623621585
transform 1 0 25944 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_282
timestamp 1623621585
transform 1 0 27048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_294
timestamp 1623621585
transform 1 0 28152 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_306
timestamp 1623621585
transform 1 0 29256 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1623621585
transform 1 0 29992 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_315
timestamp 1623621585
transform 1 0 30084 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_327
timestamp 1623621585
transform 1 0 31188 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_339
timestamp 1623621585
transform 1 0 32292 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_351
timestamp 1623621585
transform 1 0 33396 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1623621585
transform 1 0 35236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_363
timestamp 1623621585
transform 1 0 34500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_372
timestamp 1623621585
transform 1 0 35328 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1623621585
transform 1 0 37076 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_384
timestamp 1623621585
transform 1 0 36432 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_390
timestamp 1623621585
transform 1 0 36984 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_395
timestamp 1623621585
transform 1 0 37444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623621585
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1623621585
transform 1 0 37812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1623621585
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1623621585
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input362
timestamp 1623621585
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_6
timestamp 1623621585
transform 1 0 1656 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_18
timestamp 1623621585
transform 1 0 2760 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1623621585
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1623621585
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1623621585
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_54
timestamp 1623621585
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_58
timestamp 1623621585
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1623621585
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_82
timestamp 1623621585
transform 1 0 8648 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_94
timestamp 1623621585
transform 1 0 9752 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1623621585
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_106
timestamp 1623621585
transform 1 0 10856 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_115
timestamp 1623621585
transform 1 0 11684 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_127
timestamp 1623621585
transform 1 0 12788 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_139
timestamp 1623621585
transform 1 0 13892 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_151
timestamp 1623621585
transform 1 0 14996 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_163
timestamp 1623621585
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1623621585
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_172
timestamp 1623621585
transform 1 0 16928 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1623621585
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1623621585
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_208
timestamp 1623621585
transform 1 0 20240 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1623621585
transform 1 0 22080 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_220
timestamp 1623621585
transform 1 0 21344 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_229
timestamp 1623621585
transform 1 0 22172 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_241
timestamp 1623621585
transform 1 0 23276 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1623621585
transform 1 0 24380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1623621585
transform 1 0 25484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1623621585
transform 1 0 27324 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp 1623621585
transform 1 0 26588 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_286
timestamp 1623621585
transform 1 0 27416 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_298
timestamp 1623621585
transform 1 0 28520 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_310
timestamp 1623621585
transform 1 0 29624 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_322
timestamp 1623621585
transform 1 0 30728 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1623621585
transform 1 0 32568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_334
timestamp 1623621585
transform 1 0 31832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_343
timestamp 1623621585
transform 1 0 32660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_355
timestamp 1623621585
transform 1 0 33764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_367
timestamp 1623621585
transform 1 0 34868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1623621585
transform 1 0 37076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_379
timestamp 1623621585
transform 1 0 35972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1623621585
transform 1 0 37444 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1623621585
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1623621585
transform 1 0 37812 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_400
timestamp 1623621585
transform 1 0 37904 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1623621585
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1623621585
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input332
timestamp 1623621585
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_6
timestamp 1623621585
transform 1 0 1656 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_18
timestamp 1623621585
transform 1 0 2760 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1623621585
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_26
timestamp 1623621585
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1623621585
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1623621585
transform 1 0 4968 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_54
timestamp 1623621585
transform 1 0 6072 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_66
timestamp 1623621585
transform 1 0 7176 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_78
timestamp 1623621585
transform 1 0 8280 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1623621585
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1623621585
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 1623621585
transform 1 0 10212 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_111
timestamp 1623621585
transform 1 0 11316 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1623621585
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1623621585
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1623621585
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_144
timestamp 1623621585
transform 1 0 14352 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_156
timestamp 1623621585
transform 1 0 15456 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_168
timestamp 1623621585
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_180
timestamp 1623621585
transform 1 0 17664 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1623621585
transform 1 0 19504 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_192
timestamp 1623621585
transform 1 0 18768 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1623621585
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_213
timestamp 1623621585
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1623621585
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1623621585
transform 1 0 22908 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_249
timestamp 1623621585
transform 1 0 24012 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1623621585
transform 1 0 24748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_258
timestamp 1623621585
transform 1 0 24840 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_270
timestamp 1623621585
transform 1 0 25944 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_282
timestamp 1623621585
transform 1 0 27048 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_294
timestamp 1623621585
transform 1 0 28152 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_306
timestamp 1623621585
transform 1 0 29256 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1623621585
transform 1 0 29992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_315
timestamp 1623621585
transform 1 0 30084 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_327
timestamp 1623621585
transform 1 0 31188 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_339
timestamp 1623621585
transform 1 0 32292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_351
timestamp 1623621585
transform 1 0 33396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1623621585
transform 1 0 35236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_363
timestamp 1623621585
transform 1 0 34500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_372
timestamp 1623621585
transform 1 0 35328 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_384
timestamp 1623621585
transform 1 0 36432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1623621585
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1623621585
transform 1 0 37812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_396
timestamp 1623621585
transform 1 0 37536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1623621585
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1623621585
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1623621585
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1623621585
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1623621585
transform 1 0 3588 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1623621585
transform 1 0 4692 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1623621585
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_51
timestamp 1623621585
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_58
timestamp 1623621585
transform 1 0 6440 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1623621585
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_82
timestamp 1623621585
transform 1 0 8648 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_94
timestamp 1623621585
transform 1 0 9752 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1623621585
transform 1 0 11592 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_106
timestamp 1623621585
transform 1 0 10856 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1623621585
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_127
timestamp 1623621585
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_139
timestamp 1623621585
transform 1 0 13892 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_151
timestamp 1623621585
transform 1 0 14996 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_163
timestamp 1623621585
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1623621585
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_172
timestamp 1623621585
transform 1 0 16928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1623621585
transform 1 0 18032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1623621585
transform 1 0 19136 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_208
timestamp 1623621585
transform 1 0 20240 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1623621585
transform 1 0 22080 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_220
timestamp 1623621585
transform 1 0 21344 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_229
timestamp 1623621585
transform 1 0 22172 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_2  _0827_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22540 0 -1 9248
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_12_243
timestamp 1623621585
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_255
timestamp 1623621585
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_267
timestamp 1623621585
transform 1 0 25668 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1623621585
transform 1 0 27324 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_279
timestamp 1623621585
transform 1 0 26772 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_286
timestamp 1623621585
transform 1 0 27416 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_298
timestamp 1623621585
transform 1 0 28520 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_310
timestamp 1623621585
transform 1 0 29624 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_322
timestamp 1623621585
transform 1 0 30728 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1623621585
transform 1 0 32568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_334
timestamp 1623621585
transform 1 0 31832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_343
timestamp 1623621585
transform 1 0 32660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_355
timestamp 1623621585
transform 1 0 33764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_367
timestamp 1623621585
transform 1 0 34868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1623621585
transform 1 0 37076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_379
timestamp 1623621585
transform 1 0 35972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1623621585
transform 1 0 37444 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1623621585
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1623621585
transform 1 0 37812 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_400
timestamp 1623621585
transform 1 0 37904 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1623621585
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1623621585
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1623621585
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input333
timestamp 1623621585
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input334
timestamp 1623621585
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_6
timestamp 1623621585
transform 1 0 1656 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_18
timestamp 1623621585
transform 1 0 2760 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_6
timestamp 1623621585
transform 1 0 1656 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_18
timestamp 1623621585
transform 1 0 2760 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1623621585
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_26
timestamp 1623621585
transform 1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1623621585
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1623621585
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1623621585
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1623621585
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_54
timestamp 1623621585
transform 1 0 6072 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1623621585
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_54
timestamp 1623621585
transform 1 0 6072 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_58
timestamp 1623621585
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_66
timestamp 1623621585
transform 1 0 7176 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1623621585
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_70
timestamp 1623621585
transform 1 0 7544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_82
timestamp 1623621585
transform 1 0 8648 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1623621585
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_87
timestamp 1623621585
transform 1 0 9108 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_99
timestamp 1623621585
transform 1 0 10212 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_94
timestamp 1623621585
transform 1 0 9752 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1623621585
transform 1 0 11592 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_111
timestamp 1623621585
transform 1 0 11316 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1623621585
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_106
timestamp 1623621585
transform 1 0 10856 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1623621585
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1623621585
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1623621585
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_144
timestamp 1623621585
transform 1 0 14352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1623621585
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1623621585
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_156
timestamp 1623621585
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_151
timestamp 1623621585
transform 1 0 14996 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1623621585
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1623621585
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_168
timestamp 1623621585
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_180
timestamp 1623621585
transform 1 0 17664 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1623621585
transform 1 0 16928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1623621585
transform 1 0 18032 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1623621585
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_192
timestamp 1623621585
transform 1 0 18768 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_201
timestamp 1623621585
transform 1 0 19596 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_196
timestamp 1623621585
transform 1 0 19136 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_208
timestamp 1623621585
transform 1 0 20240 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1623621585
transform 1 0 22080 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_213
timestamp 1623621585
transform 1 0 20700 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1623621585
transform 1 0 21804 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_220
timestamp 1623621585
transform 1 0 21344 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_229
timestamp 1623621585
transform 1 0 22172 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1623621585
transform 1 0 22908 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_249
timestamp 1623621585
transform 1 0 24012 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_241
timestamp 1623621585
transform 1 0 23276 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1623621585
transform 1 0 24748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_258
timestamp 1623621585
transform 1 0 24840 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_270
timestamp 1623621585
transform 1 0 25944 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1623621585
transform 1 0 24380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1623621585
transform 1 0 25484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1623621585
transform 1 0 27324 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_282
timestamp 1623621585
transform 1 0 27048 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_277
timestamp 1623621585
transform 1 0 26588 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_286
timestamp 1623621585
transform 1 0 27416 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_294
timestamp 1623621585
transform 1 0 28152 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_306
timestamp 1623621585
transform 1 0 29256 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_298
timestamp 1623621585
transform 1 0 28520 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_310
timestamp 1623621585
transform 1 0 29624 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1623621585
transform 1 0 29992 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_315
timestamp 1623621585
transform 1 0 30084 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_327
timestamp 1623621585
transform 1 0 31188 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_322
timestamp 1623621585
transform 1 0 30728 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1623621585
transform 1 0 32568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_339
timestamp 1623621585
transform 1 0 32292 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_351
timestamp 1623621585
transform 1 0 33396 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_334
timestamp 1623621585
transform 1 0 31832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_343
timestamp 1623621585
transform 1 0 32660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1623621585
transform 1 0 35236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_363
timestamp 1623621585
transform 1 0 34500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_372
timestamp 1623621585
transform 1 0 35328 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_355
timestamp 1623621585
transform 1 0 33764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_367
timestamp 1623621585
transform 1 0 34868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1623621585
transform 1 0 37076 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1623621585
transform 1 0 37076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_384
timestamp 1623621585
transform 1 0 36432 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_390
timestamp 1623621585
transform 1 0 36984 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_395
timestamp 1623621585
transform 1 0 37444 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_379
timestamp 1623621585
transform 1 0 35972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_395
timestamp 1623621585
transform 1 0 37444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1623621585
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1623621585
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1623621585
transform 1 0 37812 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1623621585
transform 1 0 37812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1623621585
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_400
timestamp 1623621585
transform 1 0 37904 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1623621585
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1623621585
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1623621585
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1623621585
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1623621585
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1623621585
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1623621585
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1623621585
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_54
timestamp 1623621585
transform 1 0 6072 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_66
timestamp 1623621585
transform 1 0 7176 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1623621585
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1623621585
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_87
timestamp 1623621585
transform 1 0 9108 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_99
timestamp 1623621585
transform 1 0 10212 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_111
timestamp 1623621585
transform 1 0 11316 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1623621585
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1623621585
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_135
timestamp 1623621585
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1623621585
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1623621585
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1623621585
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_180
timestamp 1623621585
transform 1 0 17664 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1623621585
transform 1 0 19504 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_192
timestamp 1623621585
transform 1 0 18768 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_201
timestamp 1623621585
transform 1 0 19596 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_213
timestamp 1623621585
transform 1 0 20700 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1623621585
transform 1 0 21804 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1623621585
transform 1 0 22908 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_249
timestamp 1623621585
transform 1 0 24012 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1623621585
transform 1 0 24748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_258
timestamp 1623621585
transform 1 0 24840 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_270
timestamp 1623621585
transform 1 0 25944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_282
timestamp 1623621585
transform 1 0 27048 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_294
timestamp 1623621585
transform 1 0 28152 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_306
timestamp 1623621585
transform 1 0 29256 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1623621585
transform 1 0 29992 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_315
timestamp 1623621585
transform 1 0 30084 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_327
timestamp 1623621585
transform 1 0 31188 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_339
timestamp 1623621585
transform 1 0 32292 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_351
timestamp 1623621585
transform 1 0 33396 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1623621585
transform 1 0 35236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_363
timestamp 1623621585
transform 1 0 34500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_372
timestamp 1623621585
transform 1 0 35328 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_384
timestamp 1623621585
transform 1 0 36432 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1623621585
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1623621585
transform 1 0 37812 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_396
timestamp 1623621585
transform 1 0 37536 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1623621585
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1623621585
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input335
timestamp 1623621585
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_6
timestamp 1623621585
transform 1 0 1656 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_18
timestamp 1623621585
transform 1 0 2760 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1623621585
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1623621585
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1623621585
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_54
timestamp 1623621585
transform 1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_58
timestamp 1623621585
transform 1 0 6440 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1623621585
transform 1 0 7544 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_82
timestamp 1623621585
transform 1 0 8648 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_94
timestamp 1623621585
transform 1 0 9752 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1623621585
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_106
timestamp 1623621585
transform 1 0 10856 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_115
timestamp 1623621585
transform 1 0 11684 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_127
timestamp 1623621585
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1623621585
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_151
timestamp 1623621585
transform 1 0 14996 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_163
timestamp 1623621585
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1623621585
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_172
timestamp 1623621585
transform 1 0 16928 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1623621585
transform 1 0 18032 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_196
timestamp 1623621585
transform 1 0 19136 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_208
timestamp 1623621585
transform 1 0 20240 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1623621585
transform 1 0 22080 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_220
timestamp 1623621585
transform 1 0 21344 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1623621585
transform 1 0 22172 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_241
timestamp 1623621585
transform 1 0 23276 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1623621585
transform 1 0 24380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1623621585
transform 1 0 25484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1623621585
transform 1 0 27324 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_277
timestamp 1623621585
transform 1 0 26588 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_286
timestamp 1623621585
transform 1 0 27416 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_298
timestamp 1623621585
transform 1 0 28520 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_310
timestamp 1623621585
transform 1 0 29624 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_322
timestamp 1623621585
transform 1 0 30728 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1623621585
transform 1 0 32568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_334
timestamp 1623621585
transform 1 0 31832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_343
timestamp 1623621585
transform 1 0 32660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_355
timestamp 1623621585
transform 1 0 33764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_367
timestamp 1623621585
transform 1 0 34868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1623621585
transform 1 0 37076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_379
timestamp 1623621585
transform 1 0 35972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1623621585
transform 1 0 37444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1623621585
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1623621585
transform 1 0 37812 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_400
timestamp 1623621585
transform 1 0 37904 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1623621585
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1623621585
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1623621585
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1623621585
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1623621585
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1623621585
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1623621585
transform 1 0 3864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1623621585
transform 1 0 4968 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_54
timestamp 1623621585
transform 1 0 6072 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_66
timestamp 1623621585
transform 1 0 7176 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_78
timestamp 1623621585
transform 1 0 8280 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1623621585
transform 1 0 9016 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_87
timestamp 1623621585
transform 1 0 9108 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_99
timestamp 1623621585
transform 1 0 10212 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_111
timestamp 1623621585
transform 1 0 11316 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1623621585
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1623621585
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1623621585
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_144
timestamp 1623621585
transform 1 0 14352 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_156
timestamp 1623621585
transform 1 0 15456 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_168
timestamp 1623621585
transform 1 0 16560 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_180
timestamp 1623621585
transform 1 0 17664 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1623621585
transform 1 0 19504 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_192
timestamp 1623621585
transform 1 0 18768 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_201
timestamp 1623621585
transform 1 0 19596 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_213
timestamp 1623621585
transform 1 0 20700 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1623621585
transform 1 0 21804 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1623621585
transform 1 0 22908 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_249
timestamp 1623621585
transform 1 0 24012 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1623621585
transform 1 0 24748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_258
timestamp 1623621585
transform 1 0 24840 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_270
timestamp 1623621585
transform 1 0 25944 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_282
timestamp 1623621585
transform 1 0 27048 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_294
timestamp 1623621585
transform 1 0 28152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1623621585
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1623621585
transform 1 0 29992 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_315
timestamp 1623621585
transform 1 0 30084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_327
timestamp 1623621585
transform 1 0 31188 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_339
timestamp 1623621585
transform 1 0 32292 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_351
timestamp 1623621585
transform 1 0 33396 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1623621585
transform 1 0 35236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_363
timestamp 1623621585
transform 1 0 34500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_372
timestamp 1623621585
transform 1 0 35328 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1623621585
transform 1 0 37076 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_384
timestamp 1623621585
transform 1 0 36432 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_390
timestamp 1623621585
transform 1 0 36984 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_395
timestamp 1623621585
transform 1 0 37444 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1623621585
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1623621585
transform 1 0 37812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1623621585
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1623621585
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input336
timestamp 1623621585
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_6
timestamp 1623621585
transform 1 0 1656 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_18
timestamp 1623621585
transform 1 0 2760 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1623621585
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1623621585
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1623621585
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_54
timestamp 1623621585
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1623621585
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_70
timestamp 1623621585
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_82
timestamp 1623621585
transform 1 0 8648 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_94
timestamp 1623621585
transform 1 0 9752 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1623621585
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1623621585
transform 1 0 10856 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_115
timestamp 1623621585
transform 1 0 11684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1623621585
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_139
timestamp 1623621585
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1623621585
transform 1 0 14996 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1623621585
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1623621585
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_172
timestamp 1623621585
transform 1 0 16928 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_184
timestamp 1623621585
transform 1 0 18032 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_196
timestamp 1623621585
transform 1 0 19136 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_208
timestamp 1623621585
transform 1 0 20240 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1623621585
transform 1 0 22080 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_220
timestamp 1623621585
transform 1 0 21344 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_229
timestamp 1623621585
transform 1 0 22172 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_241
timestamp 1623621585
transform 1 0 23276 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1623621585
transform 1 0 24380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1623621585
transform 1 0 25484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1623621585
transform 1 0 27324 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_277
timestamp 1623621585
transform 1 0 26588 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_286
timestamp 1623621585
transform 1 0 27416 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_298
timestamp 1623621585
transform 1 0 28520 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_310
timestamp 1623621585
transform 1 0 29624 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_322
timestamp 1623621585
transform 1 0 30728 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1623621585
transform 1 0 32568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_334
timestamp 1623621585
transform 1 0 31832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_343
timestamp 1623621585
transform 1 0 32660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_355
timestamp 1623621585
transform 1 0 33764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_367
timestamp 1623621585
transform 1 0 34868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1623621585
transform 1 0 37076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_379
timestamp 1623621585
transform 1 0 35972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_395
timestamp 1623621585
transform 1 0 37444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1623621585
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1623621585
transform 1 0 37812 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_400
timestamp 1623621585
transform 1 0 37904 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1623621585
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1623621585
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1623621585
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input337
timestamp 1623621585
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_6
timestamp 1623621585
transform 1 0 1656 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_18
timestamp 1623621585
transform 1 0 2760 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1623621585
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1623621585
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1623621585
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_26
timestamp 1623621585
transform 1 0 3496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1623621585
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1623621585
transform 1 0 3588 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1623621585
transform 1 0 4692 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1623621585
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1623621585
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_54
timestamp 1623621585
transform 1 0 6072 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_51
timestamp 1623621585
transform 1 0 5796 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_58
timestamp 1623621585
transform 1 0 6440 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1623621585
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 1623621585
transform 1 0 8280 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_70
timestamp 1623621585
transform 1 0 7544 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_82
timestamp 1623621585
transform 1 0 8648 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1623621585
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_87
timestamp 1623621585
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_99
timestamp 1623621585
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_94
timestamp 1623621585
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1623621585
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_111
timestamp 1623621585
transform 1 0 11316 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1623621585
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_106
timestamp 1623621585
transform 1 0 10856 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_115
timestamp 1623621585
transform 1 0 11684 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1623621585
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1623621585
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_144
timestamp 1623621585
transform 1 0 14352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1623621585
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_139
timestamp 1623621585
transform 1 0 13892 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_156
timestamp 1623621585
transform 1 0 15456 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_151
timestamp 1623621585
transform 1 0 14996 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_163
timestamp 1623621585
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1623621585
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_168
timestamp 1623621585
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_180
timestamp 1623621585
transform 1 0 17664 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_172
timestamp 1623621585
transform 1 0 16928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1623621585
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1623621585
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_192
timestamp 1623621585
transform 1 0 18768 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_201
timestamp 1623621585
transform 1 0 19596 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1623621585
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_208
timestamp 1623621585
transform 1 0 20240 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_2  _0801_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20976 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1623621585
transform 1 0 22080 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_213
timestamp 1623621585
transform 1 0 20700 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1623621585
transform 1 0 21804 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_220
timestamp 1623621585
transform 1 0 21344 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_229
timestamp 1623621585
transform 1 0 22172 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1623621585
transform 1 0 22908 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_249
timestamp 1623621585
transform 1 0 24012 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_241
timestamp 1623621585
transform 1 0 23276 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1623621585
transform 1 0 24748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_258
timestamp 1623621585
transform 1 0 24840 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_270
timestamp 1623621585
transform 1 0 25944 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1623621585
transform 1 0 24380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1623621585
transform 1 0 25484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1623621585
transform 1 0 27324 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_282
timestamp 1623621585
transform 1 0 27048 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_277
timestamp 1623621585
transform 1 0 26588 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_286
timestamp 1623621585
transform 1 0 27416 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_294
timestamp 1623621585
transform 1 0 28152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_306
timestamp 1623621585
transform 1 0 29256 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_298
timestamp 1623621585
transform 1 0 28520 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_310
timestamp 1623621585
transform 1 0 29624 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1623621585
transform 1 0 29992 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_315
timestamp 1623621585
transform 1 0 30084 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_327
timestamp 1623621585
transform 1 0 31188 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_322
timestamp 1623621585
transform 1 0 30728 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1623621585
transform 1 0 32568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_339
timestamp 1623621585
transform 1 0 32292 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_351
timestamp 1623621585
transform 1 0 33396 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_334
timestamp 1623621585
transform 1 0 31832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_343
timestamp 1623621585
transform 1 0 32660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1623621585
transform 1 0 35236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_363
timestamp 1623621585
transform 1 0 34500 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_372
timestamp 1623621585
transform 1 0 35328 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_355
timestamp 1623621585
transform 1 0 33764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_367
timestamp 1623621585
transform 1 0 34868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1623621585
transform 1 0 37076 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_384
timestamp 1623621585
transform 1 0 36432 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_379
timestamp 1623621585
transform 1 0 35972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1623621585
transform 1 0 37444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1623621585
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1623621585
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1623621585
transform 1 0 37812 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1623621585
transform 1 0 37812 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_396
timestamp 1623621585
transform 1 0 37536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1623621585
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_400
timestamp 1623621585
transform 1 0 37904 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1623621585
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1623621585
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input338
timestamp 1623621585
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_6
timestamp 1623621585
transform 1 0 1656 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_18
timestamp 1623621585
transform 1 0 2760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1623621585
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_26
timestamp 1623621585
transform 1 0 3496 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_30
timestamp 1623621585
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1623621585
transform 1 0 4968 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_54
timestamp 1623621585
transform 1 0 6072 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_66
timestamp 1623621585
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_78
timestamp 1623621585
transform 1 0 8280 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1623621585
transform 1 0 9016 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_87
timestamp 1623621585
transform 1 0 9108 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_99
timestamp 1623621585
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_111
timestamp 1623621585
transform 1 0 11316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1623621585
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1623621585
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1623621585
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_144
timestamp 1623621585
transform 1 0 14352 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_156
timestamp 1623621585
transform 1 0 15456 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_168
timestamp 1623621585
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_180
timestamp 1623621585
transform 1 0 17664 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1623621585
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_192
timestamp 1623621585
transform 1 0 18768 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_201
timestamp 1623621585
transform 1 0 19596 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_213
timestamp 1623621585
transform 1 0 20700 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1623621585
transform 1 0 21804 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1623621585
transform 1 0 22908 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 1623621585
transform 1 0 24012 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1623621585
transform 1 0 24748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_258
timestamp 1623621585
transform 1 0 24840 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_270
timestamp 1623621585
transform 1 0 25944 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_282
timestamp 1623621585
transform 1 0 27048 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_294
timestamp 1623621585
transform 1 0 28152 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_306
timestamp 1623621585
transform 1 0 29256 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1623621585
transform 1 0 29992 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_315
timestamp 1623621585
transform 1 0 30084 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_327
timestamp 1623621585
transform 1 0 31188 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_339
timestamp 1623621585
transform 1 0 32292 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_351
timestamp 1623621585
transform 1 0 33396 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1623621585
transform 1 0 35236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_363
timestamp 1623621585
transform 1 0 34500 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_372
timestamp 1623621585
transform 1 0 35328 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1623621585
transform 1 0 37076 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_384
timestamp 1623621585
transform 1 0 36432 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_390
timestamp 1623621585
transform 1 0 36984 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_395
timestamp 1623621585
transform 1 0 37444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1623621585
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1623621585
transform 1 0 37812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1623621585
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1623621585
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input339
timestamp 1623621585
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_6
timestamp 1623621585
transform 1 0 1656 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_18
timestamp 1623621585
transform 1 0 2760 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1623621585
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1623621585
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1623621585
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_54
timestamp 1623621585
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_58
timestamp 1623621585
transform 1 0 6440 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_70
timestamp 1623621585
transform 1 0 7544 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_82
timestamp 1623621585
transform 1 0 8648 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1623621585
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1623621585
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1623621585
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1623621585
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_127
timestamp 1623621585
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_139
timestamp 1623621585
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_151
timestamp 1623621585
transform 1 0 14996 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_163
timestamp 1623621585
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1623621585
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1623621585
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1623621585
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_196
timestamp 1623621585
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_208
timestamp 1623621585
transform 1 0 20240 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1623621585
transform 1 0 22080 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_220
timestamp 1623621585
transform 1 0 21344 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_229
timestamp 1623621585
transform 1 0 22172 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_241
timestamp 1623621585
transform 1 0 23276 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1623621585
transform 1 0 24380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1623621585
transform 1 0 25484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1623621585
transform 1 0 27324 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_277
timestamp 1623621585
transform 1 0 26588 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_286
timestamp 1623621585
transform 1 0 27416 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0915_
timestamp 1623621585
transform 1 0 28980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1623621585
transform 1 0 28520 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_302
timestamp 1623621585
transform 1 0 28888 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_306
timestamp 1623621585
transform 1 0 29256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_318
timestamp 1623621585
transform 1 0 30360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_330
timestamp 1623621585
transform 1 0 31464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1623621585
transform 1 0 32568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_343
timestamp 1623621585
transform 1 0 32660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_355
timestamp 1623621585
transform 1 0 33764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_367
timestamp 1623621585
transform 1 0 34868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_379
timestamp 1623621585
transform 1 0 35972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_391
timestamp 1623621585
transform 1 0 37076 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1623621585
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1623621585
transform 1 0 37812 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_400
timestamp 1623621585
transform 1 0 37904 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1623621585
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1623621585
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1623621585
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1623621585
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1623621585
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1623621585
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_30
timestamp 1623621585
transform 1 0 3864 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1623621585
transform 1 0 4968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_54
timestamp 1623621585
transform 1 0 6072 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_66
timestamp 1623621585
transform 1 0 7176 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_78
timestamp 1623621585
transform 1 0 8280 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1623621585
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_87
timestamp 1623621585
transform 1 0 9108 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1623621585
transform 1 0 10212 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_111
timestamp 1623621585
transform 1 0 11316 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1623621585
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1623621585
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1623621585
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_144
timestamp 1623621585
transform 1 0 14352 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_156
timestamp 1623621585
transform 1 0 15456 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_164
timestamp 1623621585
transform 1 0 16192 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 16468 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0732_
timestamp 1623621585
transform 1 0 17572 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1623621585
transform 1 0 17204 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_187
timestamp 1623621585
transform 1 0 18308 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1623621585
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1623621585
transform 1 0 19412 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_201
timestamp 1623621585
transform 1 0 19596 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_213
timestamp 1623621585
transform 1 0 20700 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1623621585
transform 1 0 21804 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1623621585
transform 1 0 22908 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_249
timestamp 1623621585
transform 1 0 24012 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1623621585
transform 1 0 24748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_258
timestamp 1623621585
transform 1 0 24840 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_270
timestamp 1623621585
transform 1 0 25944 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_282
timestamp 1623621585
transform 1 0 27048 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_294
timestamp 1623621585
transform 1 0 28152 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_306
timestamp 1623621585
transform 1 0 29256 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1623621585
transform 1 0 29992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_315
timestamp 1623621585
transform 1 0 30084 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_327
timestamp 1623621585
transform 1 0 31188 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_339
timestamp 1623621585
transform 1 0 32292 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_351
timestamp 1623621585
transform 1 0 33396 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1623621585
transform 1 0 35236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_363
timestamp 1623621585
transform 1 0 34500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_372
timestamp 1623621585
transform 1 0 35328 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1623621585
transform 1 0 37260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_384
timestamp 1623621585
transform 1 0 36432 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_392
timestamp 1623621585
transform 1 0 37168 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1623621585
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1623621585
transform 1 0 37904 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_396
timestamp 1623621585
transform 1 0 37536 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1623621585
transform 1 0 38180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1623621585
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input340
timestamp 1623621585
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_6
timestamp 1623621585
transform 1 0 1656 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_18
timestamp 1623621585
transform 1 0 2760 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1623621585
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1623621585
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1623621585
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_54
timestamp 1623621585
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_58
timestamp 1623621585
transform 1 0 6440 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_70
timestamp 1623621585
transform 1 0 7544 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_82
timestamp 1623621585
transform 1 0 8648 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_94
timestamp 1623621585
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1623621585
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_106
timestamp 1623621585
transform 1 0 10856 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_115
timestamp 1623621585
transform 1 0 11684 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_127
timestamp 1623621585
transform 1 0 12788 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_139
timestamp 1623621585
transform 1 0 13892 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0741_
timestamp 1623621585
transform 1 0 15732 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_151
timestamp 1623621585
transform 1 0 14996 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0716_
timestamp 1623621585
transform 1 0 17296 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1623621585
transform 1 0 16836 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1623621585
transform 1 0 16468 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1623621585
transform 1 0 16928 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1623621585
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_196
timestamp 1623621585
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_208
timestamp 1623621585
transform 1 0 20240 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1623621585
transform 1 0 22080 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_220
timestamp 1623621585
transform 1 0 21344 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_229
timestamp 1623621585
transform 1 0 22172 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_241
timestamp 1623621585
transform 1 0 23276 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1623621585
transform 1 0 24380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1623621585
transform 1 0 25484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1623621585
transform 1 0 27324 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_277
timestamp 1623621585
transform 1 0 26588 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_286
timestamp 1623621585
transform 1 0 27416 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_298
timestamp 1623621585
transform 1 0 28520 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_310
timestamp 1623621585
transform 1 0 29624 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_322
timestamp 1623621585
transform 1 0 30728 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1623621585
transform 1 0 32568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_334
timestamp 1623621585
transform 1 0 31832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_343
timestamp 1623621585
transform 1 0 32660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_355
timestamp 1623621585
transform 1 0 33764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_367
timestamp 1623621585
transform 1 0 34868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1623621585
transform 1 0 37076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_379
timestamp 1623621585
transform 1 0 35972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_395
timestamp 1623621585
transform 1 0 37444 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1623621585
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1623621585
transform 1 0 37812 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_400
timestamp 1623621585
transform 1 0 37904 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1623621585
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1623621585
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input341
timestamp 1623621585
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_6
timestamp 1623621585
transform 1 0 1656 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_18
timestamp 1623621585
transform 1 0 2760 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1623621585
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_26
timestamp 1623621585
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_30
timestamp 1623621585
transform 1 0 3864 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_42
timestamp 1623621585
transform 1 0 4968 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_54
timestamp 1623621585
transform 1 0 6072 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_66
timestamp 1623621585
transform 1 0 7176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_78
timestamp 1623621585
transform 1 0 8280 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1623621585
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1623621585
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_99
timestamp 1623621585
transform 1 0 10212 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_111
timestamp 1623621585
transform 1 0 11316 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1623621585
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1623621585
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1623621585
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1623621585
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1623621585
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0698_
timestamp 1623621585
transform 1 0 16560 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_176
timestamp 1623621585
transform 1 0 17296 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1623621585
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_188
timestamp 1623621585
transform 1 0 18400 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_201
timestamp 1623621585
transform 1 0 19596 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_213
timestamp 1623621585
transform 1 0 20700 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1623621585
transform 1 0 21804 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1623621585
transform 1 0 22908 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1623621585
transform 1 0 24012 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1623621585
transform 1 0 24748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_258
timestamp 1623621585
transform 1 0 24840 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_270
timestamp 1623621585
transform 1 0 25944 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_282
timestamp 1623621585
transform 1 0 27048 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_294
timestamp 1623621585
transform 1 0 28152 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_306
timestamp 1623621585
transform 1 0 29256 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1623621585
transform 1 0 29992 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_315
timestamp 1623621585
transform 1 0 30084 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_327
timestamp 1623621585
transform 1 0 31188 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_339
timestamp 1623621585
transform 1 0 32292 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_351
timestamp 1623621585
transform 1 0 33396 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1623621585
transform 1 0 35236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_363
timestamp 1623621585
transform 1 0 34500 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_372
timestamp 1623621585
transform 1 0 35328 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1623621585
transform 1 0 37260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1623621585
transform 1 0 36432 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_392
timestamp 1623621585
transform 1 0 37168 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1623621585
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1623621585
transform 1 0 37904 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_396
timestamp 1623621585
transform 1 0 37536 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1623621585
transform 1 0 38180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1623621585
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1623621585
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input343
timestamp 1623621585
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1623621585
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1623621585
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_6
timestamp 1623621585
transform 1 0 1656 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_18
timestamp 1623621585
transform 1 0 2760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1623621585
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1623621585
transform 1 0 3588 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1623621585
transform 1 0 4692 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_26
timestamp 1623621585
transform 1 0 3496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_30
timestamp 1623621585
transform 1 0 3864 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1623621585
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_51
timestamp 1623621585
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_58
timestamp 1623621585
transform 1 0 6440 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_42
timestamp 1623621585
transform 1 0 4968 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_54
timestamp 1623621585
transform 1 0 6072 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_70
timestamp 1623621585
transform 1 0 7544 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_82
timestamp 1623621585
transform 1 0 8648 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_66
timestamp 1623621585
transform 1 0 7176 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_78
timestamp 1623621585
transform 1 0 8280 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1623621585
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_94
timestamp 1623621585
transform 1 0 9752 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_87
timestamp 1623621585
transform 1 0 9108 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_99
timestamp 1623621585
transform 1 0 10212 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1623621585
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_106
timestamp 1623621585
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_115
timestamp 1623621585
transform 1 0 11684 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_111
timestamp 1623621585
transform 1 0 11316 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1623621585
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1623621585
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1623621585
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1623621585
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1623621585
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1623621585
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_151
timestamp 1623621585
transform 1 0 14996 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_163
timestamp 1623621585
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1623621585
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1623621585
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1623621585
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1623621585
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1623621585
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_180
timestamp 1623621585
transform 1 0 17664 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1623621585
transform 1 0 19504 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1623621585
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_208
timestamp 1623621585
transform 1 0 20240 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_192
timestamp 1623621585
transform 1 0 18768 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_201
timestamp 1623621585
transform 1 0 19596 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _0829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 21252 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1623621585
transform 1 0 22080 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1623621585
transform 1 0 21344 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_229
timestamp 1623621585
transform 1 0 22172 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_213
timestamp 1623621585
transform 1 0 20700 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_227
timestamp 1623621585
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_241
timestamp 1623621585
transform 1 0 23276 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_239
timestamp 1623621585
transform 1 0 23092 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1623621585
transform 1 0 24748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1623621585
transform 1 0 24380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1623621585
transform 1 0 25484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_251
timestamp 1623621585
transform 1 0 24196 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_258
timestamp 1623621585
transform 1 0 24840 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_270
timestamp 1623621585
transform 1 0 25944 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1623621585
transform 1 0 27324 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1623621585
transform 1 0 26588 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_286
timestamp 1623621585
transform 1 0 27416 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_282
timestamp 1623621585
transform 1 0 27048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_298
timestamp 1623621585
transform 1 0 28520 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_310
timestamp 1623621585
transform 1 0 29624 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_294
timestamp 1623621585
transform 1 0 28152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_306
timestamp 1623621585
transform 1 0 29256 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1623621585
transform 1 0 29992 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_322
timestamp 1623621585
transform 1 0 30728 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_315
timestamp 1623621585
transform 1 0 30084 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_327
timestamp 1623621585
transform 1 0 31188 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1623621585
transform 1 0 32568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_334
timestamp 1623621585
transform 1 0 31832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_343
timestamp 1623621585
transform 1 0 32660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_339
timestamp 1623621585
transform 1 0 32292 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_351
timestamp 1623621585
transform 1 0 33396 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1623621585
transform 1 0 35236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_355
timestamp 1623621585
transform 1 0 33764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_367
timestamp 1623621585
transform 1 0 34868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_363
timestamp 1623621585
transform 1 0 34500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_372
timestamp 1623621585
transform 1 0 35328 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input161
timestamp 1623621585
transform 1 0 37260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input193
timestamp 1623621585
transform 1 0 37076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_379
timestamp 1623621585
transform 1 0 35972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1623621585
transform 1 0 37444 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_384
timestamp 1623621585
transform 1 0 36432 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_392
timestamp 1623621585
transform 1 0 37168 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1623621585
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1623621585
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1623621585
transform 1 0 37812 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1623621585
transform 1 0 37904 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_400
timestamp 1623621585
transform 1 0 37904 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1623621585
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_396
timestamp 1623621585
transform 1 0 37536 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1623621585
transform 1 0 38180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1623621585
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input344
timestamp 1623621585
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_6
timestamp 1623621585
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1623621585
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1623621585
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1623621585
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1623621585
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_54
timestamp 1623621585
transform 1 0 6072 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_58
timestamp 1623621585
transform 1 0 6440 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_70
timestamp 1623621585
transform 1 0 7544 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_82
timestamp 1623621585
transform 1 0 8648 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_94
timestamp 1623621585
transform 1 0 9752 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1623621585
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1623621585
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_115
timestamp 1623621585
transform 1 0 11684 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_127
timestamp 1623621585
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_139
timestamp 1623621585
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_151
timestamp 1623621585
transform 1 0 14996 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1623621585
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0687_
timestamp 1623621585
transform 1 0 17296 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1623621585
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1623621585
transform 1 0 16928 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1623621585
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _0986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19780 0 -1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_28_196
timestamp 1623621585
transform 1 0 19136 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_202
timestamp 1623621585
transform 1 0 19688 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1623621585
transform 1 0 22080 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_220
timestamp 1623621585
transform 1 0 21344 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_229
timestamp 1623621585
transform 1 0 22172 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_241
timestamp 1623621585
transform 1 0 23276 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1623621585
transform 1 0 24380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1623621585
transform 1 0 25484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1623621585
transform 1 0 27324 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_277
timestamp 1623621585
transform 1 0 26588 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_286
timestamp 1623621585
transform 1 0 27416 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_298
timestamp 1623621585
transform 1 0 28520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_310
timestamp 1623621585
transform 1 0 29624 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_322
timestamp 1623621585
transform 1 0 30728 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1623621585
transform 1 0 32568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_334
timestamp 1623621585
transform 1 0 31832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_343
timestamp 1623621585
transform 1 0 32660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_355
timestamp 1623621585
transform 1 0 33764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_367
timestamp 1623621585
transform 1 0 34868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input196
timestamp 1623621585
transform 1 0 37168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_379
timestamp 1623621585
transform 1 0 35972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_391
timestamp 1623621585
transform 1 0 37076 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1623621585
transform 1 0 37444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1623621585
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1623621585
transform 1 0 37812 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_400
timestamp 1623621585
transform 1 0 37904 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1623621585
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1623621585
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1623621585
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1623621585
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1623621585
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1623621585
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1623621585
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1623621585
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_54
timestamp 1623621585
transform 1 0 6072 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_66
timestamp 1623621585
transform 1 0 7176 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_78
timestamp 1623621585
transform 1 0 8280 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1623621585
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_87
timestamp 1623621585
transform 1 0 9108 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_99
timestamp 1623621585
transform 1 0 10212 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_111
timestamp 1623621585
transform 1 0 11316 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1623621585
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1623621585
transform 1 0 14260 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1623621585
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_144
timestamp 1623621585
transform 1 0 14352 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_156
timestamp 1623621585
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0678_
timestamp 1623621585
transform 1 0 16560 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_8  _0797_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17664 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_176
timestamp 1623621585
transform 1 0 17296 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0984_
timestamp 1623621585
transform 1 0 19964 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1623621585
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_196
timestamp 1623621585
transform 1 0 19136 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1623621585
transform 1 0 19596 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_222
timestamp 1623621585
transform 1 0 21528 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_234
timestamp 1623621585
transform 1 0 22632 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_246
timestamp 1623621585
transform 1 0 23736 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1623621585
transform 1 0 24748 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_254
timestamp 1623621585
transform 1 0 24472 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_258
timestamp 1623621585
transform 1 0 24840 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_270
timestamp 1623621585
transform 1 0 25944 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_282
timestamp 1623621585
transform 1 0 27048 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_294
timestamp 1623621585
transform 1 0 28152 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_306
timestamp 1623621585
transform 1 0 29256 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1623621585
transform 1 0 29992 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_315
timestamp 1623621585
transform 1 0 30084 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_327
timestamp 1623621585
transform 1 0 31188 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_339
timestamp 1623621585
transform 1 0 32292 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_351
timestamp 1623621585
transform 1 0 33396 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1623621585
transform 1 0 35236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_363
timestamp 1623621585
transform 1 0 34500 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_372
timestamp 1623621585
transform 1 0 35328 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_384
timestamp 1623621585
transform 1 0 36432 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1623621585
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1623621585
transform 1 0 37904 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_396
timestamp 1623621585
transform 1 0 37536 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1623621585
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1623621585
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input345
timestamp 1623621585
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_6
timestamp 1623621585
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_18
timestamp 1623621585
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1623621585
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1623621585
transform 1 0 6348 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1623621585
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_54
timestamp 1623621585
transform 1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_58
timestamp 1623621585
transform 1 0 6440 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_70
timestamp 1623621585
transform 1 0 7544 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_82
timestamp 1623621585
transform 1 0 8648 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_94
timestamp 1623621585
transform 1 0 9752 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1623621585
transform 1 0 11592 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_106
timestamp 1623621585
transform 1 0 10856 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_115
timestamp 1623621585
transform 1 0 11684 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_127
timestamp 1623621585
transform 1 0 12788 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_139
timestamp 1623621585
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0765_
timestamp 1623621585
transform 1 0 15732 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_151
timestamp 1623621585
transform 1 0 14996 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0662_
timestamp 1623621585
transform 1 0 17296 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1623621585
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1623621585
transform 1 0 16468 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1623621585
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1623621585
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0670_
timestamp 1623621585
transform 1 0 18400 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _0985_
timestamp 1623621585
transform 1 0 19504 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1623621585
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1623621585
transform 1 0 22080 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_217
timestamp 1623621585
transform 1 0 21068 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_225
timestamp 1623621585
transform 1 0 21804 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_229
timestamp 1623621585
transform 1 0 22172 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_241
timestamp 1623621585
transform 1 0 23276 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1623621585
transform 1 0 24380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1623621585
transform 1 0 25484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1623621585
transform 1 0 27324 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp 1623621585
transform 1 0 26588 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_286
timestamp 1623621585
transform 1 0 27416 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_298
timestamp 1623621585
transform 1 0 28520 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_310
timestamp 1623621585
transform 1 0 29624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_322
timestamp 1623621585
transform 1 0 30728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1623621585
transform 1 0 32568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_334
timestamp 1623621585
transform 1 0 31832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_343
timestamp 1623621585
transform 1 0 32660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_355
timestamp 1623621585
transform 1 0 33764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_367
timestamp 1623621585
transform 1 0 34868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input164
timestamp 1623621585
transform 1 0 37168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_379
timestamp 1623621585
transform 1 0 35972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_391
timestamp 1623621585
transform 1 0 37076 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_395
timestamp 1623621585
transform 1 0 37444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1623621585
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1623621585
transform 1 0 37812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_400
timestamp 1623621585
transform 1 0 37904 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1623621585
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1623621585
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input346
timestamp 1623621585
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_6
timestamp 1623621585
transform 1 0 1656 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_18
timestamp 1623621585
transform 1 0 2760 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1623621585
transform 1 0 3772 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_26
timestamp 1623621585
transform 1 0 3496 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_30
timestamp 1623621585
transform 1 0 3864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1623621585
transform 1 0 4968 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_54
timestamp 1623621585
transform 1 0 6072 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_66
timestamp 1623621585
transform 1 0 7176 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_78
timestamp 1623621585
transform 1 0 8280 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1623621585
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_87
timestamp 1623621585
transform 1 0 9108 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_99
timestamp 1623621585
transform 1 0 10212 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_111
timestamp 1623621585
transform 1 0 11316 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1623621585
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1623621585
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1623621585
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_144
timestamp 1623621585
transform 1 0 14352 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0749_
timestamp 1623621585
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_156
timestamp 1623621585
transform 1 0 15456 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_162
timestamp 1623621585
transform 1 0 16008 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _0644_
timestamp 1623621585
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_171
timestamp 1623621585
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_183
timestamp 1623621585
transform 1 0 17940 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1623621585
transform 1 0 19964 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1623621585
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1623621585
transform 1 0 19044 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1623621585
transform 1 0 19412 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1623621585
transform 1 0 19596 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0988_
timestamp 1623621585
transform 1 0 21896 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_31_222
timestamp 1623621585
transform 1 0 21528 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_243
timestamp 1623621585
transform 1 0 23460 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1623621585
transform 1 0 24748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_255
timestamp 1623621585
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_258
timestamp 1623621585
transform 1 0 24840 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_270
timestamp 1623621585
transform 1 0 25944 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_282
timestamp 1623621585
transform 1 0 27048 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_294
timestamp 1623621585
transform 1 0 28152 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_306
timestamp 1623621585
transform 1 0 29256 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1623621585
transform 1 0 29992 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_315
timestamp 1623621585
transform 1 0 30084 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_327
timestamp 1623621585
transform 1 0 31188 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_339
timestamp 1623621585
transform 1 0 32292 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_351
timestamp 1623621585
transform 1 0 33396 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1623621585
transform 1 0 35236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_363
timestamp 1623621585
transform 1 0 34500 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_372
timestamp 1623621585
transform 1 0 35328 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input197
timestamp 1623621585
transform 1 0 37260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1623621585
transform 1 0 36432 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_392
timestamp 1623621585
transform 1 0 37168 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1623621585
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1623621585
transform 1 0 37904 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_396
timestamp 1623621585
transform 1 0 37536 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1623621585
transform 1 0 38180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1623621585
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1623621585
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1623621585
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1623621585
transform 1 0 3588 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1623621585
transform 1 0 4692 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1623621585
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_51
timestamp 1623621585
transform 1 0 5796 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_58
timestamp 1623621585
transform 1 0 6440 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_70
timestamp 1623621585
transform 1 0 7544 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_82
timestamp 1623621585
transform 1 0 8648 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1623621585
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1623621585
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_106
timestamp 1623621585
transform 1 0 10856 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_115
timestamp 1623621585
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1623621585
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_139
timestamp 1623621585
transform 1 0 13892 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_151
timestamp 1623621585
transform 1 0 14996 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1623621585
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0757_
timestamp 1623621585
transform 1 0 17296 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1623621585
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1623621585
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1623621585
transform 1 0 18032 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1623621585
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_208
timestamp 1623621585
transform 1 0 20240 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1623621585
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1623621585
transform 1 0 21344 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_229
timestamp 1623621585
transform 1 0 22172 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_241
timestamp 1623621585
transform 1 0 23276 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1623621585
transform 1 0 24380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1623621585
transform 1 0 25484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1623621585
transform 1 0 27324 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_277
timestamp 1623621585
transform 1 0 26588 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_286
timestamp 1623621585
transform 1 0 27416 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_298
timestamp 1623621585
transform 1 0 28520 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_310
timestamp 1623621585
transform 1 0 29624 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_322
timestamp 1623621585
transform 1 0 30728 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1623621585
transform 1 0 32568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_334
timestamp 1623621585
transform 1 0 31832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_343
timestamp 1623621585
transform 1 0 32660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_355
timestamp 1623621585
transform 1 0 33764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_367
timestamp 1623621585
transform 1 0 34868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_379
timestamp 1623621585
transform 1 0 35972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_391
timestamp 1623621585
transform 1 0 37076 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1623621585
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1623621585
transform 1 0 37812 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_400
timestamp 1623621585
transform 1 0 37904 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1623621585
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1623621585
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1623621585
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input347
timestamp 1623621585
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input348
timestamp 1623621585
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_6
timestamp 1623621585
transform 1 0 1656 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_18
timestamp 1623621585
transform 1 0 2760 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_6
timestamp 1623621585
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_18
timestamp 1623621585
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1623621585
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_26
timestamp 1623621585
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1623621585
transform 1 0 3864 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1623621585
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1623621585
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1623621585
transform 1 0 4968 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_54
timestamp 1623621585
transform 1 0 6072 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1623621585
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_54
timestamp 1623621585
transform 1 0 6072 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_58
timestamp 1623621585
transform 1 0 6440 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_66
timestamp 1623621585
transform 1 0 7176 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_78
timestamp 1623621585
transform 1 0 8280 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_70
timestamp 1623621585
transform 1 0 7544 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_82
timestamp 1623621585
transform 1 0 8648 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1623621585
transform 1 0 9016 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_87
timestamp 1623621585
transform 1 0 9108 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_99
timestamp 1623621585
transform 1 0 10212 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_94
timestamp 1623621585
transform 1 0 9752 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1623621585
transform 1 0 11592 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_111
timestamp 1623621585
transform 1 0 11316 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1623621585
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_106
timestamp 1623621585
transform 1 0 10856 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_115
timestamp 1623621585
transform 1 0 11684 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1623621585
transform 1 0 14260 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1623621585
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_144
timestamp 1623621585
transform 1 0 14352 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_127
timestamp 1623621585
transform 1 0 12788 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_139
timestamp 1623621585
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1623621585
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_151
timestamp 1623621585
transform 1 0 14996 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_163
timestamp 1623621585
transform 1 0 16100 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0624_
timestamp 1623621585
transform 1 0 17756 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1623621585
transform 1 0 16836 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1623621585
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_180
timestamp 1623621585
transform 1 0 17664 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_172
timestamp 1623621585
transform 1 0 16928 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_180
timestamp 1623621585
transform 1 0 17664 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1623621585
transform 1 0 19504 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_192
timestamp 1623621585
transform 1 0 18768 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_201
timestamp 1623621585
transform 1 0 19596 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_189
timestamp 1623621585
transform 1 0 18492 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1623621585
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0694_
timestamp 1623621585
transform 1 0 20700 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1623621585
transform 1 0 22080 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_213
timestamp 1623621585
transform 1 0 20700 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1623621585
transform 1 0 21804 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_217
timestamp 1623621585
transform 1 0 21068 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_225
timestamp 1623621585
transform 1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_229
timestamp 1623621585
transform 1 0 22172 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23276 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0739_
timestamp 1623621585
transform 1 0 23092 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1623621585
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_247
timestamp 1623621585
transform 1 0 23828 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_249
timestamp 1623621585
transform 1 0 24012 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0747_
timestamp 1623621585
transform 1 0 24380 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1623621585
transform 1 0 24748 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_255
timestamp 1623621585
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_258
timestamp 1623621585
transform 1 0 24840 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_270
timestamp 1623621585
transform 1 0 25944 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_261
timestamp 1623621585
transform 1 0 25116 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1623621585
transform 1 0 27324 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_282
timestamp 1623621585
transform 1 0 27048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_273
timestamp 1623621585
transform 1 0 26220 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_286
timestamp 1623621585
transform 1 0 27416 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_294
timestamp 1623621585
transform 1 0 28152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_306
timestamp 1623621585
transform 1 0 29256 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_298
timestamp 1623621585
transform 1 0 28520 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_310
timestamp 1623621585
transform 1 0 29624 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1623621585
transform 1 0 29992 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_315
timestamp 1623621585
transform 1 0 30084 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_327
timestamp 1623621585
transform 1 0 31188 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_322
timestamp 1623621585
transform 1 0 30728 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1623621585
transform 1 0 32568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_339
timestamp 1623621585
transform 1 0 32292 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_351
timestamp 1623621585
transform 1 0 33396 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_334
timestamp 1623621585
transform 1 0 31832 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_343
timestamp 1623621585
transform 1 0 32660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1623621585
transform 1 0 35236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_363
timestamp 1623621585
transform 1 0 34500 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_372
timestamp 1623621585
transform 1 0 35328 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_355
timestamp 1623621585
transform 1 0 33764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_367
timestamp 1623621585
transform 1 0 34868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input198
timestamp 1623621585
transform 1 0 37260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1623621585
transform 1 0 36432 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_392
timestamp 1623621585
transform 1 0 37168 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_379
timestamp 1623621585
transform 1 0 35972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_391
timestamp 1623621585
transform 1 0 37076 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1623621585
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1623621585
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1623621585
transform 1 0 37812 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1623621585
transform 1 0 37904 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_396
timestamp 1623621585
transform 1 0 37536 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1623621585
transform 1 0 38180 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_400
timestamp 1623621585
transform 1 0 37904 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1623621585
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1623621585
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1623621585
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1623621585
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1623621585
transform 1 0 3772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_27
timestamp 1623621585
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_30
timestamp 1623621585
transform 1 0 3864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_42
timestamp 1623621585
transform 1 0 4968 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_54
timestamp 1623621585
transform 1 0 6072 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_66
timestamp 1623621585
transform 1 0 7176 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_78
timestamp 1623621585
transform 1 0 8280 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1623621585
transform 1 0 9016 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_87
timestamp 1623621585
transform 1 0 9108 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_99
timestamp 1623621585
transform 1 0 10212 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_111
timestamp 1623621585
transform 1 0 11316 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1623621585
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1623621585
transform 1 0 14260 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1623621585
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_144
timestamp 1623621585
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1623621585
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0616_
timestamp 1623621585
transform 1 0 17848 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1623621585
transform 1 0 16744 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_168
timestamp 1623621585
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1623621585
transform 1 0 17480 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0695_
timestamp 1623621585
transform 1 0 20056 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1623621585
transform 1 0 19504 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_190
timestamp 1623621585
transform 1 0 18584 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1623621585
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_201
timestamp 1623621585
transform 1 0 19596 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_205
timestamp 1623621585
transform 1 0 19964 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _0989_
timestamp 1623621585
transform 1 0 20792 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_35_210
timestamp 1623621585
transform 1 0 20424 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0990_
timestamp 1623621585
transform 1 0 22724 0 1 21216
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1623621585
transform 1 0 22356 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1623621585
transform 1 0 24748 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_252
timestamp 1623621585
transform 1 0 24288 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_256
timestamp 1623621585
transform 1 0 24656 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_258
timestamp 1623621585
transform 1 0 24840 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_270
timestamp 1623621585
transform 1 0 25944 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_282
timestamp 1623621585
transform 1 0 27048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_294
timestamp 1623621585
transform 1 0 28152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 1623621585
transform 1 0 29256 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1623621585
transform 1 0 29992 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_315
timestamp 1623621585
transform 1 0 30084 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_327
timestamp 1623621585
transform 1 0 31188 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_339
timestamp 1623621585
transform 1 0 32292 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_351
timestamp 1623621585
transform 1 0 33396 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1623621585
transform 1 0 35236 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_363
timestamp 1623621585
transform 1 0 34500 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_372
timestamp 1623621585
transform 1 0 35328 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1623621585
transform 1 0 37260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_384
timestamp 1623621585
transform 1 0 36432 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_392
timestamp 1623621585
transform 1 0 37168 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1623621585
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1623621585
transform 1 0 37904 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_396
timestamp 1623621585
transform 1 0 37536 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1623621585
transform 1 0 38180 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1623621585
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input349
timestamp 1623621585
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_6
timestamp 1623621585
transform 1 0 1656 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_18
timestamp 1623621585
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1623621585
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1623621585
transform 1 0 6348 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1623621585
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_54
timestamp 1623621585
transform 1 0 6072 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_58
timestamp 1623621585
transform 1 0 6440 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1623621585
transform 1 0 7544 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_82
timestamp 1623621585
transform 1 0 8648 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_94
timestamp 1623621585
transform 1 0 9752 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1623621585
transform 1 0 11592 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_106
timestamp 1623621585
transform 1 0 10856 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_115
timestamp 1623621585
transform 1 0 11684 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1623621585
transform 1 0 12788 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_139
timestamp 1623621585
transform 1 0 13892 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_151
timestamp 1623621585
transform 1 0 14996 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_163
timestamp 1623621585
transform 1 0 16100 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_4  _0779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 17388 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1623621585
transform 1 0 16836 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_172
timestamp 1623621585
transform 1 0 16928 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_176
timestamp 1623621585
transform 1 0 17296 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1623621585
transform 1 0 18216 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0608_
timestamp 1623621585
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1017_
timestamp 1623621585
transform 1 0 20148 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_36_198
timestamp 1623621585
transform 1 0 19320 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_206
timestamp 1623621585
transform 1 0 20056 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1623621585
transform 1 0 22080 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_224
timestamp 1623621585
transform 1 0 21712 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1623621585
transform 1 0 22172 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0992_
timestamp 1623621585
transform 1 0 22540 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_36_250
timestamp 1623621585
transform 1 0 24104 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0722_
timestamp 1623621585
transform 1 0 24472 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_262
timestamp 1623621585
transform 1 0 25208 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1623621585
transform 1 0 27324 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_274
timestamp 1623621585
transform 1 0 26312 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_282
timestamp 1623621585
transform 1 0 27048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_286
timestamp 1623621585
transform 1 0 27416 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_298
timestamp 1623621585
transform 1 0 28520 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_310
timestamp 1623621585
transform 1 0 29624 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_322
timestamp 1623621585
transform 1 0 30728 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1623621585
transform 1 0 32568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_334
timestamp 1623621585
transform 1 0 31832 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_343
timestamp 1623621585
transform 1 0 32660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_355
timestamp 1623621585
transform 1 0 33764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_367
timestamp 1623621585
transform 1 0 34868 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input199
timestamp 1623621585
transform 1 0 37168 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_379
timestamp 1623621585
transform 1 0 35972 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_391
timestamp 1623621585
transform 1 0 37076 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_395
timestamp 1623621585
transform 1 0 37444 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1623621585
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1623621585
transform 1 0 37812 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_400
timestamp 1623621585
transform 1 0 37904 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1623621585
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1623621585
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input350
timestamp 1623621585
transform 1 0 1380 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_6
timestamp 1623621585
transform 1 0 1656 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_18
timestamp 1623621585
transform 1 0 2760 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1623621585
transform 1 0 3772 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_26
timestamp 1623621585
transform 1 0 3496 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1623621585
transform 1 0 3864 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1623621585
transform 1 0 4968 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_54
timestamp 1623621585
transform 1 0 6072 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_66
timestamp 1623621585
transform 1 0 7176 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_78
timestamp 1623621585
transform 1 0 8280 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1623621585
transform 1 0 9016 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_87
timestamp 1623621585
transform 1 0 9108 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_99
timestamp 1623621585
transform 1 0 10212 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_111
timestamp 1623621585
transform 1 0 11316 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1623621585
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1623621585
transform 1 0 14260 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1623621585
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_144
timestamp 1623621585
transform 1 0 14352 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_156
timestamp 1623621585
transform 1 0 15456 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0590_
timestamp 1623621585
transform 1 0 17940 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_168
timestamp 1623621585
transform 1 0 16560 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_180
timestamp 1623621585
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1623621585
transform 1 0 19504 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_191
timestamp 1623621585
transform 1 0 18676 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_199
timestamp 1623621585
transform 1 0 19412 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1623621585
transform 1 0 19596 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _0991_
timestamp 1623621585
transform 1 0 21344 0 1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_37_213
timestamp 1623621585
transform 1 0 20700 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_219
timestamp 1623621585
transform 1 0 21252 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _0714_
timestamp 1623621585
transform 1 0 23552 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_237
timestamp 1623621585
transform 1 0 22908 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1623621585
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1623621585
transform 1 0 24748 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_252
timestamp 1623621585
transform 1 0 24288 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_256
timestamp 1623621585
transform 1 0 24656 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_258
timestamp 1623621585
transform 1 0 24840 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_270
timestamp 1623621585
transform 1 0 25944 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_282
timestamp 1623621585
transform 1 0 27048 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_294
timestamp 1623621585
transform 1 0 28152 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_306
timestamp 1623621585
transform 1 0 29256 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1623621585
transform 1 0 29992 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_315
timestamp 1623621585
transform 1 0 30084 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_327
timestamp 1623621585
transform 1 0 31188 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_339
timestamp 1623621585
transform 1 0 32292 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_351
timestamp 1623621585
transform 1 0 33396 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1623621585
transform 1 0 35236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_363
timestamp 1623621585
transform 1 0 34500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_372
timestamp 1623621585
transform 1 0 35328 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1623621585
transform 1 0 37260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1623621585
transform 1 0 36432 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_392
timestamp 1623621585
transform 1 0 37168 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1623621585
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1623621585
transform 1 0 37904 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_396
timestamp 1623621585
transform 1 0 37536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1623621585
transform 1 0 38180 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1623621585
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1623621585
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1623621585
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_27
timestamp 1623621585
transform 1 0 3588 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_39
timestamp 1623621585
transform 1 0 4692 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1623621585
transform 1 0 6348 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_51
timestamp 1623621585
transform 1 0 5796 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_58
timestamp 1623621585
transform 1 0 6440 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_70
timestamp 1623621585
transform 1 0 7544 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_82
timestamp 1623621585
transform 1 0 8648 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_94
timestamp 1623621585
transform 1 0 9752 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1623621585
transform 1 0 11592 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_106
timestamp 1623621585
transform 1 0 10856 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_115
timestamp 1623621585
transform 1 0 11684 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_127
timestamp 1623621585
transform 1 0 12788 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_139
timestamp 1623621585
transform 1 0 13892 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_151
timestamp 1623621585
transform 1 0 14996 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_163
timestamp 1623621585
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0532_
timestamp 1623621585
transform 1 0 18124 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0533_
timestamp 1623621585
transform 1 0 17480 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1623621585
transform 1 0 16836 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_172
timestamp 1623621585
transform 1 0 16928 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1623621585
transform 1 0 17756 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0982_
timestamp 1623621585
transform 1 0 18768 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_38_188
timestamp 1623621585
transform 1 0 18400 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0640_
timestamp 1623621585
transform 1 0 21068 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1623621585
transform 1 0 22080 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_209
timestamp 1623621585
transform 1 0 20332 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_221
timestamp 1623621585
transform 1 0 21436 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_227
timestamp 1623621585
transform 1 0 21988 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_229
timestamp 1623621585
transform 1 0 22172 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0993_
timestamp 1623621585
transform 1 0 22540 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_38_250
timestamp 1623621585
transform 1 0 24104 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_262
timestamp 1623621585
transform 1 0 25208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1623621585
transform 1 0 27324 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_274
timestamp 1623621585
transform 1 0 26312 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_282
timestamp 1623621585
transform 1 0 27048 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_286
timestamp 1623621585
transform 1 0 27416 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_298
timestamp 1623621585
transform 1 0 28520 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_310
timestamp 1623621585
transform 1 0 29624 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_322
timestamp 1623621585
transform 1 0 30728 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1623621585
transform 1 0 32568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_334
timestamp 1623621585
transform 1 0 31832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_343
timestamp 1623621585
transform 1 0 32660 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_355
timestamp 1623621585
transform 1 0 33764 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_367
timestamp 1623621585
transform 1 0 34868 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input200
timestamp 1623621585
transform 1 0 37168 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_379
timestamp 1623621585
transform 1 0 35972 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_391
timestamp 1623621585
transform 1 0 37076 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_395
timestamp 1623621585
transform 1 0 37444 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1623621585
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1623621585
transform 1 0 37812 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_400
timestamp 1623621585
transform 1 0 37904 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1623621585
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1623621585
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1623621585
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input351
timestamp 1623621585
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input352
timestamp 1623621585
transform 1 0 1748 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1623621585
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1623621585
transform 1 0 2116 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1623621585
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_11
timestamp 1623621585
transform 1 0 2116 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1623621585
transform 1 0 3772 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_23
timestamp 1623621585
transform 1 0 3220 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_30
timestamp 1623621585
transform 1 0 3864 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_23
timestamp 1623621585
transform 1 0 3220 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_35
timestamp 1623621585
transform 1 0 4324 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1623621585
transform 1 0 6348 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_42
timestamp 1623621585
transform 1 0 4968 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_54
timestamp 1623621585
transform 1 0 6072 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_47
timestamp 1623621585
transform 1 0 5428 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_55
timestamp 1623621585
transform 1 0 6164 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_58
timestamp 1623621585
transform 1 0 6440 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_66
timestamp 1623621585
transform 1 0 7176 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_78
timestamp 1623621585
transform 1 0 8280 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_70
timestamp 1623621585
transform 1 0 7544 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_82
timestamp 1623621585
transform 1 0 8648 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1623621585
transform 1 0 9016 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_87
timestamp 1623621585
transform 1 0 9108 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_99
timestamp 1623621585
transform 1 0 10212 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_94
timestamp 1623621585
transform 1 0 9752 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1623621585
transform 1 0 11592 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_111
timestamp 1623621585
transform 1 0 11316 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1623621585
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_106
timestamp 1623621585
transform 1 0 10856 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_115
timestamp 1623621585
transform 1 0 11684 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1623621585
transform 1 0 14260 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1623621585
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_144
timestamp 1623621585
transform 1 0 14352 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_127
timestamp 1623621585
transform 1 0 12788 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_139
timestamp 1623621585
transform 1 0 13892 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_156
timestamp 1623621585
transform 1 0 15456 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_151
timestamp 1623621585
transform 1 0 14996 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_163
timestamp 1623621585
transform 1 0 16100 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0570_
timestamp 1623621585
transform 1 0 17480 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1623621585
transform 1 0 16836 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_168
timestamp 1623621585
transform 1 0 16560 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_180
timestamp 1623621585
transform 1 0 17664 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_172
timestamp 1623621585
transform 1 0 16928 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_186
timestamp 1623621585
transform 1 0 18216 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0466_
timestamp 1623621585
transform 1 0 18492 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1623621585
transform 1 0 19964 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0981_
timestamp 1623621585
transform 1 0 18584 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1623621585
transform 1 0 19504 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_188
timestamp 1623621585
transform 1 0 18400 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_192
timestamp 1623621585
transform 1 0 18768 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_201
timestamp 1623621585
transform 1 0 19596 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_208
timestamp 1623621585
transform 1 0 20240 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_207
timestamp 1623621585
transform 1 0 20148 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0587_
timestamp 1623621585
transform 1 0 21344 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0641_
timestamp 1623621585
transform 1 0 21252 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1623621585
transform 1 0 22080 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1623621585
transform 1 0 21988 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_216
timestamp 1623621585
transform 1 0 20976 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_223
timestamp 1623621585
transform 1 0 21620 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_219
timestamp 1623621585
transform 1 0 21252 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1623621585
transform 1 0 21712 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1623621585
transform 1 0 22172 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_230
timestamp 1623621585
transform 1 0 22264 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_242
timestamp 1623621585
transform 1 0 23368 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_241
timestamp 1623621585
transform 1 0 23276 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1623621585
transform 1 0 24748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1623621585
transform 1 0 24472 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_254
timestamp 1623621585
transform 1 0 24472 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_258
timestamp 1623621585
transform 1 0 24840 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_270
timestamp 1623621585
transform 1 0 25944 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1623621585
transform 1 0 24380 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_257
timestamp 1623621585
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_269
timestamp 1623621585
transform 1 0 25852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1623621585
transform 1 0 27324 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_282
timestamp 1623621585
transform 1 0 27048 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_281
timestamp 1623621585
transform 1 0 26956 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_286
timestamp 1623621585
transform 1 0 27416 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_294
timestamp 1623621585
transform 1 0 28152 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_306
timestamp 1623621585
transform 1 0 29256 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_298
timestamp 1623621585
transform 1 0 28520 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_310
timestamp 1623621585
transform 1 0 29624 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1623621585
transform 1 0 29992 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_315
timestamp 1623621585
transform 1 0 30084 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_327
timestamp 1623621585
transform 1 0 31188 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_322
timestamp 1623621585
transform 1 0 30728 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1623621585
transform 1 0 32568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_339
timestamp 1623621585
transform 1 0 32292 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_351
timestamp 1623621585
transform 1 0 33396 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_334
timestamp 1623621585
transform 1 0 31832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_343
timestamp 1623621585
transform 1 0 32660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1623621585
transform 1 0 35236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_363
timestamp 1623621585
transform 1 0 34500 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_372
timestamp 1623621585
transform 1 0 35328 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_355
timestamp 1623621585
transform 1 0 33764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_367
timestamp 1623621585
transform 1 0 34868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input168
timestamp 1623621585
transform 1 0 37260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input201
timestamp 1623621585
transform 1 0 37168 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 1623621585
transform 1 0 36432 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_392
timestamp 1623621585
transform 1 0 37168 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_379
timestamp 1623621585
transform 1 0 35972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_391
timestamp 1623621585
transform 1 0 37076 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_395
timestamp 1623621585
transform 1 0 37444 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1623621585
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1623621585
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1623621585
transform 1 0 37812 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1623621585
transform 1 0 37904 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1623621585
transform 1 0 37536 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1623621585
transform 1 0 38180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_400
timestamp 1623621585
transform 1 0 37904 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1623621585
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1623621585
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1623621585
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1623621585
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1623621585
transform 1 0 3772 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_27
timestamp 1623621585
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1623621585
transform 1 0 3864 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1623621585
transform 1 0 4968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_54
timestamp 1623621585
transform 1 0 6072 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_66
timestamp 1623621585
transform 1 0 7176 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_78
timestamp 1623621585
transform 1 0 8280 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1623621585
transform 1 0 9016 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_87
timestamp 1623621585
transform 1 0 9108 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1623621585
transform 1 0 10212 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_111
timestamp 1623621585
transform 1 0 11316 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1623621585
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1623621585
transform 1 0 14260 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1623621585
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_144
timestamp 1623621585
transform 1 0 14352 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1623621585
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0562_
timestamp 1623621585
transform 1 0 17940 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0579_
timestamp 1623621585
transform 1 0 16836 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_168
timestamp 1623621585
transform 1 0 16560 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1623621585
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0468_
timestamp 1623621585
transform 1 0 19964 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1623621585
transform 1 0 19504 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_191
timestamp 1623621585
transform 1 0 18676 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_199
timestamp 1623621585
transform 1 0 19412 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1623621585
transform 1 0 19596 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0465_
timestamp 1623621585
transform 1 0 21804 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20976 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_41_209
timestamp 1623621585
transform 1 0 20332 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_215
timestamp 1623621585
transform 1 0 20884 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_221
timestamp 1623621585
transform 1 0 21436 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_229
timestamp 1623621585
transform 1 0 22172 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0586_
timestamp 1623621585
transform 1 0 22540 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0693_
timestamp 1623621585
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1623621585
transform 1 0 22908 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0676_
timestamp 1623621585
transform 1 0 25208 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1623621585
transform 1 0 24748 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_253
timestamp 1623621585
transform 1 0 24380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_258
timestamp 1623621585
transform 1 0 24840 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_270
timestamp 1623621585
transform 1 0 25944 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_282
timestamp 1623621585
transform 1 0 27048 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_294
timestamp 1623621585
transform 1 0 28152 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_306
timestamp 1623621585
transform 1 0 29256 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1623621585
transform 1 0 29992 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_315
timestamp 1623621585
transform 1 0 30084 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_327
timestamp 1623621585
transform 1 0 31188 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_339
timestamp 1623621585
transform 1 0 32292 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_351
timestamp 1623621585
transform 1 0 33396 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1623621585
transform 1 0 35236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_363
timestamp 1623621585
transform 1 0 34500 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_372
timestamp 1623621585
transform 1 0 35328 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_384
timestamp 1623621585
transform 1 0 36432 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1623621585
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1623621585
transform 1 0 37904 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_396
timestamp 1623621585
transform 1 0 37536 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1623621585
transform 1 0 38180 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1623621585
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input354
timestamp 1623621585
transform 1 0 1748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1623621585
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_11
timestamp 1623621585
transform 1 0 2116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_23
timestamp 1623621585
transform 1 0 3220 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_35
timestamp 1623621585
transform 1 0 4324 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1623621585
transform 1 0 6348 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_47
timestamp 1623621585
transform 1 0 5428 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_55
timestamp 1623621585
transform 1 0 6164 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_58
timestamp 1623621585
transform 1 0 6440 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_70
timestamp 1623621585
transform 1 0 7544 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_82
timestamp 1623621585
transform 1 0 8648 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1623621585
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1623621585
transform 1 0 11592 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 1623621585
transform 1 0 10856 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_115
timestamp 1623621585
transform 1 0 11684 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_127
timestamp 1623621585
transform 1 0 12788 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_139
timestamp 1623621585
transform 1 0 13892 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_151
timestamp 1623621585
transform 1 0 14996 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_163
timestamp 1623621585
transform 1 0 16100 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0554_
timestamp 1623621585
transform 1 0 17848 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1623621585
transform 1 0 16836 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_172
timestamp 1623621585
transform 1 0 16928 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_180
timestamp 1623621585
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _0983_
timestamp 1623621585
transform 1 0 18952 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_42_190
timestamp 1623621585
transform 1 0 18584 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0467_
timestamp 1623621585
transform 1 0 21252 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1623621585
transform 1 0 22080 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_211
timestamp 1623621585
transform 1 0 20516 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1623621585
transform 1 0 21620 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_227
timestamp 1623621585
transform 1 0 21988 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_229
timestamp 1623621585
transform 1 0 22172 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _0994_
timestamp 1623621585
transform 1 0 22540 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_42_250
timestamp 1623621585
transform 1 0 24104 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0660_
timestamp 1623621585
transform 1 0 24748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0685_
timestamp 1623621585
transform 1 0 25852 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_256
timestamp 1623621585
transform 1 0 24656 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1623621585
transform 1 0 25484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1623621585
transform 1 0 27324 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1623621585
transform 1 0 26588 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_286
timestamp 1623621585
transform 1 0 27416 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_298
timestamp 1623621585
transform 1 0 28520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_310
timestamp 1623621585
transform 1 0 29624 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_322
timestamp 1623621585
transform 1 0 30728 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1623621585
transform 1 0 32568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_334
timestamp 1623621585
transform 1 0 31832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_343
timestamp 1623621585
transform 1 0 32660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_355
timestamp 1623621585
transform 1 0 33764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_367
timestamp 1623621585
transform 1 0 34868 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1623621585
transform 1 0 37168 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_379
timestamp 1623621585
transform 1 0 35972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_391
timestamp 1623621585
transform 1 0 37076 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_395
timestamp 1623621585
transform 1 0 37444 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1623621585
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1623621585
transform 1 0 37812 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_400
timestamp 1623621585
transform 1 0 37904 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1623621585
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1623621585
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input355
timestamp 1623621585
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1623621585
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_11
timestamp 1623621585
transform 1 0 2116 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1623621585
transform 1 0 3772 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_23
timestamp 1623621585
transform 1 0 3220 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_30
timestamp 1623621585
transform 1 0 3864 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_42
timestamp 1623621585
transform 1 0 4968 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_54
timestamp 1623621585
transform 1 0 6072 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_66
timestamp 1623621585
transform 1 0 7176 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_78
timestamp 1623621585
transform 1 0 8280 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1623621585
transform 1 0 9016 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_87
timestamp 1623621585
transform 1 0 9108 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1623621585
transform 1 0 10212 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_111
timestamp 1623621585
transform 1 0 11316 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1623621585
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1623621585
transform 1 0 14260 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1623621585
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_144
timestamp 1623621585
transform 1 0 14352 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_156
timestamp 1623621585
transform 1 0 15456 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0536_
timestamp 1623621585
transform 1 0 18032 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_168
timestamp 1623621585
transform 1 0 16560 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_180
timestamp 1623621585
transform 1 0 17664 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1623621585
transform 1 0 19504 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_192
timestamp 1623621585
transform 1 0 18768 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1623621585
transform 1 0 19596 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 20884 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_43_213
timestamp 1623621585
transform 1 0 20700 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_2  _0995_
timestamp 1623621585
transform 1 0 22816 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_43_231
timestamp 1623621585
transform 1 0 22356 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_235
timestamp 1623621585
transform 1 0 22724 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1623621585
transform 1 0 25208 0 1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1623621585
transform 1 0 24748 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_253
timestamp 1623621585
transform 1 0 24380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_258
timestamp 1623621585
transform 1 0 24840 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_279
timestamp 1623621585
transform 1 0 26772 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_291
timestamp 1623621585
transform 1 0 27876 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_303
timestamp 1623621585
transform 1 0 28980 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_311
timestamp 1623621585
transform 1 0 29716 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1623621585
transform 1 0 29992 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_315
timestamp 1623621585
transform 1 0 30084 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_327
timestamp 1623621585
transform 1 0 31188 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_339
timestamp 1623621585
transform 1 0 32292 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_351
timestamp 1623621585
transform 1 0 33396 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1623621585
transform 1 0 35236 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_363
timestamp 1623621585
transform 1 0 34500 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_372
timestamp 1623621585
transform 1 0 35328 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input202
timestamp 1623621585
transform 1 0 37260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_384
timestamp 1623621585
transform 1 0 36432 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_392
timestamp 1623621585
transform 1 0 37168 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1623621585
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1623621585
transform 1 0 37904 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_396
timestamp 1623621585
transform 1 0 37536 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1623621585
transform 1 0 38180 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1623621585
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1623621585
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1623621585
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_27
timestamp 1623621585
transform 1 0 3588 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_39
timestamp 1623621585
transform 1 0 4692 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1623621585
transform 1 0 6348 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_51
timestamp 1623621585
transform 1 0 5796 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_58
timestamp 1623621585
transform 1 0 6440 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_70
timestamp 1623621585
transform 1 0 7544 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_82
timestamp 1623621585
transform 1 0 8648 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_94
timestamp 1623621585
transform 1 0 9752 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1623621585
transform 1 0 11592 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_106
timestamp 1623621585
transform 1 0 10856 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_115
timestamp 1623621585
transform 1 0 11684 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_127
timestamp 1623621585
transform 1 0 12788 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_139
timestamp 1623621585
transform 1 0 13892 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_151
timestamp 1623621585
transform 1 0 14996 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_163
timestamp 1623621585
transform 1 0 16100 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1623621585
transform 1 0 16836 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_172
timestamp 1623621585
transform 1 0 16928 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_184
timestamp 1623621585
transform 1 0 18032 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0972_
timestamp 1623621585
transform 1 0 18676 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 18492 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 1623621585
transform 1 0 18400 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_207
timestamp 1623621585
transform 1 0 20148 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0415_
timestamp 1623621585
transform 1 0 20608 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1623621585
transform 1 0 22080 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_211
timestamp 1623621585
transform 1 0 20516 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_221
timestamp 1623621585
transform 1 0 21436 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1623621585
transform 1 0 21988 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_229
timestamp 1623621585
transform 1 0 22172 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1623621585
transform 1 0 23184 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_44_237
timestamp 1623621585
transform 1 0 22908 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1623621585
transform 1 0 25116 0 -1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_44_257
timestamp 1623621585
transform 1 0 24748 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1623621585
transform 1 0 27324 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_278
timestamp 1623621585
transform 1 0 26680 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_284
timestamp 1623621585
transform 1 0 27232 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_286
timestamp 1623621585
transform 1 0 27416 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_298
timestamp 1623621585
transform 1 0 28520 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_310
timestamp 1623621585
transform 1 0 29624 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_322
timestamp 1623621585
transform 1 0 30728 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1623621585
transform 1 0 32568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_334
timestamp 1623621585
transform 1 0 31832 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_343
timestamp 1623621585
transform 1 0 32660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_355
timestamp 1623621585
transform 1 0 33764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_367
timestamp 1623621585
transform 1 0 34868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_379
timestamp 1623621585
transform 1 0 35972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_391
timestamp 1623621585
transform 1 0 37076 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1623621585
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1623621585
transform 1 0 37812 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_400
timestamp 1623621585
transform 1 0 37904 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1623621585
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1623621585
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input363
timestamp 1623621585
transform 1 0 1748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1623621585
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_11
timestamp 1623621585
transform 1 0 2116 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1623621585
transform 1 0 3772 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_23
timestamp 1623621585
transform 1 0 3220 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_30
timestamp 1623621585
transform 1 0 3864 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_42
timestamp 1623621585
transform 1 0 4968 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_54
timestamp 1623621585
transform 1 0 6072 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_66
timestamp 1623621585
transform 1 0 7176 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_78
timestamp 1623621585
transform 1 0 8280 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1623621585
transform 1 0 9016 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_87
timestamp 1623621585
transform 1 0 9108 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_99
timestamp 1623621585
transform 1 0 10212 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_111
timestamp 1623621585
transform 1 0 11316 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1623621585
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1623621585
transform 1 0 14260 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1623621585
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_144
timestamp 1623621585
transform 1 0 14352 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_156
timestamp 1623621585
transform 1 0 15456 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_168
timestamp 1623621585
transform 1 0 16560 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_180
timestamp 1623621585
transform 1 0 17664 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0973_
timestamp 1623621585
transform 1 0 19964 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1623621585
transform 1 0 19504 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_192
timestamp 1623621585
transform 1 0 18768 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_201
timestamp 1623621585
transform 1 0 19596 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0974_
timestamp 1623621585
transform 1 0 21804 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_221
timestamp 1623621585
transform 1 0 21436 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0713_
timestamp 1623621585
transform 1 0 24012 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_241
timestamp 1623621585
transform 1 0 23276 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0668_
timestamp 1623621585
transform 1 0 25208 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1623621585
transform 1 0 24748 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_253
timestamp 1623621585
transform 1 0 24380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_258
timestamp 1623621585
transform 1 0 24840 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_270
timestamp 1623621585
transform 1 0 25944 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_282
timestamp 1623621585
transform 1 0 27048 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_294
timestamp 1623621585
transform 1 0 28152 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_306
timestamp 1623621585
transform 1 0 29256 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1623621585
transform 1 0 29992 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_315
timestamp 1623621585
transform 1 0 30084 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_327
timestamp 1623621585
transform 1 0 31188 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_339
timestamp 1623621585
transform 1 0 32292 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_351
timestamp 1623621585
transform 1 0 33396 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1623621585
transform 1 0 35236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_363
timestamp 1623621585
transform 1 0 34500 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_372
timestamp 1623621585
transform 1 0 35328 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1623621585
transform 1 0 37260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_384
timestamp 1623621585
transform 1 0 36432 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_392
timestamp 1623621585
transform 1 0 37168 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1623621585
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1623621585
transform 1 0 37904 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_396
timestamp 1623621585
transform 1 0 37536 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1623621585
transform 1 0 38180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1623621585
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1623621585
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input374
timestamp 1623621585
transform 1 0 1748 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1623621585
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_11
timestamp 1623621585
transform 1 0 2116 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1623621585
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1623621585
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1623621585
transform 1 0 3772 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_23
timestamp 1623621585
transform 1 0 3220 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_35
timestamp 1623621585
transform 1 0 4324 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_27
timestamp 1623621585
transform 1 0 3588 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_30
timestamp 1623621585
transform 1 0 3864 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1623621585
transform 1 0 6348 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_47
timestamp 1623621585
transform 1 0 5428 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_55
timestamp 1623621585
transform 1 0 6164 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_58
timestamp 1623621585
transform 1 0 6440 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_42
timestamp 1623621585
transform 1 0 4968 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_54
timestamp 1623621585
transform 1 0 6072 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_70
timestamp 1623621585
transform 1 0 7544 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_82
timestamp 1623621585
transform 1 0 8648 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_66
timestamp 1623621585
transform 1 0 7176 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1623621585
transform 1 0 8280 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1623621585
transform 1 0 9016 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_94
timestamp 1623621585
transform 1 0 9752 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_87
timestamp 1623621585
transform 1 0 9108 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_99
timestamp 1623621585
transform 1 0 10212 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1623621585
transform 1 0 11592 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_106
timestamp 1623621585
transform 1 0 10856 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_115
timestamp 1623621585
transform 1 0 11684 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_111
timestamp 1623621585
transform 1 0 11316 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1623621585
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1623621585
transform 1 0 14260 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_127
timestamp 1623621585
transform 1 0 12788 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_139
timestamp 1623621585
transform 1 0 13892 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1623621585
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_144
timestamp 1623621585
transform 1 0 14352 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_151
timestamp 1623621585
transform 1 0 14996 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_163
timestamp 1623621585
transform 1 0 16100 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_156
timestamp 1623621585
transform 1 0 15456 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1623621585
transform 1 0 16836 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_172
timestamp 1623621585
transform 1 0 16928 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_184
timestamp 1623621585
transform 1 0 18032 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_168
timestamp 1623621585
transform 1 0 16560 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_180
timestamp 1623621585
transform 1 0 17664 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0416_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 19412 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0525_
timestamp 1623621585
transform 1 0 18400 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _0976_
timestamp 1623621585
transform 1 0 20240 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1623621585
transform 1 0 19504 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_196
timestamp 1623621585
transform 1 0 19136 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_204
timestamp 1623621585
transform 1 0 19872 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1623621585
transform 1 0 19136 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_201
timestamp 1623621585
transform 1 0 19596 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _0975_
timestamp 1623621585
transform 1 0 20976 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1623621585
transform 1 0 22080 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1623621585
transform 1 0 21712 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_229
timestamp 1623621585
transform 1 0 22172 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_213
timestamp 1623621585
transform 1 0 20700 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1623621585
transform 1 0 22540 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1623621585
transform 1 0 22816 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_46_249
timestamp 1623621585
transform 1 0 24012 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_232
timestamp 1623621585
transform 1 0 22448 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0417_
timestamp 1623621585
transform 1 0 24380 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _0622_
timestamp 1623621585
transform 1 0 25760 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0639_
timestamp 1623621585
transform 1 0 25576 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1623621585
transform 1 0 24748 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_262
timestamp 1623621585
transform 1 0 25208 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1623621585
transform 1 0 24288 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_256
timestamp 1623621585
transform 1 0 24656 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_258
timestamp 1623621585
transform 1 0 24840 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_266
timestamp 1623621585
transform 1 0 25576 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0659_
timestamp 1623621585
transform 1 0 26680 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0763_
timestamp 1623621585
transform 1 0 26864 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1623621585
transform 1 0 27324 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_274
timestamp 1623621585
transform 1 0 26312 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_281
timestamp 1623621585
transform 1 0 26956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_286
timestamp 1623621585
transform 1 0 27416 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1623621585
transform 1 0 26496 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_288
timestamp 1623621585
transform 1 0 27600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_298
timestamp 1623621585
transform 1 0 28520 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_310
timestamp 1623621585
transform 1 0 29624 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_300
timestamp 1623621585
transform 1 0 28704 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_312
timestamp 1623621585
transform 1 0 29808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1623621585
transform 1 0 29992 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_322
timestamp 1623621585
transform 1 0 30728 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_315
timestamp 1623621585
transform 1 0 30084 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_327
timestamp 1623621585
transform 1 0 31188 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1623621585
transform 1 0 32568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_334
timestamp 1623621585
transform 1 0 31832 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_343
timestamp 1623621585
transform 1 0 32660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_339
timestamp 1623621585
transform 1 0 32292 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_351
timestamp 1623621585
transform 1 0 33396 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1623621585
transform 1 0 35236 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_355
timestamp 1623621585
transform 1 0 33764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_367
timestamp 1623621585
transform 1 0 34868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_363
timestamp 1623621585
transform 1 0 34500 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_372
timestamp 1623621585
transform 1 0 35328 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0699_
timestamp 1623621585
transform 1 0 35972 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0743_
timestamp 1623621585
transform 1 0 35880 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1623621585
transform 1 0 37260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_382
timestamp 1623621585
transform 1 0 36248 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_394
timestamp 1623621585
transform 1 0 37352 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_386
timestamp 1623621585
transform 1 0 36616 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_392
timestamp 1623621585
transform 1 0 37168 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1623621585
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1623621585
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1623621585
transform 1 0 37812 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1623621585
transform 1 0 37904 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_398
timestamp 1623621585
transform 1 0 37720 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_400
timestamp 1623621585
transform 1 0 37904 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1623621585
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1623621585
transform 1 0 37536 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1623621585
transform 1 0 38180 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1623621585
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input385 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 1380 0 -1 28832
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_48_13
timestamp 1623621585
transform 1 0 2300 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_25
timestamp 1623621585
transform 1 0 3404 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_37
timestamp 1623621585
transform 1 0 4508 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1623621585
transform 1 0 6348 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_49
timestamp 1623621585
transform 1 0 5612 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_58
timestamp 1623621585
transform 1 0 6440 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_70
timestamp 1623621585
transform 1 0 7544 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_82
timestamp 1623621585
transform 1 0 8648 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_94
timestamp 1623621585
transform 1 0 9752 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1623621585
transform 1 0 11592 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_106
timestamp 1623621585
transform 1 0 10856 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_115
timestamp 1623621585
transform 1 0 11684 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_127
timestamp 1623621585
transform 1 0 12788 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_139
timestamp 1623621585
transform 1 0 13892 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_151
timestamp 1623621585
transform 1 0 14996 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_163
timestamp 1623621585
transform 1 0 16100 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1623621585
transform 1 0 16836 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_172
timestamp 1623621585
transform 1 0 16928 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_184
timestamp 1623621585
transform 1 0 18032 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0508_
timestamp 1623621585
transform 1 0 18676 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0516_
timestamp 1623621585
transform 1 0 19780 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_190
timestamp 1623621585
transform 1 0 18584 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_199
timestamp 1623621585
transform 1 0 19412 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1623621585
transform 1 0 22080 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_211
timestamp 1623621585
transform 1 0 20516 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1623621585
transform 1 0 21620 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_227
timestamp 1623621585
transform 1 0 21988 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_229
timestamp 1623621585
transform 1 0 22172 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1623621585
transform 1 0 22540 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_48_249
timestamp 1623621585
transform 1 0 24012 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1001_
timestamp 1623621585
transform 1 0 25208 0 -1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1623621585
transform 1 0 25116 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1623621585
transform 1 0 27324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_279
timestamp 1623621585
transform 1 0 26772 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_286
timestamp 1623621585
transform 1 0 27416 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_298
timestamp 1623621585
transform 1 0 28520 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_310
timestamp 1623621585
transform 1 0 29624 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_322
timestamp 1623621585
transform 1 0 30728 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1623621585
transform 1 0 32568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_334
timestamp 1623621585
transform 1 0 31832 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_343
timestamp 1623621585
transform 1 0 32660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_355
timestamp 1623621585
transform 1 0 33764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_367
timestamp 1623621585
transform 1 0 34868 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_375
timestamp 1623621585
transform 1 0 35604 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0734_
timestamp 1623621585
transform 1 0 35880 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input173
timestamp 1623621585
transform 1 0 37168 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_386
timestamp 1623621585
transform 1 0 36616 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_395
timestamp 1623621585
transform 1 0 37444 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1623621585
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1623621585
transform 1 0 37812 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_400
timestamp 1623621585
transform 1 0 37904 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1623621585
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1623621585
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input388
timestamp 1623621585
transform 1 0 1380 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_6
timestamp 1623621585
transform 1 0 1656 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_18
timestamp 1623621585
transform 1 0 2760 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1623621585
transform 1 0 3772 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_26
timestamp 1623621585
transform 1 0 3496 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_30
timestamp 1623621585
transform 1 0 3864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_42
timestamp 1623621585
transform 1 0 4968 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_54
timestamp 1623621585
transform 1 0 6072 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_66
timestamp 1623621585
transform 1 0 7176 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_78
timestamp 1623621585
transform 1 0 8280 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1623621585
transform 1 0 9016 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_87
timestamp 1623621585
transform 1 0 9108 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_99
timestamp 1623621585
transform 1 0 10212 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_111
timestamp 1623621585
transform 1 0 11316 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1623621585
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1623621585
transform 1 0 14260 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1623621585
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_144
timestamp 1623621585
transform 1 0 14352 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_156
timestamp 1623621585
transform 1 0 15456 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_168
timestamp 1623621585
transform 1 0 16560 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_180
timestamp 1623621585
transform 1 0 17664 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0500_
timestamp 1623621585
transform 1 0 18400 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1623621585
transform 1 0 19504 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_196
timestamp 1623621585
transform 1 0 19136 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_201
timestamp 1623621585
transform 1 0 19596 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_213
timestamp 1623621585
transform 1 0 20700 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1623621585
transform 1 0 21804 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0755_
timestamp 1623621585
transform 1 0 23552 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0824_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22356 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1623621585
transform 1 0 23184 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1623621585
transform 1 0 24748 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 25208 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_49_252
timestamp 1623621585
transform 1 0 24288 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_256
timestamp 1623621585
transform 1 0 24656 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_258
timestamp 1623621585
transform 1 0 24840 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0631_
timestamp 1623621585
transform 1 0 27416 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_282
timestamp 1623621585
transform 1 0 27048 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_294
timestamp 1623621585
transform 1 0 28152 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_306
timestamp 1623621585
transform 1 0 29256 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1623621585
transform 1 0 29992 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_315
timestamp 1623621585
transform 1 0 30084 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_327
timestamp 1623621585
transform 1 0 31188 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_339
timestamp 1623621585
transform 1 0 32292 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_351
timestamp 1623621585
transform 1 0 33396 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1623621585
transform 1 0 35236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_363
timestamp 1623621585
transform 1 0 34500 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_372
timestamp 1623621585
transform 1 0 35328 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0726_
timestamp 1623621585
transform 1 0 35880 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1623621585
transform 1 0 37260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_386
timestamp 1623621585
transform 1 0 36616 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_392
timestamp 1623621585
transform 1 0 37168 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1623621585
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1623621585
transform 1 0 37904 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_396
timestamp 1623621585
transform 1 0 37536 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1623621585
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1623621585
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1623621585
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1623621585
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_27
timestamp 1623621585
transform 1 0 3588 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_39
timestamp 1623621585
transform 1 0 4692 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1623621585
transform 1 0 6348 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_51
timestamp 1623621585
transform 1 0 5796 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_58
timestamp 1623621585
transform 1 0 6440 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_70
timestamp 1623621585
transform 1 0 7544 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_82
timestamp 1623621585
transform 1 0 8648 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_94
timestamp 1623621585
transform 1 0 9752 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1623621585
transform 1 0 11592 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_106
timestamp 1623621585
transform 1 0 10856 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_115
timestamp 1623621585
transform 1 0 11684 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_127
timestamp 1623621585
transform 1 0 12788 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_139
timestamp 1623621585
transform 1 0 13892 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_151
timestamp 1623621585
transform 1 0 14996 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_163
timestamp 1623621585
transform 1 0 16100 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1623621585
transform 1 0 16836 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_172
timestamp 1623621585
transform 1 0 16928 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_184
timestamp 1623621585
transform 1 0 18032 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0472_
timestamp 1623621585
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_200
timestamp 1623621585
transform 1 0 19504 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1623621585
transform 1 0 22080 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_212
timestamp 1623621585
transform 1 0 20608 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1623621585
transform 1 0 21712 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1623621585
transform 1 0 22172 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0771_
timestamp 1623621585
transform 1 0 22540 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1623621585
transform 1 0 23276 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1623621585
transform 1 0 24012 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1623621585
transform 1 0 24288 0 -1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_50_269
timestamp 1623621585
transform 1 0 25852 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0606_
timestamp 1623621585
transform 1 0 26220 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1623621585
transform 1 0 27324 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_281
timestamp 1623621585
transform 1 0 26956 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_286
timestamp 1623621585
transform 1 0 27416 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_298
timestamp 1623621585
transform 1 0 28520 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_310
timestamp 1623621585
transform 1 0 29624 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_322
timestamp 1623621585
transform 1 0 30728 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1623621585
transform 1 0 32568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_334
timestamp 1623621585
transform 1 0 31832 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_343
timestamp 1623621585
transform 1 0 32660 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input174
timestamp 1623621585
transform 1 0 35328 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_355
timestamp 1623621585
transform 1 0 33764 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_367
timestamp 1623621585
transform 1 0 34868 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_371
timestamp 1623621585
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_375
timestamp 1623621585
transform 1 0 35604 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0718_
timestamp 1623621585
transform 1 0 35972 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1623621585
transform 1 0 37168 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_387
timestamp 1623621585
transform 1 0 36708 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_391
timestamp 1623621585
transform 1 0 37076 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_395
timestamp 1623621585
transform 1 0 37444 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1623621585
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1623621585
transform 1 0 37812 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_400
timestamp 1623621585
transform 1 0 37904 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1623621585
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1623621585
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input389
timestamp 1623621585
transform 1 0 1380 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_6
timestamp 1623621585
transform 1 0 1656 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_18
timestamp 1623621585
transform 1 0 2760 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1623621585
transform 1 0 3772 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_26
timestamp 1623621585
transform 1 0 3496 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1623621585
transform 1 0 3864 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1623621585
transform 1 0 4968 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_54
timestamp 1623621585
transform 1 0 6072 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_66
timestamp 1623621585
transform 1 0 7176 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_78
timestamp 1623621585
transform 1 0 8280 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1623621585
transform 1 0 9016 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_87
timestamp 1623621585
transform 1 0 9108 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_99
timestamp 1623621585
transform 1 0 10212 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_111
timestamp 1623621585
transform 1 0 11316 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1623621585
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1623621585
transform 1 0 14260 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1623621585
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_144
timestamp 1623621585
transform 1 0 14352 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_156
timestamp 1623621585
transform 1 0 15456 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_168
timestamp 1623621585
transform 1 0 16560 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_180
timestamp 1623621585
transform 1 0 17664 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1623621585
transform 1 0 19504 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_192
timestamp 1623621585
transform 1 0 18768 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_201
timestamp 1623621585
transform 1 0 19596 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_213
timestamp 1623621585
transform 1 0 20700 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1623621585
transform 1 0 21804 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1623621585
transform 1 0 22908 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_249
timestamp 1623621585
transform 1 0 24012 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1623621585
transform 1 0 25208 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1623621585
transform 1 0 24748 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_258
timestamp 1623621585
transform 1 0 24840 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1623621585
transform 1 0 27140 0 1 29920
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_51_279
timestamp 1623621585
transform 1 0 26772 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_300
timestamp 1623621585
transform 1 0 28704 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_312
timestamp 1623621585
transform 1 0 29808 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1623621585
transform 1 0 29992 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_315
timestamp 1623621585
transform 1 0 30084 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_327
timestamp 1623621585
transform 1 0 31188 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_339
timestamp 1623621585
transform 1 0 32292 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_351
timestamp 1623621585
transform 1 0 33396 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1623621585
transform 1 0 35236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_363
timestamp 1623621585
transform 1 0 34500 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_372
timestamp 1623621585
transform 1 0 35328 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0704_
timestamp 1623621585
transform 1 0 35972 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_378
timestamp 1623621585
transform 1 0 35880 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_387
timestamp 1623621585
transform 1 0 36708 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_395
timestamp 1623621585
transform 1 0 37444 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 37536 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1623621585
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1623621585
transform 1 0 38180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1623621585
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1623621585
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input390
timestamp 1623621585
transform 1 0 1380 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1623621585
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1623621585
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_6
timestamp 1623621585
transform 1 0 1656 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_18
timestamp 1623621585
transform 1 0 2760 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1623621585
transform 1 0 3772 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_27
timestamp 1623621585
transform 1 0 3588 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_39
timestamp 1623621585
transform 1 0 4692 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_26
timestamp 1623621585
transform 1 0 3496 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1623621585
transform 1 0 3864 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1623621585
transform 1 0 6348 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_51
timestamp 1623621585
transform 1 0 5796 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_58
timestamp 1623621585
transform 1 0 6440 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1623621585
transform 1 0 4968 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_54
timestamp 1623621585
transform 1 0 6072 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_70
timestamp 1623621585
transform 1 0 7544 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_82
timestamp 1623621585
transform 1 0 8648 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_66
timestamp 1623621585
transform 1 0 7176 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_78
timestamp 1623621585
transform 1 0 8280 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1623621585
transform 1 0 9016 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_94
timestamp 1623621585
transform 1 0 9752 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_87
timestamp 1623621585
transform 1 0 9108 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_99
timestamp 1623621585
transform 1 0 10212 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1623621585
transform 1 0 11592 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_106
timestamp 1623621585
transform 1 0 10856 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_115
timestamp 1623621585
transform 1 0 11684 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_111
timestamp 1623621585
transform 1 0 11316 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1623621585
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1623621585
transform 1 0 14260 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_127
timestamp 1623621585
transform 1 0 12788 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_139
timestamp 1623621585
transform 1 0 13892 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1623621585
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_144
timestamp 1623621585
transform 1 0 14352 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_151
timestamp 1623621585
transform 1 0 14996 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_163
timestamp 1623621585
transform 1 0 16100 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_156
timestamp 1623621585
transform 1 0 15456 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1623621585
transform 1 0 16836 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_172
timestamp 1623621585
transform 1 0 16928 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_184
timestamp 1623621585
transform 1 0 18032 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_168
timestamp 1623621585
transform 1 0 16560 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_180
timestamp 1623621585
transform 1 0 17664 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1623621585
transform 1 0 19504 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_196
timestamp 1623621585
transform 1 0 19136 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_208
timestamp 1623621585
transform 1 0 20240 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_192
timestamp 1623621585
transform 1 0 18768 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_201
timestamp 1623621585
transform 1 0 19596 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1623621585
transform 1 0 22080 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_220
timestamp 1623621585
transform 1 0 21344 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_229
timestamp 1623621585
transform 1 0 22172 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_213
timestamp 1623621585
transform 1 0 20700 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1623621585
transform 1 0 21804 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_241
timestamp 1623621585
transform 1 0 23276 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1623621585
transform 1 0 22908 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_249
timestamp 1623621585
transform 1 0 24012 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0496_
timestamp 1623621585
transform 1 0 25208 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0614_
timestamp 1623621585
transform 1 0 25944 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1002_
timestamp 1623621585
transform 1 0 25300 0 -1 31008
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1623621585
transform 1 0 24748 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_253
timestamp 1623621585
transform 1 0 24380 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_261
timestamp 1623621585
transform 1 0 25116 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1623621585
transform 1 0 24840 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_266
timestamp 1623621585
transform 1 0 25576 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0605_
timestamp 1623621585
transform 1 0 27784 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0768_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 27048 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1623621585
transform 1 0 27324 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_280
timestamp 1623621585
transform 1 0 26864 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_284
timestamp 1623621585
transform 1 0 27232 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_286
timestamp 1623621585
transform 1 0 27416 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_278
timestamp 1623621585
transform 1 0 26680 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_290
timestamp 1623621585
transform 1 0 27784 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0551_
timestamp 1623621585
transform 1 0 28152 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_293
timestamp 1623621585
transform 1 0 28060 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_305
timestamp 1623621585
transform 1 0 29164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_297
timestamp 1623621585
transform 1 0 28428 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_309
timestamp 1623621585
transform 1 0 29532 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1623621585
transform 1 0 29992 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_317
timestamp 1623621585
transform 1 0 30268 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_329
timestamp 1623621585
transform 1 0 31372 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_313
timestamp 1623621585
transform 1 0 29900 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_315
timestamp 1623621585
transform 1 0 30084 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_327
timestamp 1623621585
transform 1 0 31188 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1623621585
transform 1 0 32568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_341
timestamp 1623621585
transform 1 0 32476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_343
timestamp 1623621585
transform 1 0 32660 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_339
timestamp 1623621585
transform 1 0 32292 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_351
timestamp 1623621585
transform 1 0 33396 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1623621585
transform 1 0 35236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_355
timestamp 1623621585
transform 1 0 33764 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_367
timestamp 1623621585
transform 1 0 34868 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_375
timestamp 1623621585
transform 1 0 35604 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_363
timestamp 1623621585
transform 1 0 34500 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_372
timestamp 1623621585
transform 1 0 35328 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0701_
timestamp 1623621585
transform 1 0 37168 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0733_
timestamp 1623621585
transform 1 0 36524 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1623621585
transform 1 0 36524 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input175
timestamp 1623621585
transform 1 0 35880 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_381
timestamp 1623621585
transform 1 0 36156 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_388
timestamp 1623621585
transform 1 0 36800 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_395
timestamp 1623621585
transform 1 0 37444 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_384
timestamp 1623621585
transform 1 0 36432 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_392
timestamp 1623621585
transform 1 0 37168 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp 1623621585
transform 1 0 37536 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1623621585
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1623621585
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1623621585
transform 1 0 37812 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_400
timestamp 1623621585
transform 1 0 37904 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1623621585
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1623621585
transform 1 0 38180 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1623621585
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input391
timestamp 1623621585
transform 1 0 1380 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1623621585
transform 1 0 1656 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_18
timestamp 1623621585
transform 1 0 2760 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1623621585
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1623621585
transform 1 0 6348 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1623621585
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_54
timestamp 1623621585
transform 1 0 6072 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_58
timestamp 1623621585
transform 1 0 6440 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_70
timestamp 1623621585
transform 1 0 7544 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_82
timestamp 1623621585
transform 1 0 8648 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_94
timestamp 1623621585
transform 1 0 9752 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1623621585
transform 1 0 11592 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_106
timestamp 1623621585
transform 1 0 10856 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_115
timestamp 1623621585
transform 1 0 11684 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_127
timestamp 1623621585
transform 1 0 12788 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_139
timestamp 1623621585
transform 1 0 13892 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_151
timestamp 1623621585
transform 1 0 14996 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_163
timestamp 1623621585
transform 1 0 16100 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1623621585
transform 1 0 16836 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_172
timestamp 1623621585
transform 1 0 16928 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_184
timestamp 1623621585
transform 1 0 18032 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_196
timestamp 1623621585
transform 1 0 19136 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_208
timestamp 1623621585
transform 1 0 20240 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1623621585
transform 1 0 22080 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_220
timestamp 1623621585
transform 1 0 21344 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_229
timestamp 1623621585
transform 1 0 22172 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0402_
timestamp 1623621585
transform 1 0 22540 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_236
timestamp 1623621585
transform 1 0 22816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_248
timestamp 1623621585
transform 1 0 23920 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0727_
timestamp 1623621585
transform 1 0 25944 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0744_
timestamp 1623621585
transform 1 0 24840 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_256
timestamp 1623621585
transform 1 0 24656 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_266
timestamp 1623621585
transform 1 0 25576 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0760_
timestamp 1623621585
transform 1 0 27784 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1623621585
transform 1 0 27324 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_278
timestamp 1623621585
transform 1 0 26680 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_284
timestamp 1623621585
transform 1 0 27232 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_286
timestamp 1623621585
transform 1 0 27416 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_298
timestamp 1623621585
transform 1 0 28520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_310
timestamp 1623621585
transform 1 0 29624 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_322
timestamp 1623621585
transform 1 0 30728 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1623621585
transform 1 0 32568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_334
timestamp 1623621585
transform 1 0 31832 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_343
timestamp 1623621585
transform 1 0 32660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input176
timestamp 1623621585
transform 1 0 35512 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_355
timestamp 1623621585
transform 1 0 33764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_367
timestamp 1623621585
transform 1 0 34868 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 1623621585
transform 1 0 35420 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1623621585
transform 1 0 36800 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1623621585
transform 1 0 36156 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_377
timestamp 1623621585
transform 1 0 35788 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_384
timestamp 1623621585
transform 1 0 36432 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_395
timestamp 1623621585
transform 1 0 37444 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1623621585
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1623621585
transform 1 0 37812 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_400
timestamp 1623621585
transform 1 0 37904 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1623621585
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1623621585
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1623621585
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1623621585
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1623621585
transform 1 0 3772 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_27
timestamp 1623621585
transform 1 0 3588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1623621585
transform 1 0 3864 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1623621585
transform 1 0 4968 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_54
timestamp 1623621585
transform 1 0 6072 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_66
timestamp 1623621585
transform 1 0 7176 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_78
timestamp 1623621585
transform 1 0 8280 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1623621585
transform 1 0 9016 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_87
timestamp 1623621585
transform 1 0 9108 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_99
timestamp 1623621585
transform 1 0 10212 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_111
timestamp 1623621585
transform 1 0 11316 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1623621585
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1623621585
transform 1 0 14260 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_135
timestamp 1623621585
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_144
timestamp 1623621585
transform 1 0 14352 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_156
timestamp 1623621585
transform 1 0 15456 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_168
timestamp 1623621585
transform 1 0 16560 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_180
timestamp 1623621585
transform 1 0 17664 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1623621585
transform 1 0 19504 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_192
timestamp 1623621585
transform 1 0 18768 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_201
timestamp 1623621585
transform 1 0 19596 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_213
timestamp 1623621585
transform 1 0 20700 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1623621585
transform 1 0 21804 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0403_
timestamp 1623621585
transform 1 0 23552 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_237
timestamp 1623621585
transform 1 0 22908 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_243
timestamp 1623621585
transform 1 0 23460 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_248
timestamp 1623621585
transform 1 0 23920 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0736_
timestamp 1623621585
transform 1 0 25392 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1623621585
transform 1 0 24748 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_256
timestamp 1623621585
transform 1 0 24656 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_258
timestamp 1623621585
transform 1 0 24840 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _0585_
timestamp 1623621585
transform 1 0 26496 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0752_
timestamp 1623621585
transform 1 0 27600 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_272
timestamp 1623621585
transform 1 0 26128 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_284
timestamp 1623621585
transform 1 0 27232 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_296
timestamp 1623621585
transform 1 0 28336 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_308
timestamp 1623621585
transform 1 0 29440 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1623621585
transform 1 0 29992 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_315
timestamp 1623621585
transform 1 0 30084 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_327
timestamp 1623621585
transform 1 0 31188 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_339
timestamp 1623621585
transform 1 0 32292 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_351
timestamp 1623621585
transform 1 0 33396 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1623621585
transform 1 0 35236 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_363
timestamp 1623621585
transform 1 0 34500 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_372
timestamp 1623621585
transform 1 0 35328 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0645_
timestamp 1623621585
transform 1 0 36064 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1623621585
transform 1 0 36892 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_383
timestamp 1623621585
transform 1 0 36340 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_392
timestamp 1623621585
transform 1 0 37168 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0703_
timestamp 1623621585
transform 1 0 37536 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1623621585
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1623621585
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1623621585
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input392
timestamp 1623621585
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1623621585
transform 1 0 1656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_18
timestamp 1623621585
transform 1 0 2760 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1623621585
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1623621585
transform 1 0 6348 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1623621585
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_54
timestamp 1623621585
transform 1 0 6072 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_58
timestamp 1623621585
transform 1 0 6440 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_70
timestamp 1623621585
transform 1 0 7544 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_82
timestamp 1623621585
transform 1 0 8648 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_94
timestamp 1623621585
transform 1 0 9752 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1623621585
transform 1 0 11592 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_106
timestamp 1623621585
transform 1 0 10856 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_115
timestamp 1623621585
transform 1 0 11684 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_127
timestamp 1623621585
transform 1 0 12788 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_139
timestamp 1623621585
transform 1 0 13892 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_151
timestamp 1623621585
transform 1 0 14996 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_163
timestamp 1623621585
transform 1 0 16100 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1623621585
transform 1 0 16836 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_172
timestamp 1623621585
transform 1 0 16928 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_184
timestamp 1623621585
transform 1 0 18032 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_196
timestamp 1623621585
transform 1 0 19136 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_208
timestamp 1623621585
transform 1 0 20240 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1623621585
transform 1 0 22080 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_220
timestamp 1623621585
transform 1 0 21344 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_229
timestamp 1623621585
transform 1 0 22172 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_241
timestamp 1623621585
transform 1 0 23276 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0719_
timestamp 1623621585
transform 1 0 25116 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 1623621585
transform 1 0 24380 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_269
timestamp 1623621585
transform 1 0 25852 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0577_
timestamp 1623621585
transform 1 0 26220 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1008_
timestamp 1623621585
transform 1 0 27784 0 -1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1623621585
transform 1 0 27324 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_281
timestamp 1623621585
transform 1 0 26956 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_286
timestamp 1623621585
transform 1 0 27416 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_307
timestamp 1623621585
transform 1 0 29348 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_319
timestamp 1623621585
transform 1 0 30452 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_331
timestamp 1623621585
transform 1 0 31556 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1623621585
transform 1 0 32568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_339
timestamp 1623621585
transform 1 0 32292 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_343
timestamp 1623621585
transform 1 0 32660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input177
timestamp 1623621585
transform 1 0 35420 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_355
timestamp 1623621585
transform 1 0 33764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_367
timestamp 1623621585
transform 1 0 34868 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0689_
timestamp 1623621585
transform 1 0 36064 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1623621585
transform 1 0 37168 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_376
timestamp 1623621585
transform 1 0 35696 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_388
timestamp 1623621585
transform 1 0 36800 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1623621585
transform 1 0 37444 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1623621585
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1623621585
transform 1 0 37812 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_400
timestamp 1623621585
transform 1 0 37904 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1623621585
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1623621585
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input393
timestamp 1623621585
transform 1 0 1748 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1623621585
transform 1 0 1380 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_11
timestamp 1623621585
transform 1 0 2116 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1623621585
transform 1 0 3772 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_23
timestamp 1623621585
transform 1 0 3220 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1623621585
transform 1 0 3864 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1623621585
transform 1 0 4968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_54
timestamp 1623621585
transform 1 0 6072 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_66
timestamp 1623621585
transform 1 0 7176 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_78
timestamp 1623621585
transform 1 0 8280 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1623621585
transform 1 0 9016 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_87
timestamp 1623621585
transform 1 0 9108 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_99
timestamp 1623621585
transform 1 0 10212 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_111
timestamp 1623621585
transform 1 0 11316 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1623621585
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1623621585
transform 1 0 14260 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1623621585
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_144
timestamp 1623621585
transform 1 0 14352 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_156
timestamp 1623621585
transform 1 0 15456 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_168
timestamp 1623621585
transform 1 0 16560 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_180
timestamp 1623621585
transform 1 0 17664 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1623621585
transform 1 0 19504 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_192
timestamp 1623621585
transform 1 0 18768 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_201
timestamp 1623621585
transform 1 0 19596 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_213
timestamp 1623621585
transform 1 0 20700 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1623621585
transform 1 0 21804 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1623621585
transform 1 0 22908 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_249
timestamp 1623621585
transform 1 0 24012 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0710_
timestamp 1623621585
transform 1 0 25208 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1623621585
transform 1 0 24748 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_258
timestamp 1623621585
transform 1 0 24840 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_270
timestamp 1623621585
transform 1 0 25944 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1004_
timestamp 1623621585
transform 1 0 26312 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_57_291
timestamp 1623621585
transform 1 0 27876 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0568_
timestamp 1623621585
transform 1 0 28244 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_303
timestamp 1623621585
transform 1 0 28980 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_311
timestamp 1623621585
transform 1 0 29716 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1623621585
transform 1 0 29992 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_315
timestamp 1623621585
transform 1 0 30084 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_327
timestamp 1623621585
transform 1 0 31188 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_339
timestamp 1623621585
transform 1 0 32292 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_351
timestamp 1623621585
transform 1 0 33396 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1623621585
transform 1 0 35236 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_363
timestamp 1623621585
transform 1 0 34500 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_372
timestamp 1623621585
transform 1 0 35328 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0680_
timestamp 1623621585
transform 1 0 36064 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1623621585
transform 1 0 37260 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1623621585
transform 1 0 36800 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_392
timestamp 1623621585
transform 1 0 37168 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1623621585
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1623621585
transform 1 0 37904 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_396
timestamp 1623621585
transform 1 0 37536 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1623621585
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1623621585
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1623621585
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1623621585
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_27
timestamp 1623621585
transform 1 0 3588 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_39
timestamp 1623621585
transform 1 0 4692 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1623621585
transform 1 0 6348 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_51
timestamp 1623621585
transform 1 0 5796 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_58
timestamp 1623621585
transform 1 0 6440 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_70
timestamp 1623621585
transform 1 0 7544 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_82
timestamp 1623621585
transform 1 0 8648 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_94
timestamp 1623621585
transform 1 0 9752 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1623621585
transform 1 0 11592 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_106
timestamp 1623621585
transform 1 0 10856 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_115
timestamp 1623621585
transform 1 0 11684 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_127
timestamp 1623621585
transform 1 0 12788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_139
timestamp 1623621585
transform 1 0 13892 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_151
timestamp 1623621585
transform 1 0 14996 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_163
timestamp 1623621585
transform 1 0 16100 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1623621585
transform 1 0 16836 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_172
timestamp 1623621585
transform 1 0 16928 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_184
timestamp 1623621585
transform 1 0 18032 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_196
timestamp 1623621585
transform 1 0 19136 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_208
timestamp 1623621585
transform 1 0 20240 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1623621585
transform 1 0 22080 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_220
timestamp 1623621585
transform 1 0 21344 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_229
timestamp 1623621585
transform 1 0 22172 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_241
timestamp 1623621585
transform 1 0 23276 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0438_
timestamp 1623621585
transform 1 0 25392 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_253
timestamp 1623621585
transform 1 0 24380 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_261
timestamp 1623621585
transform 1 0 25116 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_268
timestamp 1623621585
transform 1 0 25760 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0560_
timestamp 1623621585
transform 1 0 26220 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1006_
timestamp 1623621585
transform 1 0 27784 0 -1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1623621585
transform 1 0 27324 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_272
timestamp 1623621585
transform 1 0 26128 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_281
timestamp 1623621585
transform 1 0 26956 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1623621585
transform 1 0 27416 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0497_
timestamp 1623621585
transform 1 0 29716 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_307
timestamp 1623621585
transform 1 0 29348 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1623621585
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1623621585
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1623621585
transform 1 0 32568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_339
timestamp 1623621585
transform 1 0 32292 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_343
timestamp 1623621585
transform 1 0 32660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1623621585
transform 1 0 35420 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_355
timestamp 1623621585
transform 1 0 33764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_367
timestamp 1623621585
transform 1 0 34868 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0672_
timestamp 1623621585
transform 1 0 36064 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1623621585
transform 1 0 37168 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_376
timestamp 1623621585
transform 1 0 35696 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_388
timestamp 1623621585
transform 1 0 36800 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_395
timestamp 1623621585
transform 1 0 37444 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1623621585
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1623621585
transform 1 0 37812 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_400
timestamp 1623621585
transform 1 0 37904 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1623621585
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1623621585
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1623621585
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input364
timestamp 1623621585
transform 1 0 1380 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input394
timestamp 1623621585
transform 1 0 1380 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1623621585
transform 1 0 1656 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_18
timestamp 1623621585
transform 1 0 2760 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_6
timestamp 1623621585
transform 1 0 1656 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_18
timestamp 1623621585
transform 1 0 2760 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1623621585
transform 1 0 3772 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_26
timestamp 1623621585
transform 1 0 3496 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1623621585
transform 1 0 3864 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1623621585
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1623621585
transform 1 0 6348 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1623621585
transform 1 0 4968 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_54
timestamp 1623621585
transform 1 0 6072 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1623621585
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_54
timestamp 1623621585
transform 1 0 6072 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_58
timestamp 1623621585
transform 1 0 6440 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_66
timestamp 1623621585
transform 1 0 7176 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_78
timestamp 1623621585
transform 1 0 8280 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_70
timestamp 1623621585
transform 1 0 7544 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_82
timestamp 1623621585
transform 1 0 8648 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1623621585
transform 1 0 9016 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_87
timestamp 1623621585
transform 1 0 9108 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_99
timestamp 1623621585
transform 1 0 10212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_94
timestamp 1623621585
transform 1 0 9752 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1623621585
transform 1 0 11592 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_111
timestamp 1623621585
transform 1 0 11316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1623621585
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_106
timestamp 1623621585
transform 1 0 10856 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_115
timestamp 1623621585
transform 1 0 11684 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1623621585
transform 1 0 14260 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1623621585
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_144
timestamp 1623621585
transform 1 0 14352 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_127
timestamp 1623621585
transform 1 0 12788 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_139
timestamp 1623621585
transform 1 0 13892 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_156
timestamp 1623621585
transform 1 0 15456 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_151
timestamp 1623621585
transform 1 0 14996 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_163
timestamp 1623621585
transform 1 0 16100 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1623621585
transform 1 0 16836 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_168
timestamp 1623621585
transform 1 0 16560 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_180
timestamp 1623621585
transform 1 0 17664 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_172
timestamp 1623621585
transform 1 0 16928 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_184
timestamp 1623621585
transform 1 0 18032 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1623621585
transform 1 0 19504 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_192
timestamp 1623621585
transform 1 0 18768 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_201
timestamp 1623621585
transform 1 0 19596 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_196
timestamp 1623621585
transform 1 0 19136 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_208
timestamp 1623621585
transform 1 0 20240 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1623621585
transform 1 0 22080 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_213
timestamp 1623621585
transform 1 0 20700 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1623621585
transform 1 0 21804 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_220
timestamp 1623621585
transform 1 0 21344 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_229
timestamp 1623621585
transform 1 0 22172 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0405_
timestamp 1623621585
transform 1 0 23368 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1623621585
transform 1 0 22908 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1623621585
transform 1 0 24012 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_241
timestamp 1623621585
transform 1 0 23276 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_245
timestamp 1623621585
transform 1 0 23644 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1623621585
transform 1 0 24748 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1623621585
transform 1 0 25208 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_258
timestamp 1623621585
transform 1 0 24840 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_265
timestamp 1623621585
transform 1 0 25484 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_257
timestamp 1623621585
transform 1 0 24748 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_269
timestamp 1623621585
transform 1 0 25852 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1005_
timestamp 1623621585
transform 1 0 26680 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1007_
timestamp 1623621585
transform 1 0 27784 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1623621585
transform 1 0 27324 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1623621585
transform 1 0 26036 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_274
timestamp 1623621585
transform 1 0 26312 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_281
timestamp 1623621585
transform 1 0 26956 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1623621585
transform 1 0 27416 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0552_
timestamp 1623621585
transform 1 0 28612 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_295
timestamp 1623621585
transform 1 0 28244 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_307
timestamp 1623621585
transform 1 0 29348 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_307
timestamp 1623621585
transform 1 0 29348 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1623621585
transform 1 0 29992 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_313
timestamp 1623621585
transform 1 0 29900 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_315
timestamp 1623621585
transform 1 0 30084 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_327
timestamp 1623621585
transform 1 0 31188 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_319
timestamp 1623621585
transform 1 0 30452 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_331
timestamp 1623621585
transform 1 0 31556 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1623621585
transform 1 0 32568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_339
timestamp 1623621585
transform 1 0 32292 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_351
timestamp 1623621585
transform 1 0 33396 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_339
timestamp 1623621585
transform 1 0 32292 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_343
timestamp 1623621585
transform 1 0 32660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0473_
timestamp 1623621585
transform 1 0 35328 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1623621585
transform 1 0 35236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input178
timestamp 1623621585
transform 1 0 34592 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_363
timestamp 1623621585
transform 1 0 34500 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1623621585
transform 1 0 34868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_372
timestamp 1623621585
transform 1 0 35328 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_355
timestamp 1623621585
transform 1 0 33764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_367
timestamp 1623621585
transform 1 0 34868 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_371
timestamp 1623621585
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0647_
timestamp 1623621585
transform 1 0 37168 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0650_
timestamp 1623621585
transform 1 0 36064 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0664_
timestamp 1623621585
transform 1 0 36064 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_388
timestamp 1623621585
transform 1 0 36800 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_376
timestamp 1623621585
transform 1 0 35696 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_388
timestamp 1623621585
transform 1 0 36800 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_395
timestamp 1623621585
transform 1 0 37444 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0688_
timestamp 1623621585
transform 1 0 37536 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1623621585
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1623621585
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1623621585
transform 1 0 37812 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1623621585
transform 1 0 38180 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_400
timestamp 1623621585
transform 1 0 37904 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1623621585
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1623621585
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1623621585
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1623621585
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1623621585
transform 1 0 3772 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_27
timestamp 1623621585
transform 1 0 3588 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1623621585
transform 1 0 3864 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1623621585
transform 1 0 4968 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_54
timestamp 1623621585
transform 1 0 6072 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_66
timestamp 1623621585
transform 1 0 7176 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_78
timestamp 1623621585
transform 1 0 8280 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1623621585
transform 1 0 9016 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_87
timestamp 1623621585
transform 1 0 9108 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_99
timestamp 1623621585
transform 1 0 10212 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_111
timestamp 1623621585
transform 1 0 11316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1623621585
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1623621585
transform 1 0 14260 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1623621585
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_144
timestamp 1623621585
transform 1 0 14352 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_156
timestamp 1623621585
transform 1 0 15456 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_168
timestamp 1623621585
transform 1 0 16560 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_180
timestamp 1623621585
transform 1 0 17664 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1623621585
transform 1 0 19504 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_192
timestamp 1623621585
transform 1 0 18768 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_201
timestamp 1623621585
transform 1 0 19596 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_213
timestamp 1623621585
transform 1 0 20700 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1623621585
transform 1 0 21804 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0404_
timestamp 1623621585
transform 1 0 23920 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0408_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22632 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_233
timestamp 1623621585
transform 1 0 22540 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_238
timestamp 1623621585
transform 1 0 23000 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_246
timestamp 1623621585
transform 1 0 23736 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1623621585
transform 1 0 24748 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_251
timestamp 1623621585
transform 1 0 24196 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_258
timestamp 1623621585
transform 1 0 24840 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_270
timestamp 1623621585
transform 1 0 25944 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_282
timestamp 1623621585
transform 1 0 27048 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_294
timestamp 1623621585
transform 1 0 28152 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_306
timestamp 1623621585
transform 1 0 29256 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1623621585
transform 1 0 29992 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_315
timestamp 1623621585
transform 1 0 30084 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_327
timestamp 1623621585
transform 1 0 31188 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_339
timestamp 1623621585
transform 1 0 32292 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_351
timestamp 1623621585
transform 1 0 33396 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1623621585
transform 1 0 35236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1623621585
transform 1 0 34592 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_363
timestamp 1623621585
transform 1 0 34500 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_367
timestamp 1623621585
transform 1 0 34868 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_372
timestamp 1623621585
transform 1 0 35328 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0751_
timestamp 1623621585
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0759_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 35880 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_61_387
timestamp 1623621585
transform 1 0 36708 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1623621585
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_399
timestamp 1623621585
transform 1 0 37812 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1623621585
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input365
timestamp 1623621585
transform 1 0 1380 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_6
timestamp 1623621585
transform 1 0 1656 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_18
timestamp 1623621585
transform 1 0 2760 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1623621585
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1623621585
transform 1 0 6348 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1623621585
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_54
timestamp 1623621585
transform 1 0 6072 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_58
timestamp 1623621585
transform 1 0 6440 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_70
timestamp 1623621585
transform 1 0 7544 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_82
timestamp 1623621585
transform 1 0 8648 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_94
timestamp 1623621585
transform 1 0 9752 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1623621585
transform 1 0 11592 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_106
timestamp 1623621585
transform 1 0 10856 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_115
timestamp 1623621585
transform 1 0 11684 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_127
timestamp 1623621585
transform 1 0 12788 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_139
timestamp 1623621585
transform 1 0 13892 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_151
timestamp 1623621585
transform 1 0 14996 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_163
timestamp 1623621585
transform 1 0 16100 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1623621585
transform 1 0 16836 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_172
timestamp 1623621585
transform 1 0 16928 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_184
timestamp 1623621585
transform 1 0 18032 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_196
timestamp 1623621585
transform 1 0 19136 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_208
timestamp 1623621585
transform 1 0 20240 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0406_
timestamp 1623621585
transform 1 0 21436 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1623621585
transform 1 0 22080 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_220
timestamp 1623621585
transform 1 0 21344 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_224
timestamp 1623621585
transform 1 0 21712 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_229
timestamp 1623621585
transform 1 0 22172 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1623621585
transform 1 0 23092 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_62_237
timestamp 1623621585
transform 1 0 22908 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_255
timestamp 1623621585
transform 1 0 24564 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_267
timestamp 1623621585
transform 1 0 25668 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0690_
timestamp 1623621585
transform 1 0 26220 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1623621585
transform 1 0 27324 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_281
timestamp 1623621585
transform 1 0 26956 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_286
timestamp 1623621585
transform 1 0 27416 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_298
timestamp 1623621585
transform 1 0 28520 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_310
timestamp 1623621585
transform 1 0 29624 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_322
timestamp 1623621585
transform 1 0 30728 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1623621585
transform 1 0 32568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_334
timestamp 1623621585
transform 1 0 31832 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_343
timestamp 1623621585
transform 1 0 32660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1623621585
transform 1 0 35236 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input179
timestamp 1623621585
transform 1 0 34592 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1623621585
transform 1 0 33764 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1623621585
transform 1 0 34500 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_367
timestamp 1623621585
transform 1 0 34868 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_374
timestamp 1623621585
transform 1 0 35512 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0591_
timestamp 1623621585
transform 1 0 37076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_2  _0767_
timestamp 1623621585
transform 1 0 35880 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_62_387
timestamp 1623621585
transform 1 0 36708 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1623621585
transform 1 0 37444 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1623621585
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1623621585
transform 1 0 37812 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_400
timestamp 1623621585
transform 1 0 37904 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1623621585
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1623621585
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input366
timestamp 1623621585
transform 1 0 1380 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_6
timestamp 1623621585
transform 1 0 1656 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_18
timestamp 1623621585
transform 1 0 2760 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1623621585
transform 1 0 3772 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_26
timestamp 1623621585
transform 1 0 3496 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1623621585
transform 1 0 3864 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1623621585
transform 1 0 4968 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_54
timestamp 1623621585
transform 1 0 6072 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_66
timestamp 1623621585
transform 1 0 7176 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_78
timestamp 1623621585
transform 1 0 8280 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1623621585
transform 1 0 9016 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_87
timestamp 1623621585
transform 1 0 9108 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_99
timestamp 1623621585
transform 1 0 10212 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_111
timestamp 1623621585
transform 1 0 11316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1623621585
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1623621585
transform 1 0 14260 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1623621585
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_144
timestamp 1623621585
transform 1 0 14352 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_156
timestamp 1623621585
transform 1 0 15456 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_168
timestamp 1623621585
transform 1 0 16560 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_180
timestamp 1623621585
transform 1 0 17664 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1623621585
transform 1 0 19504 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_192
timestamp 1623621585
transform 1 0 18768 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_201
timestamp 1623621585
transform 1 0 19596 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1016_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 21252 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_63_213
timestamp 1623621585
transform 1 0 20700 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 23460 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1623621585
transform 1 0 23000 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_242
timestamp 1623621585
transform 1 0 23368 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_250
timestamp 1623621585
transform 1 0 24104 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1623621585
transform 1 0 24748 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_256
timestamp 1623621585
transform 1 0 24656 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_258
timestamp 1623621585
transform 1 0 24840 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_270
timestamp 1623621585
transform 1 0 25944 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0682_
timestamp 1623621585
transform 1 0 26220 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1623621585
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0523_
timestamp 1623621585
transform 1 0 28152 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_293
timestamp 1623621585
transform 1 0 28060 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_302
timestamp 1623621585
transform 1 0 28888 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1623621585
transform 1 0 29992 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_315
timestamp 1623621585
transform 1 0 30084 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_327
timestamp 1623621585
transform 1 0 31188 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_339
timestamp 1623621585
transform 1 0 32292 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_351
timestamp 1623621585
transform 1 0 33396 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1623621585
transform 1 0 35236 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_363
timestamp 1623621585
transform 1 0 34500 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_372
timestamp 1623621585
transform 1 0 35328 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0679_
timestamp 1623621585
transform 1 0 36524 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0700_
timestamp 1623621585
transform 1 0 35788 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_376
timestamp 1623621585
transform 1 0 35696 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_381
timestamp 1623621585
transform 1 0 36156 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_392
timestamp 1623621585
transform 1 0 37168 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0663_
timestamp 1623621585
transform 1 0 37536 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1623621585
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1623621585
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1623621585
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1623621585
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1623621585
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_27
timestamp 1623621585
transform 1 0 3588 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_39
timestamp 1623621585
transform 1 0 4692 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1623621585
transform 1 0 6348 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_51
timestamp 1623621585
transform 1 0 5796 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_58
timestamp 1623621585
transform 1 0 6440 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_70
timestamp 1623621585
transform 1 0 7544 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_82
timestamp 1623621585
transform 1 0 8648 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1623621585
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1623621585
transform 1 0 11592 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_106
timestamp 1623621585
transform 1 0 10856 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_115
timestamp 1623621585
transform 1 0 11684 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_127
timestamp 1623621585
transform 1 0 12788 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_139
timestamp 1623621585
transform 1 0 13892 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_151
timestamp 1623621585
transform 1 0 14996 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_163
timestamp 1623621585
transform 1 0 16100 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1623621585
transform 1 0 16836 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_172
timestamp 1623621585
transform 1 0 16928 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_184
timestamp 1623621585
transform 1 0 18032 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_196
timestamp 1623621585
transform 1 0 19136 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_208
timestamp 1623621585
transform 1 0 20240 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1623621585
transform 1 0 22080 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_220
timestamp 1623621585
transform 1 0 21344 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_229
timestamp 1623621585
transform 1 0 22172 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0407_
timestamp 1623621585
transform 1 0 22908 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 24104 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_64_246
timestamp 1623621585
transform 1 0 23736 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_255
timestamp 1623621585
transform 1 0 24564 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_267
timestamp 1623621585
transform 1 0 25668 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0673_
timestamp 1623621585
transform 1 0 26220 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1623621585
transform 1 0 27324 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_281
timestamp 1623621585
transform 1 0 26956 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_286
timestamp 1623621585
transform 1 0 27416 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0514_
timestamp 1623621585
transform 1 0 28336 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0531_
timestamp 1623621585
transform 1 0 29440 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_294
timestamp 1623621585
transform 1 0 28152 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1623621585
transform 1 0 29072 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_316
timestamp 1623621585
transform 1 0 30176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_328
timestamp 1623621585
transform 1 0 31280 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1623621585
transform 1 0 32568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_340
timestamp 1623621585
transform 1 0 32384 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_343
timestamp 1623621585
transform 1 0 32660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input180
timestamp 1623621585
transform 1 0 35512 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_355
timestamp 1623621585
transform 1 0 33764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_367
timestamp 1623621585
transform 1 0 34868 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_373
timestamp 1623621585
transform 1 0 35420 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0671_
timestamp 1623621585
transform 1 0 36800 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1623621585
transform 1 0 36156 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 1623621585
transform 1 0 35788 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_384
timestamp 1623621585
transform 1 0 36432 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1623621585
transform 1 0 37444 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1623621585
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1623621585
transform 1 0 37812 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_400
timestamp 1623621585
transform 1 0 37904 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_406
timestamp 1623621585
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1623621585
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input367
timestamp 1623621585
transform 1 0 1748 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1623621585
transform 1 0 1380 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_11
timestamp 1623621585
transform 1 0 2116 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1623621585
transform 1 0 3772 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_23
timestamp 1623621585
transform 1 0 3220 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_30
timestamp 1623621585
transform 1 0 3864 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_42
timestamp 1623621585
transform 1 0 4968 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_54
timestamp 1623621585
transform 1 0 6072 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_66
timestamp 1623621585
transform 1 0 7176 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_78
timestamp 1623621585
transform 1 0 8280 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1623621585
transform 1 0 9016 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_87
timestamp 1623621585
transform 1 0 9108 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_99
timestamp 1623621585
transform 1 0 10212 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_111
timestamp 1623621585
transform 1 0 11316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1623621585
transform 1 0 12420 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1623621585
transform 1 0 14260 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_135
timestamp 1623621585
transform 1 0 13524 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_144
timestamp 1623621585
transform 1 0 14352 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_156
timestamp 1623621585
transform 1 0 15456 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_168
timestamp 1623621585
transform 1 0 16560 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_180
timestamp 1623621585
transform 1 0 17664 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1623621585
transform 1 0 19504 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_192
timestamp 1623621585
transform 1 0 18768 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_201
timestamp 1623621585
transform 1 0 19596 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0441_
timestamp 1623621585
transform 1 0 21712 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_213
timestamp 1623621585
transform 1 0 20700 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_221
timestamp 1623621585
transform 1 0 21436 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0413_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 24104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0449_
timestamp 1623621585
transform 1 0 22816 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_232
timestamp 1623621585
transform 1 0 22448 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_244
timestamp 1623621585
transform 1 0 23552 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1623621585
transform 1 0 24748 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_253
timestamp 1623621585
transform 1 0 24380 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_258
timestamp 1623621585
transform 1 0 24840 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_270
timestamp 1623621585
transform 1 0 25944 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0665_
timestamp 1623621585
transform 1 0 26220 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1623621585
transform 1 0 26956 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0506_
timestamp 1623621585
transform 1 0 28520 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_293
timestamp 1623621585
transform 1 0 28060 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_297
timestamp 1623621585
transform 1 0 28428 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_306
timestamp 1623621585
transform 1 0 29256 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1623621585
transform 1 0 29992 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_315
timestamp 1623621585
transform 1 0 30084 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_327
timestamp 1623621585
transform 1 0 31188 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_339
timestamp 1623621585
transform 1 0 32292 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_351
timestamp 1623621585
transform 1 0 33396 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1623621585
transform 1 0 35236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_363
timestamp 1623621585
transform 1 0 34500 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_372
timestamp 1623621585
transform 1 0 35328 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0702_
timestamp 1623621585
transform 1 0 36800 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1623621585
transform 1 0 36156 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_380
timestamp 1623621585
transform 1 0 36064 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_384
timestamp 1623621585
transform 1 0 36432 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_392
timestamp 1623621585
transform 1 0 37168 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0649_
timestamp 1623621585
transform 1 0 37536 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1623621585
transform -1 0 38824 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1623621585
transform 1 0 38180 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1623621585
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1623621585
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input368
timestamp 1623621585
transform 1 0 1748 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1623621585
transform 1 0 1380 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_11
timestamp 1623621585
transform 1 0 2116 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1623621585
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1623621585
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1623621585
transform 1 0 3772 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_23
timestamp 1623621585
transform 1 0 3220 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_35
timestamp 1623621585
transform 1 0 4324 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_27
timestamp 1623621585
transform 1 0 3588 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1623621585
transform 1 0 3864 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1623621585
transform 1 0 6348 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_47
timestamp 1623621585
transform 1 0 5428 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_55
timestamp 1623621585
transform 1 0 6164 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_58
timestamp 1623621585
transform 1 0 6440 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1623621585
transform 1 0 4968 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_54
timestamp 1623621585
transform 1 0 6072 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_70
timestamp 1623621585
transform 1 0 7544 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_82
timestamp 1623621585
transform 1 0 8648 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_66
timestamp 1623621585
transform 1 0 7176 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_78
timestamp 1623621585
transform 1 0 8280 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1623621585
transform 1 0 9016 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_94
timestamp 1623621585
transform 1 0 9752 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_87
timestamp 1623621585
transform 1 0 9108 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_99
timestamp 1623621585
transform 1 0 10212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1623621585
transform 1 0 11592 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_106
timestamp 1623621585
transform 1 0 10856 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_115
timestamp 1623621585
transform 1 0 11684 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_111
timestamp 1623621585
transform 1 0 11316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_123
timestamp 1623621585
transform 1 0 12420 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1623621585
transform 1 0 14260 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_127
timestamp 1623621585
transform 1 0 12788 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_139
timestamp 1623621585
transform 1 0 13892 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_135
timestamp 1623621585
transform 1 0 13524 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_144
timestamp 1623621585
transform 1 0 14352 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_151
timestamp 1623621585
transform 1 0 14996 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_163
timestamp 1623621585
transform 1 0 16100 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_156
timestamp 1623621585
transform 1 0 15456 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1623621585
transform 1 0 16836 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_172
timestamp 1623621585
transform 1 0 16928 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_184
timestamp 1623621585
transform 1 0 18032 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_168
timestamp 1623621585
transform 1 0 16560 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_180
timestamp 1623621585
transform 1 0 17664 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1623621585
transform 1 0 19504 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_196
timestamp 1623621585
transform 1 0 19136 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_208
timestamp 1623621585
transform 1 0 20240 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_192
timestamp 1623621585
transform 1 0 18768 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_201
timestamp 1623621585
transform 1 0 19596 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0458_
timestamp 1623621585
transform 1 0 21620 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1623621585
transform 1 0 22080 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_220
timestamp 1623621585
transform 1 0 21344 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_229
timestamp 1623621585
transform 1 0 22172 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_213
timestamp 1623621585
transform 1 0 20700 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_221
timestamp 1623621585
transform 1 0 21436 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _0418_
timestamp 1623621585
transform 1 0 23000 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0423_
timestamp 1623621585
transform 1 0 22540 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1623621585
transform 1 0 23828 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_241
timestamp 1623621585
transform 1 0 23276 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_231
timestamp 1623621585
transform 1 0 22356 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_237
timestamp 1623621585
transform 1 0 22908 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1623621585
transform 1 0 23644 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0414_
timestamp 1623621585
transform 1 0 25208 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1623621585
transform 1 0 24748 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_263
timestamp 1623621585
transform 1 0 25300 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_258
timestamp 1623621585
transform 1 0 24840 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_265
timestamp 1623621585
transform 1 0 25484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0656_
timestamp 1623621585
transform 1 0 26220 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1623621585
transform 1 0 27324 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_271
timestamp 1623621585
transform 1 0 26036 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_281
timestamp 1623621585
transform 1 0 26956 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_286
timestamp 1623621585
transform 1 0 27416 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_277
timestamp 1623621585
transform 1 0 26588 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_289
timestamp 1623621585
transform 1 0 27692 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _0498_
timestamp 1623621585
transform 1 0 28704 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0708_
timestamp 1623621585
transform 1 0 28520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0709_
timestamp 1623621585
transform 1 0 29256 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_298
timestamp 1623621585
transform 1 0 28520 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_308
timestamp 1623621585
transform 1 0 29440 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_297
timestamp 1623621585
transform 1 0 28428 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_302
timestamp 1623621585
transform 1 0 28888 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_310
timestamp 1623621585
transform 1 0 29624 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1623621585
transform 1 0 29992 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_320
timestamp 1623621585
transform 1 0 30544 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_332
timestamp 1623621585
transform 1 0 31648 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_315
timestamp 1623621585
transform 1 0 30084 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_327
timestamp 1623621585
transform 1 0 31188 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1623621585
transform 1 0 32568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_340
timestamp 1623621585
transform 1 0 32384 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_343
timestamp 1623621585
transform 1 0 32660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_339
timestamp 1623621585
transform 1 0 32292 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_351
timestamp 1623621585
transform 1 0 33396 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_363
timestamp 1623621585
transform 1 0 34500 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_363
timestamp 1623621585
transform 1 0 34500 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_355
timestamp 1623621585
transform 1 0 33764 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_367
timestamp 1623621585
transform 1 0 34868 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_369
timestamp 1623621585
transform 1 0 35052 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input181
timestamp 1623621585
transform 1 0 34592 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1623621585
transform 1 0 34776 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1623621585
transform 1 0 35236 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_372
timestamp 1623621585
transform 1 0 35328 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1623621585
transform 1 0 35420 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0477_
timestamp 1623621585
transform 1 0 36064 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0635_
timestamp 1623621585
transform 1 0 36248 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0766_
timestamp 1623621585
transform 1 0 36800 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_66_376
timestamp 1623621585
transform 1 0 35696 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_384
timestamp 1623621585
transform 1 0 36432 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_395
timestamp 1623621585
transform 1 0 37444 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_380
timestamp 1623621585
transform 1 0 36064 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_390
timestamp 1623621585
transform 1 0 36984 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0750_
timestamp 1623621585
transform 1 0 37536 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1623621585
transform -1 0 38824 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1623621585
transform -1 0 38824 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1623621585
transform 1 0 37812 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_400
timestamp 1623621585
transform 1 0 37904 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_406
timestamp 1623621585
transform 1 0 38456 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_403
timestamp 1623621585
transform 1 0 38180 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1623621585
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input369
timestamp 1623621585
transform 1 0 1748 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_3
timestamp 1623621585
transform 1 0 1380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_11
timestamp 1623621585
transform 1 0 2116 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_23
timestamp 1623621585
transform 1 0 3220 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_35
timestamp 1623621585
transform 1 0 4324 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1623621585
transform 1 0 6348 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_47
timestamp 1623621585
transform 1 0 5428 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_55
timestamp 1623621585
transform 1 0 6164 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_58
timestamp 1623621585
transform 1 0 6440 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_70
timestamp 1623621585
transform 1 0 7544 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_82
timestamp 1623621585
transform 1 0 8648 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_94
timestamp 1623621585
transform 1 0 9752 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1623621585
transform 1 0 11592 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_106
timestamp 1623621585
transform 1 0 10856 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_115
timestamp 1623621585
transform 1 0 11684 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_127
timestamp 1623621585
transform 1 0 12788 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_139
timestamp 1623621585
transform 1 0 13892 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_151
timestamp 1623621585
transform 1 0 14996 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_163
timestamp 1623621585
transform 1 0 16100 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1623621585
transform 1 0 16836 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_172
timestamp 1623621585
transform 1 0 16928 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_184
timestamp 1623621585
transform 1 0 18032 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_196
timestamp 1623621585
transform 1 0 19136 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_208
timestamp 1623621585
transform 1 0 20240 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1623621585
transform 1 0 22080 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_220
timestamp 1623621585
transform 1 0 21344 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_229
timestamp 1623621585
transform 1 0 22172 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_241
timestamp 1623621585
transform 1 0 23276 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1623621585
transform 1 0 24380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1623621585
transform 1 0 25484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1623621585
transform 1 0 27324 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_277
timestamp 1623621585
transform 1 0 26588 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_286
timestamp 1623621585
transform 1 0 27416 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_2  _1009_
timestamp 1623621585
transform 1 0 28152 0 -1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_68_311
timestamp 1623621585
transform 1 0 29716 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_2  _1010_
timestamp 1623621585
transform 1 0 30084 0 -1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_68_332
timestamp 1623621585
transform 1 0 31648 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1623621585
transform 1 0 32568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_340
timestamp 1623621585
transform 1 0 32384 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_343
timestamp 1623621585
transform 1 0 32660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0593_
timestamp 1623621585
transform 1 0 34868 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0646_
timestamp 1623621585
transform 1 0 35512 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1623621585
transform 1 0 34224 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_355
timestamp 1623621585
transform 1 0 33764 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_359
timestamp 1623621585
transform 1 0 34132 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_363
timestamp 1623621585
transform 1 0 34500 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_370
timestamp 1623621585
transform 1 0 35144 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0626_
timestamp 1623621585
transform 1 0 36248 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_378
timestamp 1623621585
transform 1 0 35880 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_390
timestamp 1623621585
transform 1 0 36984 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1623621585
transform -1 0 38824 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1623621585
transform 1 0 37812 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_398
timestamp 1623621585
transform 1 0 37720 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_400
timestamp 1623621585
transform 1 0 37904 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_406
timestamp 1623621585
transform 1 0 38456 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1623621585
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input370
timestamp 1623621585
transform 1 0 1748 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1623621585
transform 1 0 1380 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_11
timestamp 1623621585
transform 1 0 2116 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1623621585
transform 1 0 3772 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_23
timestamp 1623621585
transform 1 0 3220 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1623621585
transform 1 0 3864 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1623621585
transform 1 0 4968 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_54
timestamp 1623621585
transform 1 0 6072 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1623621585
transform 1 0 8004 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_69_66
timestamp 1623621585
transform 1 0 7176 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_74
timestamp 1623621585
transform 1 0 7912 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_80
timestamp 1623621585
transform 1 0 8464 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1623621585
transform 1 0 9016 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_87
timestamp 1623621585
transform 1 0 9108 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_99
timestamp 1623621585
transform 1 0 10212 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_111
timestamp 1623621585
transform 1 0 11316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_123
timestamp 1623621585
transform 1 0 12420 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1623621585
transform 1 0 14260 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_135
timestamp 1623621585
transform 1 0 13524 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_144
timestamp 1623621585
transform 1 0 14352 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_156
timestamp 1623621585
transform 1 0 15456 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_168
timestamp 1623621585
transform 1 0 16560 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_180
timestamp 1623621585
transform 1 0 17664 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1623621585
transform 1 0 19504 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_192
timestamp 1623621585
transform 1 0 18768 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_201
timestamp 1623621585
transform 1 0 19596 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_213
timestamp 1623621585
transform 1 0 20700 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1623621585
transform 1 0 21804 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1623621585
transform 1 0 22908 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_249
timestamp 1623621585
transform 1 0 24012 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1623621585
transform 1 0 24748 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_258
timestamp 1623621585
transform 1 0 24840 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_270
timestamp 1623621585
transform 1 0 25944 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_282
timestamp 1623621585
transform 1 0 27048 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_290
timestamp 1623621585
transform 1 0 27784 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  _1012_
timestamp 1623621585
transform 1 0 28060 0 1 39712
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_69_310
timestamp 1623621585
transform 1 0 29624 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1623621585
transform 1 0 29992 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_315
timestamp 1623621585
transform 1 0 30084 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_327
timestamp 1623621585
transform 1 0 31188 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_339
timestamp 1623621585
transform 1 0 32292 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_351
timestamp 1623621585
transform 1 0 33396 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1623621585
transform 1 0 35236 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input183
timestamp 1623621585
transform 1 0 34592 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_363
timestamp 1623621585
transform 1 0 34500 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_367
timestamp 1623621585
transform 1 0 34868 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_372
timestamp 1623621585
transform 1 0 35328 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0618_
timestamp 1623621585
transform 1 0 36248 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_380
timestamp 1623621585
transform 1 0 36064 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_390
timestamp 1623621585
transform 1 0 36984 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0758_
timestamp 1623621585
transform 1 0 37536 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1623621585
transform -1 0 38824 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_403
timestamp 1623621585
transform 1 0 38180 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1623621585
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1623621585
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1623621585
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_27
timestamp 1623621585
transform 1 0 3588 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_39
timestamp 1623621585
transform 1 0 4692 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1623621585
transform 1 0 6348 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_51
timestamp 1623621585
transform 1 0 5796 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_58
timestamp 1623621585
transform 1 0 6440 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0740_
timestamp 1623621585
transform 1 0 7820 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1623621585
transform 1 0 8648 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_70_70
timestamp 1623621585
transform 1 0 7544 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_78
timestamp 1623621585
transform 1 0 8280 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_87
timestamp 1623621585
transform 1 0 9108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_99
timestamp 1623621585
transform 1 0 10212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1623621585
transform 1 0 11592 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_111
timestamp 1623621585
transform 1 0 11316 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_115
timestamp 1623621585
transform 1 0 11684 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_127
timestamp 1623621585
transform 1 0 12788 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_139
timestamp 1623621585
transform 1 0 13892 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_151
timestamp 1623621585
transform 1 0 14996 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_163
timestamp 1623621585
transform 1 0 16100 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1623621585
transform 1 0 16836 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_172
timestamp 1623621585
transform 1 0 16928 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_184
timestamp 1623621585
transform 1 0 18032 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_196
timestamp 1623621585
transform 1 0 19136 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_208
timestamp 1623621585
transform 1 0 20240 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1623621585
transform 1 0 22080 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_220
timestamp 1623621585
transform 1 0 21344 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_229
timestamp 1623621585
transform 1 0 22172 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1013_
timestamp 1623621585
transform 1 0 22540 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0420_
timestamp 1623621585
transform 1 0 24656 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_252
timestamp 1623621585
transform 1 0 24288 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_260
timestamp 1623621585
transform 1 0 25024 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1623621585
transform 1 0 27324 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_272
timestamp 1623621585
transform 1 0 26128 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_284
timestamp 1623621585
transform 1 0 27232 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_286
timestamp 1623621585
transform 1 0 27416 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1011_
timestamp 1623621585
transform 1 0 28704 0 -1 40800
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_70_298
timestamp 1623621585
transform 1 0 28520 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_317
timestamp 1623621585
transform 1 0 30268 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_329
timestamp 1623621585
transform 1 0 31372 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1623621585
transform 1 0 32568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_341
timestamp 1623621585
transform 1 0 32476 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_343
timestamp 1623621585
transform 1 0 32660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1623621585
transform 1 0 35604 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1623621585
transform 1 0 34960 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_355
timestamp 1623621585
transform 1 0 33764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_367
timestamp 1623621585
transform 1 0 34868 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_371
timestamp 1623621585
transform 1 0 35236 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0596_
timestamp 1623621585
transform 1 0 36248 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_378
timestamp 1623621585
transform 1 0 35880 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_390
timestamp 1623621585
transform 1 0 36984 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1623621585
transform -1 0 38824 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1623621585
transform 1 0 37812 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_398
timestamp 1623621585
transform 1 0 37720 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_400
timestamp 1623621585
transform 1 0 37904 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_406
timestamp 1623621585
transform 1 0 38456 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1623621585
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input371
timestamp 1623621585
transform 1 0 1748 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1623621585
transform 1 0 1380 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_11
timestamp 1623621585
transform 1 0 2116 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1623621585
transform 1 0 3772 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_23
timestamp 1623621585
transform 1 0 3220 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1623621585
transform 1 0 3864 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1623621585
transform 1 0 4968 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_54
timestamp 1623621585
transform 1 0 6072 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0731_
timestamp 1623621585
transform 1 0 7820 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_71_66
timestamp 1623621585
transform 1 0 7176 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_72
timestamp 1623621585
transform 1 0 7728 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_78
timestamp 1623621585
transform 1 0 8280 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1623621585
transform 1 0 9476 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1623621585
transform 1 0 9016 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_87
timestamp 1623621585
transform 1 0 9108 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_96
timestamp 1623621585
transform 1 0 9936 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_108
timestamp 1623621585
transform 1 0 11040 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_120
timestamp 1623621585
transform 1 0 12144 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1623621585
transform 1 0 14260 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_132
timestamp 1623621585
transform 1 0 13248 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_140
timestamp 1623621585
transform 1 0 13984 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_144
timestamp 1623621585
transform 1 0 14352 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_156
timestamp 1623621585
transform 1 0 15456 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_168
timestamp 1623621585
transform 1 0 16560 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_180
timestamp 1623621585
transform 1 0 17664 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1623621585
transform 1 0 19504 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_192
timestamp 1623621585
transform 1 0 18768 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_201
timestamp 1623621585
transform 1 0 19596 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_213
timestamp 1623621585
transform 1 0 20700 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1623621585
transform 1 0 21804 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1623621585
transform 1 0 22908 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1623621585
transform 1 0 24012 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1623621585
transform 1 0 24748 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_258
timestamp 1623621585
transform 1 0 24840 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_270
timestamp 1623621585
transform 1 0 25944 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0636_
timestamp 1623621585
transform 1 0 26496 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_284
timestamp 1623621585
transform 1 0 27232 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0655_
timestamp 1623621585
transform 1 0 28612 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_71_296
timestamp 1623621585
transform 1 0 28336 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_303
timestamp 1623621585
transform 1 0 28980 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_311
timestamp 1623621585
transform 1 0 29716 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1623621585
transform 1 0 29992 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_315
timestamp 1623621585
transform 1 0 30084 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_327
timestamp 1623621585
transform 1 0 31188 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_339
timestamp 1623621585
transform 1 0 32292 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_351
timestamp 1623621585
transform 1 0 33396 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1623621585
transform 1 0 35236 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input184
timestamp 1623621585
transform 1 0 34592 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_363
timestamp 1623621585
transform 1 0 34500 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_367
timestamp 1623621585
transform 1 0 34868 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_372
timestamp 1623621585
transform 1 0 35328 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0610_
timestamp 1623621585
transform 1 0 36248 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_380
timestamp 1623621585
transform 1 0 36064 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_390
timestamp 1623621585
transform 1 0 36984 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0634_
timestamp 1623621585
transform 1 0 37536 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1623621585
transform -1 0 38824 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_403
timestamp 1623621585
transform 1 0 38180 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1623621585
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1623621585
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input372
timestamp 1623621585
transform 1 0 1748 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_3
timestamp 1623621585
transform 1 0 1380 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_11
timestamp 1623621585
transform 1 0 2116 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1623621585
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1623621585
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1623621585
transform 1 0 3772 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_23
timestamp 1623621585
transform 1 0 3220 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_35
timestamp 1623621585
transform 1 0 4324 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1623621585
transform 1 0 3588 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_30
timestamp 1623621585
transform 1 0 3864 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1623621585
transform 1 0 6348 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_47
timestamp 1623621585
transform 1 0 5428 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_55
timestamp 1623621585
transform 1 0 6164 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_58
timestamp 1623621585
transform 1 0 6440 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_42
timestamp 1623621585
transform 1 0 4968 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_54
timestamp 1623621585
transform 1 0 6072 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1623621585
transform 1 0 7912 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1623621585
transform 1 0 8740 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0723_
timestamp 1623621585
transform 1 0 7912 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_72_70
timestamp 1623621585
transform 1 0 7544 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_79
timestamp 1623621585
transform 1 0 8372 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_66
timestamp 1623621585
transform 1 0 7176 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_79
timestamp 1623621585
transform 1 0 8372 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1623621585
transform 1 0 9016 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_88
timestamp 1623621585
transform 1 0 9200 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_100
timestamp 1623621585
transform 1 0 10304 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_85
timestamp 1623621585
transform 1 0 8924 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_87
timestamp 1623621585
transform 1 0 9108 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_99
timestamp 1623621585
transform 1 0 10212 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1623621585
transform 1 0 11592 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_112
timestamp 1623621585
transform 1 0 11408 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_115
timestamp 1623621585
transform 1 0 11684 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_111
timestamp 1623621585
transform 1 0 11316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1623621585
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1623621585
transform 1 0 14260 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_127
timestamp 1623621585
transform 1 0 12788 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_139
timestamp 1623621585
transform 1 0 13892 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_135
timestamp 1623621585
transform 1 0 13524 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_144
timestamp 1623621585
transform 1 0 14352 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_151
timestamp 1623621585
transform 1 0 14996 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_163
timestamp 1623621585
transform 1 0 16100 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_156
timestamp 1623621585
transform 1 0 15456 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1623621585
transform 1 0 16836 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_172
timestamp 1623621585
transform 1 0 16928 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_184
timestamp 1623621585
transform 1 0 18032 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_168
timestamp 1623621585
transform 1 0 16560 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_180
timestamp 1623621585
transform 1 0 17664 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1623621585
transform 1 0 19504 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_196
timestamp 1623621585
transform 1 0 19136 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_208
timestamp 1623621585
transform 1 0 20240 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_192
timestamp 1623621585
transform 1 0 18768 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_201
timestamp 1623621585
transform 1 0 19596 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1623621585
transform 1 0 22080 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_220
timestamp 1623621585
transform 1 0 21344 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_229
timestamp 1623621585
transform 1 0 22172 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_213
timestamp 1623621585
transform 1 0 20700 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1623621585
transform 1 0 21804 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_241
timestamp 1623621585
transform 1 0 23276 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1623621585
transform 1 0 22908 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_249
timestamp 1623621585
transform 1 0 24012 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0546_
timestamp 1623621585
transform 1 0 25760 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1623621585
transform 1 0 24748 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1623621585
transform 1 0 24380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1623621585
transform 1 0 25484 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_258
timestamp 1623621585
transform 1 0 24840 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_266
timestamp 1623621585
transform 1 0 25576 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0547_
timestamp 1623621585
transform 1 0 26496 0 1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _0619_
timestamp 1623621585
transform 1 0 27784 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0628_
timestamp 1623621585
transform 1 0 26220 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1623621585
transform 1 0 27324 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_281
timestamp 1623621585
transform 1 0 26956 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_286
timestamp 1623621585
transform 1 0 27416 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_272
timestamp 1623621585
transform 1 0 26128 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_286
timestamp 1623621585
transform 1 0 27416 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0489_
timestamp 1623621585
transform 1 0 28704 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0491_
timestamp 1623621585
transform 1 0 29440 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0654_
timestamp 1623621585
transform 1 0 28888 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_298
timestamp 1623621585
transform 1 0 28520 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1623621585
transform 1 0 29072 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_312
timestamp 1623621585
transform 1 0 29808 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_298
timestamp 1623621585
transform 1 0 28520 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_306
timestamp 1623621585
transform 1 0 29256 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1623621585
transform 1 0 29992 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_324
timestamp 1623621585
transform 1 0 30912 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_315
timestamp 1623621585
transform 1 0 30084 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_327
timestamp 1623621585
transform 1 0 31188 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1623621585
transform 1 0 32568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_336
timestamp 1623621585
transform 1 0 32016 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_343
timestamp 1623621585
transform 1 0 32660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_339
timestamp 1623621585
transform 1 0 32292 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_351
timestamp 1623621585
transform 1 0 33396 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_363
timestamp 1623621585
transform 1 0 34500 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1623621585
transform 1 0 34500 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_355
timestamp 1623621585
transform 1 0 33764 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_367
timestamp 1623621585
transform 1 0 34868 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_367
timestamp 1623621585
transform 1 0 34868 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1623621585
transform 1 0 34592 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1623621585
transform 1 0 34592 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1623621585
transform 1 0 35236 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1623621585
transform 1 0 35236 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_372
timestamp 1623621585
transform 1 0 35328 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_374
timestamp 1623621585
transform 1 0 35512 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0475_
timestamp 1623621585
transform 1 0 36616 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0537_
timestamp 1623621585
transform 1 0 35880 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0625_
timestamp 1623621585
transform 1 0 36248 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0648_
timestamp 1623621585
transform 1 0 37260 0 1 41888
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_72_382
timestamp 1623621585
transform 1 0 36248 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_390
timestamp 1623621585
transform 1 0 36984 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_380
timestamp 1623621585
transform 1 0 36064 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_389
timestamp 1623621585
transform 1 0 36892 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1623621585
transform -1 0 38824 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1623621585
transform -1 0 38824 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1623621585
transform 1 0 37812 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_398
timestamp 1623621585
transform 1 0 37720 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_400
timestamp 1623621585
transform 1 0 37904 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_406
timestamp 1623621585
transform 1 0 38456 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_403
timestamp 1623621585
transform 1 0 38180 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1623621585
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input373
timestamp 1623621585
transform 1 0 1748 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_3
timestamp 1623621585
transform 1 0 1380 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_11
timestamp 1623621585
transform 1 0 2116 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_23
timestamp 1623621585
transform 1 0 3220 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_35
timestamp 1623621585
transform 1 0 4324 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1623621585
transform 1 0 6348 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_47
timestamp 1623621585
transform 1 0 5428 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_55
timestamp 1623621585
transform 1 0 6164 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_58
timestamp 1623621585
transform 1 0 6440 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_70
timestamp 1623621585
transform 1 0 7544 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_82
timestamp 1623621585
transform 1 0 8648 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_94
timestamp 1623621585
transform 1 0 9752 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1623621585
transform 1 0 11592 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_106
timestamp 1623621585
transform 1 0 10856 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_115
timestamp 1623621585
transform 1 0 11684 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_127
timestamp 1623621585
transform 1 0 12788 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_139
timestamp 1623621585
transform 1 0 13892 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_151
timestamp 1623621585
transform 1 0 14996 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_163
timestamp 1623621585
transform 1 0 16100 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1623621585
transform 1 0 16836 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_172
timestamp 1623621585
transform 1 0 16928 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_184
timestamp 1623621585
transform 1 0 18032 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_196
timestamp 1623621585
transform 1 0 19136 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_208
timestamp 1623621585
transform 1 0 20240 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1623621585
transform 1 0 22080 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_220
timestamp 1623621585
transform 1 0 21344 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_229
timestamp 1623621585
transform 1 0 22172 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_241
timestamp 1623621585
transform 1 0 23276 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1623621585
transform 1 0 24380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1623621585
transform 1 0 25484 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0611_
timestamp 1623621585
transform 1 0 26220 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1623621585
transform 1 0 27324 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_281
timestamp 1623621585
transform 1 0 26956 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_286
timestamp 1623621585
transform 1 0 27416 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_298
timestamp 1623621585
transform 1 0 28520 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_310
timestamp 1623621585
transform 1 0 29624 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_322
timestamp 1623621585
transform 1 0 30728 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1623621585
transform 1 0 32568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_334
timestamp 1623621585
transform 1 0 31832 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_343
timestamp 1623621585
transform 1 0 32660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1623621585
transform 1 0 35512 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input185
timestamp 1623621585
transform 1 0 34868 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_355
timestamp 1623621585
transform 1 0 33764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_370
timestamp 1623621585
transform 1 0 35144 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0592_
timestamp 1623621585
transform 1 0 36156 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0617_
timestamp 1623621585
transform 1 0 36800 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_74_377
timestamp 1623621585
transform 1 0 35788 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_384
timestamp 1623621585
transform 1 0 36432 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_395
timestamp 1623621585
transform 1 0 37444 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1623621585
transform -1 0 38824 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1623621585
transform 1 0 37812 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_400
timestamp 1623621585
transform 1 0 37904 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_406
timestamp 1623621585
transform 1 0 38456 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1623621585
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input375
timestamp 1623621585
transform 1 0 1748 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_3
timestamp 1623621585
transform 1 0 1380 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_11
timestamp 1623621585
transform 1 0 2116 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1623621585
transform 1 0 3772 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_23
timestamp 1623621585
transform 1 0 3220 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1623621585
transform 1 0 3864 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1623621585
transform 1 0 4968 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_54
timestamp 1623621585
transform 1 0 6072 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_66
timestamp 1623621585
transform 1 0 7176 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_78
timestamp 1623621585
transform 1 0 8280 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1623621585
transform 1 0 9016 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_87
timestamp 1623621585
transform 1 0 9108 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_99
timestamp 1623621585
transform 1 0 10212 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_111
timestamp 1623621585
transform 1 0 11316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_123
timestamp 1623621585
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1623621585
transform 1 0 14260 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_135
timestamp 1623621585
transform 1 0 13524 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_144
timestamp 1623621585
transform 1 0 14352 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_156
timestamp 1623621585
transform 1 0 15456 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_168
timestamp 1623621585
transform 1 0 16560 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_180
timestamp 1623621585
transform 1 0 17664 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1623621585
transform 1 0 19504 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_192
timestamp 1623621585
transform 1 0 18768 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_201
timestamp 1623621585
transform 1 0 19596 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_213
timestamp 1623621585
transform 1 0 20700 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1623621585
transform 1 0 21804 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1623621585
transform 1 0 22908 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1623621585
transform 1 0 24012 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1623621585
transform 1 0 24748 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_258
timestamp 1623621585
transform 1 0 24840 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_270
timestamp 1623621585
transform 1 0 25944 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0602_
timestamp 1623621585
transform 1 0 26496 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_284
timestamp 1623621585
transform 1 0 27232 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0464_
timestamp 1623621585
transform 1 0 28888 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_75_296
timestamp 1623621585
transform 1 0 28336 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_310
timestamp 1623621585
transform 1 0 29624 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1623621585
transform 1 0 29992 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_315
timestamp 1623621585
transform 1 0 30084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_327
timestamp 1623621585
transform 1 0 31188 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_339
timestamp 1623621585
transform 1 0 32292 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_351
timestamp 1623621585
transform 1 0 33396 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1623621585
transform 1 0 35236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input153
timestamp 1623621585
transform 1 0 34592 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_363
timestamp 1623621585
transform 1 0 34500 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_367
timestamp 1623621585
transform 1 0 34868 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_372
timestamp 1623621585
transform 1 0 35328 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0424_
timestamp 1623621585
transform 1 0 35696 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0474_
timestamp 1623621585
transform 1 0 36616 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_380
timestamp 1623621585
transform 1 0 36064 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_75_390
timestamp 1623621585
transform 1 0 36984 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0609_
timestamp 1623621585
transform 1 0 37536 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1623621585
transform -1 0 38824 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1623621585
transform 1 0 38180 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1623621585
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1623621585
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1623621585
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_27
timestamp 1623621585
transform 1 0 3588 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_39
timestamp 1623621585
transform 1 0 4692 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1623621585
transform 1 0 6348 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_51
timestamp 1623621585
transform 1 0 5796 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_58
timestamp 1623621585
transform 1 0 6440 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp 1623621585
transform 1 0 8188 0 -1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_76_70
timestamp 1623621585
transform 1 0 7544 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_76
timestamp 1623621585
transform 1 0 8096 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_82
timestamp 1623621585
transform 1 0 8648 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1623621585
transform 1 0 9016 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_89
timestamp 1623621585
transform 1 0 9292 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_101
timestamp 1623621585
transform 1 0 10396 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1623621585
transform 1 0 11592 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_113
timestamp 1623621585
transform 1 0 11500 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_115
timestamp 1623621585
transform 1 0 11684 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_127
timestamp 1623621585
transform 1 0 12788 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_139
timestamp 1623621585
transform 1 0 13892 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_151
timestamp 1623621585
transform 1 0 14996 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_163
timestamp 1623621585
transform 1 0 16100 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1623621585
transform 1 0 16836 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_172
timestamp 1623621585
transform 1 0 16928 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_184
timestamp 1623621585
transform 1 0 18032 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_196
timestamp 1623621585
transform 1 0 19136 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_208
timestamp 1623621585
transform 1 0 20240 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1623621585
transform 1 0 22080 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_220
timestamp 1623621585
transform 1 0 21344 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_229
timestamp 1623621585
transform 1 0 22172 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_241
timestamp 1623621585
transform 1 0 23276 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1623621585
transform 1 0 24380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1623621585
transform 1 0 25484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1623621585
transform 1 0 27324 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_277
timestamp 1623621585
transform 1 0 26588 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_286
timestamp 1623621585
transform 1 0 27416 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0456_
timestamp 1623621585
transform 1 0 29348 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_298
timestamp 1623621585
transform 1 0 28520 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_306
timestamp 1623621585
transform 1 0 29256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_315
timestamp 1623621585
transform 1 0 30084 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_327
timestamp 1623621585
transform 1 0 31188 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1623621585
transform 1 0 32568 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_339
timestamp 1623621585
transform 1 0 32292 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_343
timestamp 1623621585
transform 1 0 32660 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input186
timestamp 1623621585
transform 1 0 35052 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_355
timestamp 1623621585
transform 1 0 33764 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_367
timestamp 1623621585
transform 1 0 34868 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_372
timestamp 1623621585
transform 1 0 35328 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0581_
timestamp 1623621585
transform 1 0 36340 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1623621585
transform 1 0 35696 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_379
timestamp 1623621585
transform 1 0 35972 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_391
timestamp 1623621585
transform 1 0 37076 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1623621585
transform -1 0 38824 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1623621585
transform 1 0 37812 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_400
timestamp 1623621585
transform 1 0 37904 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_406
timestamp 1623621585
transform 1 0 38456 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1623621585
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input376
timestamp 1623621585
transform 1 0 1748 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1623621585
transform 1 0 1380 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_11
timestamp 1623621585
transform 1 0 2116 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1623621585
transform 1 0 3772 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_23
timestamp 1623621585
transform 1 0 3220 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_30
timestamp 1623621585
transform 1 0 3864 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1623621585
transform 1 0 4968 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_54
timestamp 1623621585
transform 1 0 6072 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0661_
timestamp 1623621585
transform 1 0 8188 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0677_
timestamp 1623621585
transform 1 0 7360 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_77_66
timestamp 1623621585
transform 1 0 7176 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_73
timestamp 1623621585
transform 1 0 7820 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_82
timestamp 1623621585
transform 1 0 8648 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1623621585
transform 1 0 9476 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1623621585
transform 1 0 9016 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_87
timestamp 1623621585
transform 1 0 9108 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_96
timestamp 1623621585
transform 1 0 9936 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_108
timestamp 1623621585
transform 1 0 11040 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_120
timestamp 1623621585
transform 1 0 12144 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1623621585
transform 1 0 14260 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_132
timestamp 1623621585
transform 1 0 13248 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_140
timestamp 1623621585
transform 1 0 13984 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_144
timestamp 1623621585
transform 1 0 14352 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_156
timestamp 1623621585
transform 1 0 15456 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_168
timestamp 1623621585
transform 1 0 16560 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_180
timestamp 1623621585
transform 1 0 17664 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1623621585
transform 1 0 19504 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_192
timestamp 1623621585
transform 1 0 18768 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_201
timestamp 1623621585
transform 1 0 19596 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_213
timestamp 1623621585
transform 1 0 20700 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1623621585
transform 1 0 21804 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1623621585
transform 1 0 22908 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_249
timestamp 1623621585
transform 1 0 24012 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1623621585
transform 1 0 24748 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_258
timestamp 1623621585
transform 1 0 24840 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_270
timestamp 1623621585
transform 1 0 25944 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0490_
timestamp 1623621585
transform 1 0 26772 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_278
timestamp 1623621585
transform 1 0 26680 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_283
timestamp 1623621585
transform 1 0 27140 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_291
timestamp 1623621585
transform 1 0 27876 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0447_
timestamp 1623621585
transform 1 0 28888 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0601_
timestamp 1623621585
transform 1 0 28152 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_298
timestamp 1623621585
transform 1 0 28520 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_310
timestamp 1623621585
transform 1 0 29624 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1623621585
transform 1 0 29992 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_315
timestamp 1623621585
transform 1 0 30084 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_327
timestamp 1623621585
transform 1 0 31188 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_339
timestamp 1623621585
transform 1 0 32292 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_351
timestamp 1623621585
transform 1 0 33396 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1623621585
transform 1 0 35236 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1623621585
transform 1 0 34592 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_363
timestamp 1623621585
transform 1 0 34500 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_367
timestamp 1623621585
transform 1 0 34868 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_372
timestamp 1623621585
transform 1 0 35328 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0476_
timestamp 1623621585
transform 1 0 35696 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0572_
timestamp 1623621585
transform 1 0 36432 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_380
timestamp 1623621585
transform 1 0 36064 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_392
timestamp 1623621585
transform 1 0 37168 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0595_
timestamp 1623621585
transform 1 0 37536 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1623621585
transform -1 0 38824 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_403
timestamp 1623621585
transform 1 0 38180 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1623621585
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input377
timestamp 1623621585
transform 1 0 1748 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1623621585
transform 1 0 1380 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_11
timestamp 1623621585
transform 1 0 2116 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_23
timestamp 1623621585
transform 1 0 3220 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_35
timestamp 1623621585
transform 1 0 4324 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1623621585
transform 1 0 6348 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_47
timestamp 1623621585
transform 1 0 5428 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_55
timestamp 1623621585
transform 1 0 6164 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_58
timestamp 1623621585
transform 1 0 6440 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0535_
timestamp 1623621585
transform 1 0 8648 0 -1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0569_
timestamp 1623621585
transform 1 0 7820 0 -1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_78_70
timestamp 1623621585
transform 1 0 7544 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_78
timestamp 1623621585
transform 1 0 8280 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0553_
timestamp 1623621585
transform 1 0 9476 0 -1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0578_
timestamp 1623621585
transform 1 0 10304 0 -1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_78_87
timestamp 1623621585
transform 1 0 9108 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_96
timestamp 1623621585
transform 1 0 9936 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1623621585
transform 1 0 11592 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_105
timestamp 1623621585
transform 1 0 10764 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_113
timestamp 1623621585
transform 1 0 11500 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_115
timestamp 1623621585
transform 1 0 11684 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_127
timestamp 1623621585
transform 1 0 12788 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_139
timestamp 1623621585
transform 1 0 13892 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_151
timestamp 1623621585
transform 1 0 14996 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_163
timestamp 1623621585
transform 1 0 16100 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1623621585
transform 1 0 16836 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_172
timestamp 1623621585
transform 1 0 16928 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_184
timestamp 1623621585
transform 1 0 18032 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_196
timestamp 1623621585
transform 1 0 19136 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_208
timestamp 1623621585
transform 1 0 20240 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1623621585
transform 1 0 22080 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_220
timestamp 1623621585
transform 1 0 21344 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_229
timestamp 1623621585
transform 1 0 22172 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0419_
timestamp 1623621585
transform 1 0 24012 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_241
timestamp 1623621585
transform 1 0 23276 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1623621585
transform 1 0 24380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1623621585
transform 1 0 25484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0492_
timestamp 1623621585
transform 1 0 26588 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1623621585
transform 1 0 27324 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_281
timestamp 1623621585
transform 1 0 26956 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_286
timestamp 1623621585
transform 1 0 27416 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__o32a_1  _0439_
timestamp 1623621585
transform 1 0 29532 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0600_
timestamp 1623621585
transform 1 0 28796 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_298
timestamp 1623621585
transform 1 0 28520 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_305
timestamp 1623621585
transform 1 0 29164 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_317
timestamp 1623621585
transform 1 0 30268 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_329
timestamp 1623621585
transform 1 0 31372 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1623621585
transform 1 0 32568 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_341
timestamp 1623621585
transform 1 0 32476 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_343
timestamp 1623621585
transform 1 0 32660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0594_
timestamp 1623621585
transform 1 0 35144 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input187
timestamp 1623621585
transform 1 0 34500 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_355
timestamp 1623621585
transform 1 0 33764 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_366
timestamp 1623621585
transform 1 0 34776 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_373
timestamp 1623621585
transform 1 0 35420 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1623621585
transform 1 0 35788 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0564_
timestamp 1623621585
transform 1 0 36432 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_380
timestamp 1623621585
transform 1 0 36064 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_392
timestamp 1623621585
transform 1 0 37168 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1623621585
transform -1 0 38824 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1623621585
transform 1 0 37812 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_398
timestamp 1623621585
transform 1 0 37720 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_400
timestamp 1623621585
transform 1 0 37904 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_406
timestamp 1623621585
transform 1 0 38456 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1623621585
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1623621585
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input378
timestamp 1623621585
transform 1 0 1748 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1623621585
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1623621585
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_3
timestamp 1623621585
transform 1 0 1380 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_11
timestamp 1623621585
transform 1 0 2116 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1623621585
transform 1 0 3772 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_27
timestamp 1623621585
transform 1 0 3588 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1623621585
transform 1 0 3864 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_23
timestamp 1623621585
transform 1 0 3220 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_35
timestamp 1623621585
transform 1 0 4324 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1623621585
transform 1 0 6348 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1623621585
transform 1 0 4968 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_54
timestamp 1623621585
transform 1 0 6072 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_47
timestamp 1623621585
transform 1 0 5428 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_55
timestamp 1623621585
transform 1 0 6164 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_58
timestamp 1623621585
transform 1 0 6440 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0470_
timestamp 1623621585
transform 1 0 7544 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0643_
timestamp 1623621585
transform 1 0 8188 0 1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_79_66
timestamp 1623621585
transform 1 0 7176 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_73
timestamp 1623621585
transform 1 0 7820 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_82
timestamp 1623621585
transform 1 0 8648 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_70
timestamp 1623621585
transform 1 0 7544 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_82
timestamp 1623621585
transform 1 0 8648 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0515_
timestamp 1623621585
transform 1 0 8924 0 -1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0561_
timestamp 1623621585
transform 1 0 9476 0 1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1623621585
transform 1 0 9016 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_87
timestamp 1623621585
transform 1 0 9108 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_96
timestamp 1623621585
transform 1 0 9936 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_90
timestamp 1623621585
transform 1 0 9384 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_102
timestamp 1623621585
transform 1 0 10488 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1623621585
transform 1 0 11592 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_108
timestamp 1623621585
transform 1 0 11040 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_120
timestamp 1623621585
transform 1 0 12144 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_115
timestamp 1623621585
transform 1 0 11684 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1623621585
transform 1 0 14260 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_132
timestamp 1623621585
transform 1 0 13248 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_140
timestamp 1623621585
transform 1 0 13984 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_144
timestamp 1623621585
transform 1 0 14352 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_127
timestamp 1623621585
transform 1 0 12788 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_139
timestamp 1623621585
transform 1 0 13892 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_156
timestamp 1623621585
transform 1 0 15456 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_151
timestamp 1623621585
transform 1 0 14996 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_163
timestamp 1623621585
transform 1 0 16100 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1623621585
transform 1 0 16836 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_168
timestamp 1623621585
transform 1 0 16560 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_180
timestamp 1623621585
transform 1 0 17664 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_172
timestamp 1623621585
transform 1 0 16928 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_184
timestamp 1623621585
transform 1 0 18032 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1623621585
transform 1 0 19504 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_192
timestamp 1623621585
transform 1 0 18768 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_201
timestamp 1623621585
transform 1 0 19596 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_196
timestamp 1623621585
transform 1 0 19136 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_208
timestamp 1623621585
transform 1 0 20240 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1623621585
transform 1 0 22080 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_213
timestamp 1623621585
transform 1 0 20700 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1623621585
transform 1 0 21804 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_220
timestamp 1623621585
transform 1 0 21344 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_229
timestamp 1623621585
transform 1 0 22172 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1623621585
transform 1 0 22908 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_249
timestamp 1623621585
transform 1 0 24012 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_241
timestamp 1623621585
transform 1 0 23276 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1623621585
transform 1 0 24748 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_258
timestamp 1623621585
transform 1 0 24840 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_270
timestamp 1623621585
transform 1 0 25944 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1623621585
transform 1 0 24380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_265
timestamp 1623621585
transform 1 0 25484 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0574_
timestamp 1623621585
transform 1 0 26220 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0582_
timestamp 1623621585
transform 1 0 26312 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1623621585
transform 1 0 27324 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_282
timestamp 1623621585
transform 1 0 27048 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_281
timestamp 1623621585
transform 1 0 26956 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_286
timestamp 1623621585
transform 1 0 27416 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_294
timestamp 1623621585
transform 1 0 28152 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_306
timestamp 1623621585
transform 1 0 29256 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_298
timestamp 1623621585
transform 1 0 28520 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_310
timestamp 1623621585
transform 1 0 29624 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1623621585
transform 1 0 29992 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_315
timestamp 1623621585
transform 1 0 30084 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_327
timestamp 1623621585
transform 1 0 31188 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_322
timestamp 1623621585
transform 1 0 30728 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1623621585
transform 1 0 32568 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_339
timestamp 1623621585
transform 1 0 32292 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_351
timestamp 1623621585
transform 1 0 33396 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_334
timestamp 1623621585
transform 1 0 31832 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_343
timestamp 1623621585
transform 1 0 32660 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1623621585
transform 1 0 35236 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1623621585
transform 1 0 35236 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_363
timestamp 1623621585
transform 1 0 34500 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_372
timestamp 1623621585
transform 1 0 35328 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_355
timestamp 1623621585
transform 1 0 33764 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_367
timestamp 1623621585
transform 1 0 34868 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_374
timestamp 1623621585
transform 1 0 35512 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0540_
timestamp 1623621585
transform 1 0 35788 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _0542_
timestamp 1623621585
transform 1 0 36524 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0556_
timestamp 1623621585
transform 1 0 36432 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1623621585
transform 1 0 35880 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_79_376
timestamp 1623621585
transform 1 0 35696 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_380
timestamp 1623621585
transform 1 0 36064 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_393
timestamp 1623621585
transform 1 0 37260 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_381
timestamp 1623621585
transform 1 0 36156 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_394
timestamp 1623621585
transform 1 0 37352 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0479_
timestamp 1623621585
transform 1 0 37628 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1623621585
transform -1 0 38824 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1623621585
transform -1 0 38824 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1623621585
transform 1 0 37812 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_401
timestamp 1623621585
transform 1 0 37996 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_398
timestamp 1623621585
transform 1 0 37720 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_80_400
timestamp 1623621585
transform 1 0 37904 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_406
timestamp 1623621585
transform 1 0 38456 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1623621585
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input379
timestamp 1623621585
transform 1 0 1380 0 1 46240
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_81_13
timestamp 1623621585
transform 1 0 2300 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1623621585
transform 1 0 3772 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_25
timestamp 1623621585
transform 1 0 3404 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1623621585
transform 1 0 3864 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1623621585
transform 1 0 4968 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_54
timestamp 1623621585
transform 1 0 6072 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_62
timestamp 1623621585
transform 1 0 6808 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__and2_1  _0524_
timestamp 1623621585
transform 1 0 8188 0 1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0696_
timestamp 1623621585
transform 1 0 6992 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_67
timestamp 1623621585
transform 1 0 7268 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_75
timestamp 1623621585
transform 1 0 8004 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_82
timestamp 1623621585
transform 1 0 8648 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0471_
timestamp 1623621585
transform 1 0 9476 0 1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1623621585
transform 1 0 9016 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_87
timestamp 1623621585
transform 1 0 9108 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_96
timestamp 1623621585
transform 1 0 9936 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_108
timestamp 1623621585
transform 1 0 11040 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_120
timestamp 1623621585
transform 1 0 12144 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1623621585
transform 1 0 14260 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_132
timestamp 1623621585
transform 1 0 13248 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_140
timestamp 1623621585
transform 1 0 13984 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_144
timestamp 1623621585
transform 1 0 14352 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_156
timestamp 1623621585
transform 1 0 15456 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_168
timestamp 1623621585
transform 1 0 16560 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_180
timestamp 1623621585
transform 1 0 17664 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1623621585
transform 1 0 19504 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_192
timestamp 1623621585
transform 1 0 18768 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_201
timestamp 1623621585
transform 1 0 19596 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_213
timestamp 1623621585
transform 1 0 20700 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1623621585
transform 1 0 21804 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1623621585
transform 1 0 22908 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_249
timestamp 1623621585
transform 1 0 24012 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1623621585
transform 1 0 24748 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_258
timestamp 1623621585
transform 1 0 24840 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_270
timestamp 1623621585
transform 1 0 25944 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0565_
timestamp 1623621585
transform 1 0 26312 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_282
timestamp 1623621585
transform 1 0 27048 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_294
timestamp 1623621585
transform 1 0 28152 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_306
timestamp 1623621585
transform 1 0 29256 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1623621585
transform 1 0 29992 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_315
timestamp 1623621585
transform 1 0 30084 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_327
timestamp 1623621585
transform 1 0 31188 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_339
timestamp 1623621585
transform 1 0 32292 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_351
timestamp 1623621585
transform 1 0 33396 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1623621585
transform 1 0 35236 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_363
timestamp 1623621585
transform 1 0 34500 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_81_372
timestamp 1623621585
transform 1 0 35328 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0478_
timestamp 1623621585
transform 1 0 36800 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1623621585
transform 1 0 36156 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_380
timestamp 1623621585
transform 1 0 36064 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_384
timestamp 1623621585
transform 1 0 36432 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_392
timestamp 1623621585
transform 1 0 37168 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0580_
timestamp 1623621585
transform 1 0 37536 0 1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1623621585
transform -1 0 38824 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1623621585
transform 1 0 38180 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1623621585
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1623621585
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1623621585
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_27
timestamp 1623621585
transform 1 0 3588 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_39
timestamp 1623621585
transform 1 0 4692 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1623621585
transform 1 0 6348 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_51
timestamp 1623621585
transform 1 0 5796 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_58
timestamp 1623621585
transform 1 0 6440 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0615_
timestamp 1623621585
transform 1 0 8188 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0632_
timestamp 1623621585
transform 1 0 7360 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_82_66
timestamp 1623621585
transform 1 0 7176 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_73
timestamp 1623621585
transform 1 0 7820 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_82
timestamp 1623621585
transform 1 0 8648 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0499_
timestamp 1623621585
transform 1 0 9016 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0507_
timestamp 1623621585
transform 1 0 9844 0 -1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_82_91
timestamp 1623621585
transform 1 0 9476 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_100
timestamp 1623621585
transform 1 0 10304 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1623621585
transform 1 0 11592 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_112
timestamp 1623621585
transform 1 0 11408 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_115
timestamp 1623621585
transform 1 0 11684 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_127
timestamp 1623621585
transform 1 0 12788 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_139
timestamp 1623621585
transform 1 0 13892 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_151
timestamp 1623621585
transform 1 0 14996 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_163
timestamp 1623621585
transform 1 0 16100 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1623621585
transform 1 0 16836 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_172
timestamp 1623621585
transform 1 0 16928 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_184
timestamp 1623621585
transform 1 0 18032 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_196
timestamp 1623621585
transform 1 0 19136 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_208
timestamp 1623621585
transform 1 0 20240 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1623621585
transform 1 0 22080 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_220
timestamp 1623621585
transform 1 0 21344 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_229
timestamp 1623621585
transform 1 0 22172 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_241
timestamp 1623621585
transform 1 0 23276 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1623621585
transform 1 0 24380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_265
timestamp 1623621585
transform 1 0 25484 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0557_
timestamp 1623621585
transform 1 0 26220 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1623621585
transform 1 0 27324 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_281
timestamp 1623621585
transform 1 0 26956 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_286
timestamp 1623621585
transform 1 0 27416 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_298
timestamp 1623621585
transform 1 0 28520 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_310
timestamp 1623621585
transform 1 0 29624 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_322
timestamp 1623621585
transform 1 0 30728 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1623621585
transform 1 0 32568 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_334
timestamp 1623621585
transform 1 0 31832 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_343
timestamp 1623621585
transform 1 0 32660 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input188
timestamp 1623621585
transform 1 0 35236 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_355
timestamp 1623621585
transform 1 0 33764 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_367
timestamp 1623621585
transform 1 0 34868 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_374
timestamp 1623621585
transform 1 0 35512 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0426_
timestamp 1623621585
transform 1 0 36524 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input156
timestamp 1623621585
transform 1 0 35880 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_381
timestamp 1623621585
transform 1 0 36156 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_389
timestamp 1623621585
transform 1 0 36892 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1623621585
transform -1 0 38824 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1623621585
transform 1 0 37812 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_397
timestamp 1623621585
transform 1 0 37628 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_400
timestamp 1623621585
transform 1 0 37904 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_406
timestamp 1623621585
transform 1 0 38456 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1623621585
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input380
timestamp 1623621585
transform 1 0 1380 0 1 47328
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_83_13
timestamp 1623621585
transform 1 0 2300 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1623621585
transform 1 0 3772 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_25
timestamp 1623621585
transform 1 0 3404 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_30
timestamp 1623621585
transform 1 0 3864 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1623621585
transform 1 0 4968 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_54
timestamp 1623621585
transform 1 0 6072 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_62
timestamp 1623621585
transform 1 0 6808 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0469_
timestamp 1623621585
transform 1 0 7084 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0589_
timestamp 1623621585
transform 1 0 8188 0 1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_83_68
timestamp 1623621585
transform 1 0 7360 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_76
timestamp 1623621585
transform 1 0 8096 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_82
timestamp 1623621585
transform 1 0 8648 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1623621585
transform 1 0 9476 0 1 47328
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1623621585
transform 1 0 9016 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_87
timestamp 1623621585
transform 1 0 9108 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_96
timestamp 1623621585
transform 1 0 9936 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_108
timestamp 1623621585
transform 1 0 11040 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_120
timestamp 1623621585
transform 1 0 12144 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1623621585
transform 1 0 14260 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_132
timestamp 1623621585
transform 1 0 13248 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_140
timestamp 1623621585
transform 1 0 13984 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_144
timestamp 1623621585
transform 1 0 14352 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_156
timestamp 1623621585
transform 1 0 15456 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_168
timestamp 1623621585
transform 1 0 16560 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_180
timestamp 1623621585
transform 1 0 17664 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1623621585
transform 1 0 19504 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_192
timestamp 1623621585
transform 1 0 18768 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_201
timestamp 1623621585
transform 1 0 19596 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_213
timestamp 1623621585
transform 1 0 20700 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_225
timestamp 1623621585
transform 1 0 21804 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_237
timestamp 1623621585
transform 1 0 22908 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1623621585
transform 1 0 24012 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1623621585
transform 1 0 24748 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_258
timestamp 1623621585
transform 1 0 24840 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_270
timestamp 1623621585
transform 1 0 25944 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _0548_
timestamp 1623621585
transform 1 0 26312 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_282
timestamp 1623621585
transform 1 0 27048 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_294
timestamp 1623621585
transform 1 0 28152 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_306
timestamp 1623621585
transform 1 0 29256 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1623621585
transform 1 0 29992 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_315
timestamp 1623621585
transform 1 0 30084 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_327
timestamp 1623621585
transform 1 0 31188 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_339
timestamp 1623621585
transform 1 0 32292 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_351
timestamp 1623621585
transform 1 0 33396 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1623621585
transform 1 0 35236 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_363
timestamp 1623621585
transform 1 0 34500 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_83_372
timestamp 1623621585
transform 1 0 35328 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0571_
timestamp 1623621585
transform 1 0 36524 0 1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input189
timestamp 1623621585
transform 1 0 35880 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_381
timestamp 1623621585
transform 1 0 36156 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_392
timestamp 1623621585
transform 1 0 37168 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0555_
timestamp 1623621585
transform 1 0 37536 0 1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1623621585
transform -1 0 38824 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_403
timestamp 1623621585
transform 1 0 38180 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1623621585
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input381
timestamp 1623621585
transform 1 0 1748 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_3
timestamp 1623621585
transform 1 0 1380 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_11
timestamp 1623621585
transform 1 0 2116 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_23
timestamp 1623621585
transform 1 0 3220 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_35
timestamp 1623621585
transform 1 0 4324 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1623621585
transform 1 0 6348 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_47
timestamp 1623621585
transform 1 0 5428 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_55
timestamp 1623621585
transform 1 0 6164 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_58
timestamp 1623621585
transform 1 0 6440 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0607_
timestamp 1623621585
transform 1 0 8556 0 -1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_84_70
timestamp 1623621585
transform 1 0 7544 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_78
timestamp 1623621585
transform 1 0 8280 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_86
timestamp 1623621585
transform 1 0 9016 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_98
timestamp 1623621585
transform 1 0 10120 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1623621585
transform 1 0 11592 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_110
timestamp 1623621585
transform 1 0 11224 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_115
timestamp 1623621585
transform 1 0 11684 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_127
timestamp 1623621585
transform 1 0 12788 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_139
timestamp 1623621585
transform 1 0 13892 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_151
timestamp 1623621585
transform 1 0 14996 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_163
timestamp 1623621585
transform 1 0 16100 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1623621585
transform 1 0 16836 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_172
timestamp 1623621585
transform 1 0 16928 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_184
timestamp 1623621585
transform 1 0 18032 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_196
timestamp 1623621585
transform 1 0 19136 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_208
timestamp 1623621585
transform 1 0 20240 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1623621585
transform 1 0 22080 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_220
timestamp 1623621585
transform 1 0 21344 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_229
timestamp 1623621585
transform 1 0 22172 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_241
timestamp 1623621585
transform 1 0 23276 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_253
timestamp 1623621585
transform 1 0 24380 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_265
timestamp 1623621585
transform 1 0 25484 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1623621585
transform 1 0 27324 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_277
timestamp 1623621585
transform 1 0 26588 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_286
timestamp 1623621585
transform 1 0 27416 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_298
timestamp 1623621585
transform 1 0 28520 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_310
timestamp 1623621585
transform 1 0 29624 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_322
timestamp 1623621585
transform 1 0 30728 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1623621585
transform 1 0 32568 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_334
timestamp 1623621585
transform 1 0 31832 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_343
timestamp 1623621585
transform 1 0 32660 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input190
timestamp 1623621585
transform 1 0 35512 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_355
timestamp 1623621585
transform 1 0 33764 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_367
timestamp 1623621585
transform 1 0 34868 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_373
timestamp 1623621585
transform 1 0 35420 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0563_
timestamp 1623621585
transform 1 0 36800 0 -1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1623621585
transform 1 0 36156 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_377
timestamp 1623621585
transform 1 0 35788 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_384
timestamp 1623621585
transform 1 0 36432 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_395
timestamp 1623621585
transform 1 0 37444 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1623621585
transform -1 0 38824 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1623621585
transform 1 0 37812 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_400
timestamp 1623621585
transform 1 0 37904 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_406
timestamp 1623621585
transform 1 0 38456 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1623621585
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1623621585
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input382
timestamp 1623621585
transform 1 0 1748 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1623621585
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1623621585
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1623621585
transform 1 0 1380 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_11
timestamp 1623621585
transform 1 0 2116 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1623621585
transform 1 0 3772 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_27
timestamp 1623621585
transform 1 0 3588 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_30
timestamp 1623621585
transform 1 0 3864 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_23
timestamp 1623621585
transform 1 0 3220 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_35
timestamp 1623621585
transform 1 0 4324 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1623621585
transform 1 0 6348 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_42
timestamp 1623621585
transform 1 0 4968 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_54
timestamp 1623621585
transform 1 0 6072 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_47
timestamp 1623621585
transform 1 0 5428 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_55
timestamp 1623621585
transform 1 0 6164 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_58
timestamp 1623621585
transform 1 0 6440 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0642_
timestamp 1623621585
transform 1 0 7176 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1623621585
transform 1 0 7452 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_81
timestamp 1623621585
transform 1 0 8556 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_70
timestamp 1623621585
transform 1 0 7544 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_82
timestamp 1623621585
transform 1 0 8648 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1623621585
transform 1 0 9016 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_85
timestamp 1623621585
transform 1 0 8924 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_87
timestamp 1623621585
transform 1 0 9108 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_99
timestamp 1623621585
transform 1 0 10212 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_94
timestamp 1623621585
transform 1 0 9752 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1623621585
transform 1 0 11592 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_111
timestamp 1623621585
transform 1 0 11316 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_123
timestamp 1623621585
transform 1 0 12420 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_106
timestamp 1623621585
transform 1 0 10856 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_115
timestamp 1623621585
transform 1 0 11684 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1623621585
transform 1 0 14260 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_135
timestamp 1623621585
transform 1 0 13524 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_144
timestamp 1623621585
transform 1 0 14352 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_127
timestamp 1623621585
transform 1 0 12788 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_139
timestamp 1623621585
transform 1 0 13892 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_156
timestamp 1623621585
transform 1 0 15456 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_151
timestamp 1623621585
transform 1 0 14996 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_163
timestamp 1623621585
transform 1 0 16100 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1623621585
transform 1 0 16836 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_168
timestamp 1623621585
transform 1 0 16560 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_180
timestamp 1623621585
transform 1 0 17664 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_172
timestamp 1623621585
transform 1 0 16928 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_184
timestamp 1623621585
transform 1 0 18032 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1623621585
transform 1 0 19504 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_192
timestamp 1623621585
transform 1 0 18768 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_201
timestamp 1623621585
transform 1 0 19596 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_196
timestamp 1623621585
transform 1 0 19136 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_208
timestamp 1623621585
transform 1 0 20240 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1623621585
transform 1 0 22080 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_213
timestamp 1623621585
transform 1 0 20700 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_225
timestamp 1623621585
transform 1 0 21804 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_220
timestamp 1623621585
transform 1 0 21344 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_86_229
timestamp 1623621585
transform 1 0 22172 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22816 0 -1 49504
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_85_237
timestamp 1623621585
transform 1 0 22908 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_249
timestamp 1623621585
transform 1 0 24012 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_235
timestamp 1623621585
transform 1 0 22724 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1623621585
transform 1 0 24748 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_258
timestamp 1623621585
transform 1 0 24840 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_270
timestamp 1623621585
transform 1 0 25944 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_253
timestamp 1623621585
transform 1 0 24380 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_265
timestamp 1623621585
transform 1 0 25484 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1623621585
transform 1 0 27324 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_282
timestamp 1623621585
transform 1 0 27048 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_277
timestamp 1623621585
transform 1 0 26588 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_286
timestamp 1623621585
transform 1 0 27416 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_294
timestamp 1623621585
transform 1 0 28152 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_306
timestamp 1623621585
transform 1 0 29256 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_298
timestamp 1623621585
transform 1 0 28520 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_310
timestamp 1623621585
transform 1 0 29624 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1623621585
transform 1 0 29992 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_315
timestamp 1623621585
transform 1 0 30084 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_327
timestamp 1623621585
transform 1 0 31188 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_322
timestamp 1623621585
transform 1 0 30728 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1623621585
transform 1 0 32568 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_339
timestamp 1623621585
transform 1 0 32292 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_351
timestamp 1623621585
transform 1 0 33396 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_334
timestamp 1623621585
transform 1 0 31832 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_343
timestamp 1623621585
transform 1 0 32660 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 1623621585
transform 1 0 35604 0 -1 49504
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1623621585
transform 1 0 35236 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_363
timestamp 1623621585
transform 1 0 34500 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_85_372
timestamp 1623621585
transform 1 0 35328 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_86_355
timestamp 1623621585
transform 1 0 33764 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_367
timestamp 1623621585
transform 1 0 34868 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0518_
timestamp 1623621585
transform 1 0 36616 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0527_
timestamp 1623621585
transform 1 0 36616 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input157
timestamp 1623621585
transform 1 0 35972 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_85_378
timestamp 1623621585
transform 1 0 35880 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_382
timestamp 1623621585
transform 1 0 36248 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_394
timestamp 1623621585
transform 1 0 37352 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_382
timestamp 1623621585
transform 1 0 36248 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_394
timestamp 1623621585
transform 1 0 37352 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0480_
timestamp 1623621585
transform 1 0 37812 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1623621585
transform -1 0 38824 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1623621585
transform -1 0 38824 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1623621585
transform 1 0 37812 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_398
timestamp 1623621585
transform 1 0 37720 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_403
timestamp 1623621585
transform 1 0 38180 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_398
timestamp 1623621585
transform 1 0 37720 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_400
timestamp 1623621585
transform 1 0 37904 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_406
timestamp 1623621585
transform 1 0 38456 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1623621585
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input383
timestamp 1623621585
transform 1 0 1748 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_3
timestamp 1623621585
transform 1 0 1380 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_11
timestamp 1623621585
transform 1 0 2116 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1623621585
transform 1 0 3772 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_23
timestamp 1623621585
transform 1 0 3220 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1623621585
transform 1 0 3864 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1623621585
transform 1 0 4968 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_54
timestamp 1623621585
transform 1 0 6072 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_66
timestamp 1623621585
transform 1 0 7176 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_78
timestamp 1623621585
transform 1 0 8280 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1623621585
transform 1 0 9016 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_87
timestamp 1623621585
transform 1 0 9108 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_99
timestamp 1623621585
transform 1 0 10212 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_111
timestamp 1623621585
transform 1 0 11316 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_123
timestamp 1623621585
transform 1 0 12420 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1623621585
transform 1 0 14260 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_135
timestamp 1623621585
transform 1 0 13524 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_144
timestamp 1623621585
transform 1 0 14352 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_156
timestamp 1623621585
transform 1 0 15456 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_168
timestamp 1623621585
transform 1 0 16560 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_180
timestamp 1623621585
transform 1 0 17664 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1623621585
transform 1 0 19504 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_192
timestamp 1623621585
transform 1 0 18768 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_201
timestamp 1623621585
transform 1 0 19596 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_213
timestamp 1623621585
transform 1 0 20700 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_225
timestamp 1623621585
transform 1 0 21804 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_237
timestamp 1623621585
transform 1 0 22908 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_249
timestamp 1623621585
transform 1 0 24012 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1623621585
transform 1 0 24748 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_258
timestamp 1623621585
transform 1 0 24840 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_270
timestamp 1623621585
transform 1 0 25944 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0528_
timestamp 1623621585
transform 1 0 26496 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_284
timestamp 1623621585
transform 1 0 27232 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_296
timestamp 1623621585
transform 1 0 28336 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_308
timestamp 1623621585
transform 1 0 29440 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1623621585
transform 1 0 29992 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_315
timestamp 1623621585
transform 1 0 30084 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_327
timestamp 1623621585
transform 1 0 31188 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_339
timestamp 1623621585
transform 1 0 32292 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_351
timestamp 1623621585
transform 1 0 33396 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1623621585
transform 1 0 35236 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_363
timestamp 1623621585
transform 1 0 34500 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_87_372
timestamp 1623621585
transform 1 0 35328 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0510_
timestamp 1623621585
transform 1 0 36708 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1623621585
transform 1 0 36064 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_383
timestamp 1623621585
transform 1 0 36340 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_395
timestamp 1623621585
transform 1 0 37444 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1623621585
transform -1 0 38824 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1623621585
transform 1 0 37904 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_87_399
timestamp 1623621585
transform 1 0 37812 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_403
timestamp 1623621585
transform 1 0 38180 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1623621585
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1623621585
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1623621585
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_27
timestamp 1623621585
transform 1 0 3588 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_39
timestamp 1623621585
transform 1 0 4692 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1623621585
transform 1 0 6348 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_51
timestamp 1623621585
transform 1 0 5796 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_88_58
timestamp 1623621585
transform 1 0 6440 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0588_
timestamp 1623621585
transform 1 0 7268 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_88_66
timestamp 1623621585
transform 1 0 7176 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_70
timestamp 1623621585
transform 1 0 7544 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_82
timestamp 1623621585
transform 1 0 8648 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_94
timestamp 1623621585
transform 1 0 9752 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1623621585
transform 1 0 11592 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_106
timestamp 1623621585
transform 1 0 10856 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_115
timestamp 1623621585
transform 1 0 11684 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_127
timestamp 1623621585
transform 1 0 12788 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_139
timestamp 1623621585
transform 1 0 13892 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_151
timestamp 1623621585
transform 1 0 14996 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_163
timestamp 1623621585
transform 1 0 16100 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1623621585
transform 1 0 16836 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_172
timestamp 1623621585
transform 1 0 16928 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_184
timestamp 1623621585
transform 1 0 18032 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_196
timestamp 1623621585
transform 1 0 19136 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_208
timestamp 1623621585
transform 1 0 20240 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1623621585
transform 1 0 22080 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_220
timestamp 1623621585
transform 1 0 21344 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_229
timestamp 1623621585
transform 1 0 22172 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_241
timestamp 1623621585
transform 1 0 23276 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0937_
timestamp 1623621585
transform 1 0 25116 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1623621585
transform 1 0 24380 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_267
timestamp 1623621585
transform 1 0 25668 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1623621585
transform 1 0 27324 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_279
timestamp 1623621585
transform 1 0 26772 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_88_286
timestamp 1623621585
transform 1 0 27416 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_298
timestamp 1623621585
transform 1 0 28520 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_310
timestamp 1623621585
transform 1 0 29624 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_322
timestamp 1623621585
transform 1 0 30728 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1623621585
transform 1 0 32568 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_334
timestamp 1623621585
transform 1 0 31832 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_343
timestamp 1623621585
transform 1 0 32660 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_355
timestamp 1623621585
transform 1 0 33764 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_367
timestamp 1623621585
transform 1 0 34868 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0502_
timestamp 1623621585
transform 1 0 36708 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input191
timestamp 1623621585
transform 1 0 36064 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_88_379
timestamp 1623621585
transform 1 0 35972 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_383
timestamp 1623621585
transform 1 0 36340 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_395
timestamp 1623621585
transform 1 0 37444 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1623621585
transform -1 0 38824 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1623621585
transform 1 0 37812 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_400
timestamp 1623621585
transform 1 0 37904 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_406
timestamp 1623621585
transform 1 0 38456 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1623621585
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input384
timestamp 1623621585
transform 1 0 1748 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_3
timestamp 1623621585
transform 1 0 1380 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_11
timestamp 1623621585
transform 1 0 2116 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1623621585
transform 1 0 3772 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_23
timestamp 1623621585
transform 1 0 3220 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_30
timestamp 1623621585
transform 1 0 3864 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1623621585
transform 1 0 4968 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_54
timestamp 1623621585
transform 1 0 6072 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_66
timestamp 1623621585
transform 1 0 7176 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_78
timestamp 1623621585
transform 1 0 8280 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1623621585
transform 1 0 9016 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_87
timestamp 1623621585
transform 1 0 9108 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_99
timestamp 1623621585
transform 1 0 10212 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_111
timestamp 1623621585
transform 1 0 11316 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_123
timestamp 1623621585
transform 1 0 12420 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1623621585
transform 1 0 14260 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_135
timestamp 1623621585
transform 1 0 13524 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_144
timestamp 1623621585
transform 1 0 14352 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_156
timestamp 1623621585
transform 1 0 15456 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_168
timestamp 1623621585
transform 1 0 16560 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_180
timestamp 1623621585
transform 1 0 17664 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1623621585
transform 1 0 19504 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_192
timestamp 1623621585
transform 1 0 18768 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_89_201
timestamp 1623621585
transform 1 0 19596 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0929_
timestamp 1623621585
transform 1 0 20332 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_215
timestamp 1623621585
transform 1 0 20884 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_227
timestamp 1623621585
transform 1 0 21988 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1623621585
transform 1 0 23368 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0932_
timestamp 1623621585
transform 1 0 22356 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_237
timestamp 1623621585
transform 1 0 22908 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_241
timestamp 1623621585
transform 1 0 23276 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_248
timestamp 1623621585
transform 1 0 23920 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0924_
timestamp 1623621585
transform 1 0 25208 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1623621585
transform 1 0 24748 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_256
timestamp 1623621585
transform 1 0 24656 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_258
timestamp 1623621585
transform 1 0 24840 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_268
timestamp 1623621585
transform 1 0 25760 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0520_
timestamp 1623621585
transform 1 0 26496 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_89_284
timestamp 1623621585
transform 1 0 27232 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _0817_
timestamp 1623621585
transform 1 0 28244 0 1 50592
box -38 -48 958 592
use sky130_fd_sc_hd__decap_3  FILLER_89_292
timestamp 1623621585
transform 1 0 27968 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_305
timestamp 1623621585
transform 1 0 29164 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0947_
timestamp 1623621585
transform 1 0 30452 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1623621585
transform 1 0 29992 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_313
timestamp 1623621585
transform 1 0 29900 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_315
timestamp 1623621585
transform 1 0 30084 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_325
timestamp 1623621585
transform 1 0 31004 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0953_
timestamp 1623621585
transform 1 0 32660 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_89_337
timestamp 1623621585
transform 1 0 32108 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_349
timestamp 1623621585
transform 1 0 33212 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1623621585
transform 1 0 35236 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_361
timestamp 1623621585
transform 1 0 34316 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_369
timestamp 1623621585
transform 1 0 35052 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_372
timestamp 1623621585
transform 1 0 35328 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0482_
timestamp 1623621585
transform 1 0 36708 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_384
timestamp 1623621585
transform 1 0 36432 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_395
timestamp 1623621585
transform 1 0 37444 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1623621585
transform -1 0 38824 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1623621585
transform 1 0 37904 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_89_399
timestamp 1623621585
transform 1 0 37812 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_403
timestamp 1623621585
transform 1 0 38180 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1623621585
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1623621585
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1623621585
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_27
timestamp 1623621585
transform 1 0 3588 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_39
timestamp 1623621585
transform 1 0 4692 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1623621585
transform 1 0 6348 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_51
timestamp 1623621585
transform 1 0 5796 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_58
timestamp 1623621585
transform 1 0 6440 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_70
timestamp 1623621585
transform 1 0 7544 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_82
timestamp 1623621585
transform 1 0 8648 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_94
timestamp 1623621585
transform 1 0 9752 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1623621585
transform 1 0 11592 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_106
timestamp 1623621585
transform 1 0 10856 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_115
timestamp 1623621585
transform 1 0 11684 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_127
timestamp 1623621585
transform 1 0 12788 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_139
timestamp 1623621585
transform 1 0 13892 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_151
timestamp 1623621585
transform 1 0 14996 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_163
timestamp 1623621585
transform 1 0 16100 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1623621585
transform 1 0 16836 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_172
timestamp 1623621585
transform 1 0 16928 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_184
timestamp 1623621585
transform 1 0 18032 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0960_
timestamp 1623621585
transform 1 0 19412 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_90_196
timestamp 1623621585
transform 1 0 19136 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_205
timestamp 1623621585
transform 1 0 19964 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1623621585
transform 1 0 22080 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_217
timestamp 1623621585
transform 1 0 21068 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_225
timestamp 1623621585
transform 1 0 21804 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_229
timestamp 1623621585
transform 1 0 22172 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0933_
timestamp 1623621585
transform 1 0 22908 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_243
timestamp 1623621585
transform 1 0 23460 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0936_
timestamp 1623621585
transform 1 0 24564 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_261
timestamp 1623621585
transform 1 0 25116 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0511_
timestamp 1623621585
transform 1 0 26220 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0942_
timestamp 1623621585
transform 1 0 27784 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1623621585
transform 1 0 27324 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_281
timestamp 1623621585
transform 1 0 26956 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_286
timestamp 1623621585
transform 1 0 27416 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0944_
timestamp 1623621585
transform 1 0 28704 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0946_
timestamp 1623621585
transform 1 0 29624 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_296
timestamp 1623621585
transform 1 0 28336 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_306
timestamp 1623621585
transform 1 0 29256 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_316
timestamp 1623621585
transform 1 0 30176 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_328
timestamp 1623621585
transform 1 0 31280 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1623621585
transform 1 0 32568 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_340
timestamp 1623621585
transform 1 0 32384 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_90_343
timestamp 1623621585
transform 1 0 32660 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0957_
timestamp 1623621585
transform 1 0 34500 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_90_355
timestamp 1623621585
transform 1 0 33764 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_369
timestamp 1623621585
transform 1 0 35052 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input159
timestamp 1623621585
transform 1 0 37168 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input192
timestamp 1623621585
transform 1 0 36524 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_381
timestamp 1623621585
transform 1 0 36156 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_388
timestamp 1623621585
transform 1 0 36800 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_395
timestamp 1623621585
transform 1 0 37444 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1623621585
transform -1 0 38824 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1623621585
transform 1 0 37812 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_90_400
timestamp 1623621585
transform 1 0 37904 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_406
timestamp 1623621585
transform 1 0 38456 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1623621585
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input386
timestamp 1623621585
transform 1 0 1748 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_3
timestamp 1623621585
transform 1 0 1380 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_11
timestamp 1623621585
transform 1 0 2116 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1623621585
transform 1 0 3772 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_23
timestamp 1623621585
transform 1 0 3220 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_91_30
timestamp 1623621585
transform 1 0 3864 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_42
timestamp 1623621585
transform 1 0 4968 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_54
timestamp 1623621585
transform 1 0 6072 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_66
timestamp 1623621585
transform 1 0 7176 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_78
timestamp 1623621585
transform 1 0 8280 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1623621585
transform 1 0 9016 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_87
timestamp 1623621585
transform 1 0 9108 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_99
timestamp 1623621585
transform 1 0 10212 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_111
timestamp 1623621585
transform 1 0 11316 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_123
timestamp 1623621585
transform 1 0 12420 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1623621585
transform 1 0 14260 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_135
timestamp 1623621585
transform 1 0 13524 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_144
timestamp 1623621585
transform 1 0 14352 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_156
timestamp 1623621585
transform 1 0 15456 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_168
timestamp 1623621585
transform 1 0 16560 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_180
timestamp 1623621585
transform 1 0 17664 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1623621585
transform 1 0 19504 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_192
timestamp 1623621585
transform 1 0 18768 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_201
timestamp 1623621585
transform 1 0 19596 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_213
timestamp 1623621585
transform 1 0 20700 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_225
timestamp 1623621585
transform 1 0 21804 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_237
timestamp 1623621585
transform 1 0 22908 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_249
timestamp 1623621585
transform 1 0 24012 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1623621585
transform 1 0 24748 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_258
timestamp 1623621585
transform 1 0 24840 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_270
timestamp 1623621585
transform 1 0 25944 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0503_
timestamp 1623621585
transform 1 0 26496 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_284
timestamp 1623621585
transform 1 0 27232 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_296
timestamp 1623621585
transform 1 0 28336 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_308
timestamp 1623621585
transform 1 0 29440 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1623621585
transform 1 0 29992 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_315
timestamp 1623621585
transform 1 0 30084 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_327
timestamp 1623621585
transform 1 0 31188 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_339
timestamp 1623621585
transform 1 0 32292 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_351
timestamp 1623621585
transform 1 0 33396 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1623621585
transform 1 0 35236 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_363
timestamp 1623621585
transform 1 0 34500 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_372
timestamp 1623621585
transform 1 0 35328 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_384
timestamp 1623621585
transform 1 0 36432 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0526_
timestamp 1623621585
transform 1 0 37536 0 1 51680
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1623621585
transform -1 0 38824 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_403
timestamp 1623621585
transform 1 0 38180 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1623621585
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1623621585
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input387
timestamp 1623621585
transform 1 0 1748 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_3
timestamp 1623621585
transform 1 0 1380 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_11
timestamp 1623621585
transform 1 0 2116 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1623621585
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1623621585
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1623621585
transform 1 0 3772 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_23
timestamp 1623621585
transform 1 0 3220 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_35
timestamp 1623621585
transform 1 0 4324 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_27
timestamp 1623621585
transform 1 0 3588 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_30
timestamp 1623621585
transform 1 0 3864 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1623621585
transform 1 0 6348 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_47
timestamp 1623621585
transform 1 0 5428 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_55
timestamp 1623621585
transform 1 0 6164 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_58
timestamp 1623621585
transform 1 0 6440 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_42
timestamp 1623621585
transform 1 0 4968 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_54
timestamp 1623621585
transform 1 0 6072 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_70
timestamp 1623621585
transform 1 0 7544 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_82
timestamp 1623621585
transform 1 0 8648 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_66
timestamp 1623621585
transform 1 0 7176 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_78
timestamp 1623621585
transform 1 0 8280 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1623621585
transform 1 0 9016 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_94
timestamp 1623621585
transform 1 0 9752 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_87
timestamp 1623621585
transform 1 0 9108 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_99
timestamp 1623621585
transform 1 0 10212 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1623621585
transform 1 0 11592 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_106
timestamp 1623621585
transform 1 0 10856 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_115
timestamp 1623621585
transform 1 0 11684 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_111
timestamp 1623621585
transform 1 0 11316 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_123
timestamp 1623621585
transform 1 0 12420 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1623621585
transform 1 0 14260 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_127
timestamp 1623621585
transform 1 0 12788 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_139
timestamp 1623621585
transform 1 0 13892 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_135
timestamp 1623621585
transform 1 0 13524 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_144
timestamp 1623621585
transform 1 0 14352 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_151
timestamp 1623621585
transform 1 0 14996 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_163
timestamp 1623621585
transform 1 0 16100 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_156
timestamp 1623621585
transform 1 0 15456 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1623621585
transform 1 0 16836 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_172
timestamp 1623621585
transform 1 0 16928 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_184
timestamp 1623621585
transform 1 0 18032 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_168
timestamp 1623621585
transform 1 0 16560 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_180
timestamp 1623621585
transform 1 0 17664 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1623621585
transform 1 0 19504 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_196
timestamp 1623621585
transform 1 0 19136 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_208
timestamp 1623621585
transform 1 0 20240 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_192
timestamp 1623621585
transform 1 0 18768 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_201
timestamp 1623621585
transform 1 0 19596 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1623621585
transform 1 0 22080 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_220
timestamp 1623621585
transform 1 0 21344 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_229
timestamp 1623621585
transform 1 0 22172 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_213
timestamp 1623621585
transform 1 0 20700 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_225
timestamp 1623621585
transform 1 0 21804 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_241
timestamp 1623621585
transform 1 0 23276 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_237
timestamp 1623621585
transform 1 0 22908 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_249
timestamp 1623621585
transform 1 0 24012 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1623621585
transform 1 0 24748 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_253
timestamp 1623621585
transform 1 0 24380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_265
timestamp 1623621585
transform 1 0 25484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_258
timestamp 1623621585
transform 1 0 24840 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_270
timestamp 1623621585
transform 1 0 25944 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0493_
timestamp 1623621585
transform 1 0 26496 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1623621585
transform 1 0 27324 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_277
timestamp 1623621585
transform 1 0 26588 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_286
timestamp 1623621585
transform 1 0 27416 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_284
timestamp 1623621585
transform 1 0 27232 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_298
timestamp 1623621585
transform 1 0 28520 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_310
timestamp 1623621585
transform 1 0 29624 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_296
timestamp 1623621585
transform 1 0 28336 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_308
timestamp 1623621585
transform 1 0 29440 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1623621585
transform 1 0 29992 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_322
timestamp 1623621585
transform 1 0 30728 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_315
timestamp 1623621585
transform 1 0 30084 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_327
timestamp 1623621585
transform 1 0 31188 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1623621585
transform 1 0 32568 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_334
timestamp 1623621585
transform 1 0 31832 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_343
timestamp 1623621585
transform 1 0 32660 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_339
timestamp 1623621585
transform 1 0 32292 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_351
timestamp 1623621585
transform 1 0 33396 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1623621585
transform 1 0 35236 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_355
timestamp 1623621585
transform 1 0 33764 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_367
timestamp 1623621585
transform 1 0 34868 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_363
timestamp 1623621585
transform 1 0 34500 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_93_372
timestamp 1623621585
transform 1 0 35328 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0517_
timestamp 1623621585
transform 1 0 36524 0 1 52768
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1623621585
transform 1 0 37168 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1623621585
transform 1 0 36524 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input194
timestamp 1623621585
transform 1 0 35880 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_379
timestamp 1623621585
transform 1 0 35972 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_388
timestamp 1623621585
transform 1 0 36800 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_395
timestamp 1623621585
transform 1 0 37444 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_381
timestamp 1623621585
transform 1 0 36156 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_392
timestamp 1623621585
transform 1 0 37168 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0509_
timestamp 1623621585
transform 1 0 37536 0 1 52768
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1623621585
transform -1 0 38824 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1623621585
transform -1 0 38824 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1623621585
transform 1 0 37812 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_400
timestamp 1623621585
transform 1 0 37904 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_406
timestamp 1623621585
transform 1 0 38456 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_403
timestamp 1623621585
transform 1 0 38180 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1623621585
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input395
timestamp 1623621585
transform 1 0 1380 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_6
timestamp 1623621585
transform 1 0 1656 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_18
timestamp 1623621585
transform 1 0 2760 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_30
timestamp 1623621585
transform 1 0 3864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1623621585
transform 1 0 6348 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_42
timestamp 1623621585
transform 1 0 4968 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_54
timestamp 1623621585
transform 1 0 6072 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_58
timestamp 1623621585
transform 1 0 6440 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_70
timestamp 1623621585
transform 1 0 7544 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_82
timestamp 1623621585
transform 1 0 8648 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_94
timestamp 1623621585
transform 1 0 9752 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1623621585
transform 1 0 11592 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_106
timestamp 1623621585
transform 1 0 10856 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_115
timestamp 1623621585
transform 1 0 11684 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_127
timestamp 1623621585
transform 1 0 12788 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_139
timestamp 1623621585
transform 1 0 13892 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_151
timestamp 1623621585
transform 1 0 14996 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_163
timestamp 1623621585
transform 1 0 16100 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1623621585
transform 1 0 16836 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_172
timestamp 1623621585
transform 1 0 16928 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_184
timestamp 1623621585
transform 1 0 18032 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_196
timestamp 1623621585
transform 1 0 19136 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_208
timestamp 1623621585
transform 1 0 20240 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1623621585
transform 1 0 22080 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_220
timestamp 1623621585
transform 1 0 21344 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_229
timestamp 1623621585
transform 1 0 22172 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_241
timestamp 1623621585
transform 1 0 23276 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_253
timestamp 1623621585
transform 1 0 24380 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_265
timestamp 1623621585
transform 1 0 25484 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1623621585
transform 1 0 27324 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_277
timestamp 1623621585
transform 1 0 26588 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_286
timestamp 1623621585
transform 1 0 27416 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_298
timestamp 1623621585
transform 1 0 28520 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_310
timestamp 1623621585
transform 1 0 29624 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_322
timestamp 1623621585
transform 1 0 30728 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1623621585
transform 1 0 32568 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_334
timestamp 1623621585
transform 1 0 31832 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_343
timestamp 1623621585
transform 1 0 32660 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_355
timestamp 1623621585
transform 1 0 33764 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_367
timestamp 1623621585
transform 1 0 34868 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1623621585
transform 1 0 37168 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input162
timestamp 1623621585
transform 1 0 36524 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_94_379
timestamp 1623621585
transform 1 0 35972 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_388
timestamp 1623621585
transform 1 0 36800 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_395
timestamp 1623621585
transform 1 0 37444 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1623621585
transform -1 0 38824 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1623621585
transform 1 0 37812 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_400
timestamp 1623621585
transform 1 0 37904 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_406
timestamp 1623621585
transform 1 0 38456 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1623621585
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input406
timestamp 1623621585
transform 1 0 1380 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_6
timestamp 1623621585
transform 1 0 1656 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_18
timestamp 1623621585
transform 1 0 2760 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1623621585
transform 1 0 3772 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_26
timestamp 1623621585
transform 1 0 3496 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_30
timestamp 1623621585
transform 1 0 3864 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_42
timestamp 1623621585
transform 1 0 4968 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_54
timestamp 1623621585
transform 1 0 6072 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_66
timestamp 1623621585
transform 1 0 7176 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_78
timestamp 1623621585
transform 1 0 8280 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1623621585
transform 1 0 9016 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_87
timestamp 1623621585
transform 1 0 9108 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_99
timestamp 1623621585
transform 1 0 10212 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_111
timestamp 1623621585
transform 1 0 11316 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_123
timestamp 1623621585
transform 1 0 12420 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1623621585
transform 1 0 14260 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_135
timestamp 1623621585
transform 1 0 13524 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_144
timestamp 1623621585
transform 1 0 14352 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_156
timestamp 1623621585
transform 1 0 15456 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_168
timestamp 1623621585
transform 1 0 16560 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_180
timestamp 1623621585
transform 1 0 17664 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1623621585
transform 1 0 19504 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_192
timestamp 1623621585
transform 1 0 18768 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_201
timestamp 1623621585
transform 1 0 19596 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_213
timestamp 1623621585
transform 1 0 20700 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_225
timestamp 1623621585
transform 1 0 21804 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_237
timestamp 1623621585
transform 1 0 22908 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_249
timestamp 1623621585
transform 1 0 24012 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1623621585
transform 1 0 24748 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_258
timestamp 1623621585
transform 1 0 24840 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_270
timestamp 1623621585
transform 1 0 25944 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_282
timestamp 1623621585
transform 1 0 27048 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_294
timestamp 1623621585
transform 1 0 28152 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_306
timestamp 1623621585
transform 1 0 29256 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1623621585
transform 1 0 29992 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_315
timestamp 1623621585
transform 1 0 30084 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_327
timestamp 1623621585
transform 1 0 31188 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_339
timestamp 1623621585
transform 1 0 32292 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_351
timestamp 1623621585
transform 1 0 33396 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1623621585
transform 1 0 35236 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_363
timestamp 1623621585
transform 1 0 34500 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_95_372
timestamp 1623621585
transform 1 0 35328 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1623621585
transform 1 0 36892 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1623621585
transform 1 0 36248 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_380
timestamp 1623621585
transform 1 0 36064 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_385
timestamp 1623621585
transform 1 0 36524 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_392
timestamp 1623621585
transform 1 0 37168 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0501_
timestamp 1623621585
transform 1 0 37536 0 1 53856
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1623621585
transform -1 0 38824 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_403
timestamp 1623621585
transform 1 0 38180 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1623621585
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1623621585
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1623621585
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_27
timestamp 1623621585
transform 1 0 3588 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_39
timestamp 1623621585
transform 1 0 4692 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1623621585
transform 1 0 6348 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_51
timestamp 1623621585
transform 1 0 5796 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_58
timestamp 1623621585
transform 1 0 6440 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_70
timestamp 1623621585
transform 1 0 7544 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_82
timestamp 1623621585
transform 1 0 8648 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_94
timestamp 1623621585
transform 1 0 9752 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1623621585
transform 1 0 11592 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_106
timestamp 1623621585
transform 1 0 10856 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_115
timestamp 1623621585
transform 1 0 11684 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_127
timestamp 1623621585
transform 1 0 12788 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_139
timestamp 1623621585
transform 1 0 13892 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_151
timestamp 1623621585
transform 1 0 14996 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_163
timestamp 1623621585
transform 1 0 16100 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1623621585
transform 1 0 16836 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_172
timestamp 1623621585
transform 1 0 16928 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_184
timestamp 1623621585
transform 1 0 18032 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_196
timestamp 1623621585
transform 1 0 19136 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_208
timestamp 1623621585
transform 1 0 20240 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1623621585
transform 1 0 22080 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_220
timestamp 1623621585
transform 1 0 21344 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_229
timestamp 1623621585
transform 1 0 22172 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_241
timestamp 1623621585
transform 1 0 23276 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_253
timestamp 1623621585
transform 1 0 24380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_265
timestamp 1623621585
transform 1 0 25484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1623621585
transform 1 0 27324 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_277
timestamp 1623621585
transform 1 0 26588 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_286
timestamp 1623621585
transform 1 0 27416 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_298
timestamp 1623621585
transform 1 0 28520 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_310
timestamp 1623621585
transform 1 0 29624 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_322
timestamp 1623621585
transform 1 0 30728 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1623621585
transform 1 0 32568 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_334
timestamp 1623621585
transform 1 0 31832 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_343
timestamp 1623621585
transform 1 0 32660 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input195
timestamp 1623621585
transform 1 0 35512 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_355
timestamp 1623621585
transform 1 0 33764 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_367
timestamp 1623621585
transform 1 0 34868 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_373
timestamp 1623621585
transform 1 0 35420 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _0460_
timestamp 1623621585
transform 1 0 36156 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_96_377
timestamp 1623621585
transform 1 0 35788 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_389
timestamp 1623621585
transform 1 0 36892 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1623621585
transform -1 0 38824 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1623621585
transform 1 0 37812 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_397
timestamp 1623621585
transform 1 0 37628 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_400
timestamp 1623621585
transform 1 0 37904 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_406
timestamp 1623621585
transform 1 0 38456 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1623621585
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input417
timestamp 1623621585
transform 1 0 1380 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_6
timestamp 1623621585
transform 1 0 1656 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_18
timestamp 1623621585
transform 1 0 2760 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1623621585
transform 1 0 3772 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_97_26
timestamp 1623621585
transform 1 0 3496 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_30
timestamp 1623621585
transform 1 0 3864 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_42
timestamp 1623621585
transform 1 0 4968 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_54
timestamp 1623621585
transform 1 0 6072 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_66
timestamp 1623621585
transform 1 0 7176 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_78
timestamp 1623621585
transform 1 0 8280 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1623621585
transform 1 0 9016 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_87
timestamp 1623621585
transform 1 0 9108 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_99
timestamp 1623621585
transform 1 0 10212 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_111
timestamp 1623621585
transform 1 0 11316 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_123
timestamp 1623621585
transform 1 0 12420 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1623621585
transform 1 0 14260 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_135
timestamp 1623621585
transform 1 0 13524 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_144
timestamp 1623621585
transform 1 0 14352 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_156
timestamp 1623621585
transform 1 0 15456 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_168
timestamp 1623621585
transform 1 0 16560 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_180
timestamp 1623621585
transform 1 0 17664 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1623621585
transform 1 0 19504 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_192
timestamp 1623621585
transform 1 0 18768 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_201
timestamp 1623621585
transform 1 0 19596 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_213
timestamp 1623621585
transform 1 0 20700 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_225
timestamp 1623621585
transform 1 0 21804 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_237
timestamp 1623621585
transform 1 0 22908 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_249
timestamp 1623621585
transform 1 0 24012 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1623621585
transform 1 0 24748 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_258
timestamp 1623621585
transform 1 0 24840 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_270
timestamp 1623621585
transform 1 0 25944 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_282
timestamp 1623621585
transform 1 0 27048 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0434_
timestamp 1623621585
transform 1 0 28980 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_294
timestamp 1623621585
transform 1 0 28152 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_302
timestamp 1623621585
transform 1 0 28888 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_307
timestamp 1623621585
transform 1 0 29348 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1623621585
transform 1 0 29992 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_313
timestamp 1623621585
transform 1 0 29900 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_315
timestamp 1623621585
transform 1 0 30084 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_327
timestamp 1623621585
transform 1 0 31188 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_339
timestamp 1623621585
transform 1 0 32292 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_351
timestamp 1623621585
transform 1 0 33396 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1623621585
transform 1 0 35236 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input203
timestamp 1623621585
transform 1 0 34592 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_97_363
timestamp 1623621585
transform 1 0 34500 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_367
timestamp 1623621585
transform 1 0 34868 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_372
timestamp 1623621585
transform 1 0 35328 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0451_
timestamp 1623621585
transform 1 0 36156 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_380
timestamp 1623621585
transform 1 0 36064 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_389
timestamp 1623621585
transform 1 0 36892 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_395
timestamp 1623621585
transform 1 0 37444 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _0481_
timestamp 1623621585
transform 1 0 37536 0 1 54944
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1623621585
transform -1 0 38824 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_403
timestamp 1623621585
transform 1 0 38180 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1623621585
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input420
timestamp 1623621585
transform 1 0 1380 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_6
timestamp 1623621585
transform 1 0 1656 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_18
timestamp 1623621585
transform 1 0 2760 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_30
timestamp 1623621585
transform 1 0 3864 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1623621585
transform 1 0 6348 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_42
timestamp 1623621585
transform 1 0 4968 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_54
timestamp 1623621585
transform 1 0 6072 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_58
timestamp 1623621585
transform 1 0 6440 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_70
timestamp 1623621585
transform 1 0 7544 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_82
timestamp 1623621585
transform 1 0 8648 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_94
timestamp 1623621585
transform 1 0 9752 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1623621585
transform 1 0 11592 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_106
timestamp 1623621585
transform 1 0 10856 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_115
timestamp 1623621585
transform 1 0 11684 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_127
timestamp 1623621585
transform 1 0 12788 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_139
timestamp 1623621585
transform 1 0 13892 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_151
timestamp 1623621585
transform 1 0 14996 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_163
timestamp 1623621585
transform 1 0 16100 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1623621585
transform 1 0 16836 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_172
timestamp 1623621585
transform 1 0 16928 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_184
timestamp 1623621585
transform 1 0 18032 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_196
timestamp 1623621585
transform 1 0 19136 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_208
timestamp 1623621585
transform 1 0 20240 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1623621585
transform 1 0 22080 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_220
timestamp 1623621585
transform 1 0 21344 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_229
timestamp 1623621585
transform 1 0 22172 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_241
timestamp 1623621585
transform 1 0 23276 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_253
timestamp 1623621585
transform 1 0 24380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_265
timestamp 1623621585
transform 1 0 25484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1623621585
transform 1 0 27324 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_277
timestamp 1623621585
transform 1 0 26588 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_286
timestamp 1623621585
transform 1 0 27416 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_298
timestamp 1623621585
transform 1 0 28520 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_310
timestamp 1623621585
transform 1 0 29624 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_322
timestamp 1623621585
transform 1 0 30728 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1623621585
transform 1 0 32568 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_334
timestamp 1623621585
transform 1 0 31832 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_343
timestamp 1623621585
transform 1 0 32660 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0425_
timestamp 1623621585
transform 1 0 35420 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input214
timestamp 1623621585
transform 1 0 34776 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_355
timestamp 1623621585
transform 1 0 33764 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_363
timestamp 1623621585
transform 1 0 34500 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_369
timestamp 1623621585
transform 1 0 35052 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0429_
timestamp 1623621585
transform 1 0 36156 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_377
timestamp 1623621585
transform 1 0 35788 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_389
timestamp 1623621585
transform 1 0 36892 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1623621585
transform -1 0 38824 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1623621585
transform 1 0 37812 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_397
timestamp 1623621585
transform 1 0 37628 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_400
timestamp 1623621585
transform 1 0 37904 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_406
timestamp 1623621585
transform 1 0 38456 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1623621585
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1623621585
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input421
timestamp 1623621585
transform 1 0 1380 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1623621585
transform 1 0 1380 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1623621585
transform 1 0 2484 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_6
timestamp 1623621585
transform 1 0 1656 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_18
timestamp 1623621585
transform 1 0 2760 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1623621585
transform 1 0 3772 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_27
timestamp 1623621585
transform 1 0 3588 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_30
timestamp 1623621585
transform 1 0 3864 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_30
timestamp 1623621585
transform 1 0 3864 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1623621585
transform 1 0 6348 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_42
timestamp 1623621585
transform 1 0 4968 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_54
timestamp 1623621585
transform 1 0 6072 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_42
timestamp 1623621585
transform 1 0 4968 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_54
timestamp 1623621585
transform 1 0 6072 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_58
timestamp 1623621585
transform 1 0 6440 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_66
timestamp 1623621585
transform 1 0 7176 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_78
timestamp 1623621585
transform 1 0 8280 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_70
timestamp 1623621585
transform 1 0 7544 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_82
timestamp 1623621585
transform 1 0 8648 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1623621585
transform 1 0 9016 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_87
timestamp 1623621585
transform 1 0 9108 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_99
timestamp 1623621585
transform 1 0 10212 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_94
timestamp 1623621585
transform 1 0 9752 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1623621585
transform 1 0 11592 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_111
timestamp 1623621585
transform 1 0 11316 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_123
timestamp 1623621585
transform 1 0 12420 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_106
timestamp 1623621585
transform 1 0 10856 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_115
timestamp 1623621585
transform 1 0 11684 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1623621585
transform 1 0 14260 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_135
timestamp 1623621585
transform 1 0 13524 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_144
timestamp 1623621585
transform 1 0 14352 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_127
timestamp 1623621585
transform 1 0 12788 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_139
timestamp 1623621585
transform 1 0 13892 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_156
timestamp 1623621585
transform 1 0 15456 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_151
timestamp 1623621585
transform 1 0 14996 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_163
timestamp 1623621585
transform 1 0 16100 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1623621585
transform 1 0 16836 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_168
timestamp 1623621585
transform 1 0 16560 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_180
timestamp 1623621585
transform 1 0 17664 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_172
timestamp 1623621585
transform 1 0 16928 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_184
timestamp 1623621585
transform 1 0 18032 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1623621585
transform 1 0 19504 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_192
timestamp 1623621585
transform 1 0 18768 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_201
timestamp 1623621585
transform 1 0 19596 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_196
timestamp 1623621585
transform 1 0 19136 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_208
timestamp 1623621585
transform 1 0 20240 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1623621585
transform 1 0 22080 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_213
timestamp 1623621585
transform 1 0 20700 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_225
timestamp 1623621585
transform 1 0 21804 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_220
timestamp 1623621585
transform 1 0 21344 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_229
timestamp 1623621585
transform 1 0 22172 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_237
timestamp 1623621585
transform 1 0 22908 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_249
timestamp 1623621585
transform 1 0 24012 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_241
timestamp 1623621585
transform 1 0 23276 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1623621585
transform 1 0 24748 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_258
timestamp 1623621585
transform 1 0 24840 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_270
timestamp 1623621585
transform 1 0 25944 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_253
timestamp 1623621585
transform 1 0 24380 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_265
timestamp 1623621585
transform 1 0 25484 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0453_
timestamp 1623621585
transform 1 0 26312 0 -1 57120
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0461_
timestamp 1623621585
transform 1 0 26680 0 1 56032
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1623621585
transform 1 0 27324 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_285
timestamp 1623621585
transform 1 0 27324 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_273
timestamp 1623621585
transform 1 0 26220 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_281
timestamp 1623621585
transform 1 0 26956 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_286
timestamp 1623621585
transform 1 0 27416 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_297
timestamp 1623621585
transform 1 0 28428 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_309
timestamp 1623621585
transform 1 0 29532 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_298
timestamp 1623621585
transform 1 0 28520 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_310
timestamp 1623621585
transform 1 0 29624 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1623621585
transform 1 0 29992 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_313
timestamp 1623621585
transform 1 0 29900 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_315
timestamp 1623621585
transform 1 0 30084 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_327
timestamp 1623621585
transform 1 0 31188 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_322
timestamp 1623621585
transform 1 0 30728 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1623621585
transform 1 0 32568 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_339
timestamp 1623621585
transform 1 0 32292 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_351
timestamp 1623621585
transform 1 0 33396 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_334
timestamp 1623621585
transform 1 0 31832 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_343
timestamp 1623621585
transform 1 0 32660 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1623621585
transform 1 0 35236 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_363
timestamp 1623621585
transform 1 0 34500 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_99_372
timestamp 1623621585
transform 1 0 35328 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_355
timestamp 1623621585
transform 1 0 33764 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_367
timestamp 1623621585
transform 1 0 34868 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0427_
timestamp 1623621585
transform 1 0 37260 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0443_
timestamp 1623621585
transform 1 0 36156 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1623621585
transform 1 0 37076 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1623621585
transform 1 0 36340 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_380
timestamp 1623621585
transform 1 0 36064 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_389
timestamp 1623621585
transform 1 0 36892 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_379
timestamp 1623621585
transform 1 0 35972 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_387
timestamp 1623621585
transform 1 0 36708 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_395
timestamp 1623621585
transform 1 0 37444 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1623621585
transform -1 0 38824 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1623621585
transform -1 0 38824 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1623621585
transform 1 0 37812 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_397
timestamp 1623621585
transform 1 0 37628 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_405
timestamp 1623621585
transform 1 0 38364 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_100_400
timestamp 1623621585
transform 1 0 37904 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_406
timestamp 1623621585
transform 1 0 38456 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1623621585
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input422
timestamp 1623621585
transform 1 0 1380 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_6
timestamp 1623621585
transform 1 0 1656 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_18
timestamp 1623621585
transform 1 0 2760 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1623621585
transform 1 0 3772 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_26
timestamp 1623621585
transform 1 0 3496 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_30
timestamp 1623621585
transform 1 0 3864 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_42
timestamp 1623621585
transform 1 0 4968 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_54
timestamp 1623621585
transform 1 0 6072 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_66
timestamp 1623621585
transform 1 0 7176 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_78
timestamp 1623621585
transform 1 0 8280 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1623621585
transform 1 0 9016 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_87
timestamp 1623621585
transform 1 0 9108 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_99
timestamp 1623621585
transform 1 0 10212 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_111
timestamp 1623621585
transform 1 0 11316 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_123
timestamp 1623621585
transform 1 0 12420 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1623621585
transform 1 0 14260 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_135
timestamp 1623621585
transform 1 0 13524 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_144
timestamp 1623621585
transform 1 0 14352 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_156
timestamp 1623621585
transform 1 0 15456 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_168
timestamp 1623621585
transform 1 0 16560 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_180
timestamp 1623621585
transform 1 0 17664 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1623621585
transform 1 0 19504 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_192
timestamp 1623621585
transform 1 0 18768 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_201
timestamp 1623621585
transform 1 0 19596 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_213
timestamp 1623621585
transform 1 0 20700 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_225
timestamp 1623621585
transform 1 0 21804 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_237
timestamp 1623621585
transform 1 0 22908 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_249
timestamp 1623621585
transform 1 0 24012 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1623621585
transform 1 0 24748 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_258
timestamp 1623621585
transform 1 0 24840 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_270
timestamp 1623621585
transform 1 0 25944 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0444_
timestamp 1623621585
transform 1 0 26588 0 1 57120
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_101_276
timestamp 1623621585
transform 1 0 26496 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_284
timestamp 1623621585
transform 1 0 27232 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0433_
timestamp 1623621585
transform 1 0 28888 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_296
timestamp 1623621585
transform 1 0 28336 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_306
timestamp 1623621585
transform 1 0 29256 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1623621585
transform 1 0 29992 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_315
timestamp 1623621585
transform 1 0 30084 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_327
timestamp 1623621585
transform 1 0 31188 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_339
timestamp 1623621585
transform 1 0 32292 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_351
timestamp 1623621585
transform 1 0 33396 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1623621585
transform 1 0 35236 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_363
timestamp 1623621585
transform 1 0 34500 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_372
timestamp 1623621585
transform 1 0 35328 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input225
timestamp 1623621585
transform 1 0 36892 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_384
timestamp 1623621585
transform 1 0 36432 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_388
timestamp 1623621585
transform 1 0 36800 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_392
timestamp 1623621585
transform 1 0 37168 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0459_
timestamp 1623621585
transform 1 0 37536 0 1 57120
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1623621585
transform -1 0 38824 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_403
timestamp 1623621585
transform 1 0 38180 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1623621585
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1623621585
transform 1 0 1380 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_15
timestamp 1623621585
transform 1 0 2484 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_27
timestamp 1623621585
transform 1 0 3588 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_39
timestamp 1623621585
transform 1 0 4692 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1623621585
transform 1 0 6348 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_51
timestamp 1623621585
transform 1 0 5796 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_102_58
timestamp 1623621585
transform 1 0 6440 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_70
timestamp 1623621585
transform 1 0 7544 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_82
timestamp 1623621585
transform 1 0 8648 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_94
timestamp 1623621585
transform 1 0 9752 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0457_
timestamp 1623621585
transform 1 0 12052 0 -1 58208
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1623621585
transform 1 0 11592 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_106
timestamp 1623621585
transform 1 0 10856 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_102_115
timestamp 1623621585
transform 1 0 11684 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_124
timestamp 1623621585
transform 1 0 12512 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_136
timestamp 1623621585
transform 1 0 13616 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_148
timestamp 1623621585
transform 1 0 14720 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_160
timestamp 1623621585
transform 1 0 15824 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1623621585
transform 1 0 16836 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_102_168
timestamp 1623621585
transform 1 0 16560 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_172
timestamp 1623621585
transform 1 0 16928 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_184
timestamp 1623621585
transform 1 0 18032 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_196
timestamp 1623621585
transform 1 0 19136 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_208
timestamp 1623621585
transform 1 0 20240 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1623621585
transform 1 0 22080 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_220
timestamp 1623621585
transform 1 0 21344 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_229
timestamp 1623621585
transform 1 0 22172 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_241
timestamp 1623621585
transform 1 0 23276 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_253
timestamp 1623621585
transform 1 0 24380 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_265
timestamp 1623621585
transform 1 0 25484 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1623621585
transform 1 0 27324 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_277
timestamp 1623621585
transform 1 0 26588 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_286
timestamp 1623621585
transform 1 0 27416 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_298
timestamp 1623621585
transform 1 0 28520 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_310
timestamp 1623621585
transform 1 0 29624 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_322
timestamp 1623621585
transform 1 0 30728 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1623621585
transform 1 0 32568 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_334
timestamp 1623621585
transform 1 0 31832 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_343
timestamp 1623621585
transform 1 0 32660 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_355
timestamp 1623621585
transform 1 0 33764 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_367
timestamp 1623621585
transform 1 0 34868 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1623621585
transform 1 0 37076 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1623621585
transform 1 0 36340 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_379
timestamp 1623621585
transform 1 0 35972 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_387
timestamp 1623621585
transform 1 0 36708 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_395
timestamp 1623621585
transform 1 0 37444 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1623621585
transform -1 0 38824 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1623621585
transform 1 0 37812 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_400
timestamp 1623621585
transform 1 0 37904 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_406
timestamp 1623621585
transform 1 0 38456 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1623621585
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input423
timestamp 1623621585
transform 1 0 1380 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_6
timestamp 1623621585
transform 1 0 1656 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_18
timestamp 1623621585
transform 1 0 2760 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1623621585
transform 1 0 3772 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_103_26
timestamp 1623621585
transform 1 0 3496 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_30
timestamp 1623621585
transform 1 0 3864 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_42
timestamp 1623621585
transform 1 0 4968 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_54
timestamp 1623621585
transform 1 0 6072 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_66
timestamp 1623621585
transform 1 0 7176 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_78
timestamp 1623621585
transform 1 0 8280 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1623621585
transform 1 0 9016 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_87
timestamp 1623621585
transform 1 0 9108 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_99
timestamp 1623621585
transform 1 0 10212 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0422_
timestamp 1623621585
transform 1 0 11960 0 1 58208
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_103_111
timestamp 1623621585
transform 1 0 11316 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_117
timestamp 1623621585
transform 1 0 11868 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_123
timestamp 1623621585
transform 1 0 12420 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0440_
timestamp 1623621585
transform 1 0 12788 0 1 58208
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1623621585
transform 1 0 14260 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_132
timestamp 1623621585
transform 1 0 13248 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_140
timestamp 1623621585
transform 1 0 13984 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_144
timestamp 1623621585
transform 1 0 14352 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_156
timestamp 1623621585
transform 1 0 15456 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_168
timestamp 1623621585
transform 1 0 16560 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_180
timestamp 1623621585
transform 1 0 17664 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1623621585
transform 1 0 19504 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_192
timestamp 1623621585
transform 1 0 18768 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_201
timestamp 1623621585
transform 1 0 19596 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_213
timestamp 1623621585
transform 1 0 20700 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_225
timestamp 1623621585
transform 1 0 21804 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_237
timestamp 1623621585
transform 1 0 22908 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_249
timestamp 1623621585
transform 1 0 24012 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1623621585
transform 1 0 24748 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_258
timestamp 1623621585
transform 1 0 24840 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_270
timestamp 1623621585
transform 1 0 25944 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0435_
timestamp 1623621585
transform 1 0 26588 0 1 58208
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_103_276
timestamp 1623621585
transform 1 0 26496 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_284
timestamp 1623621585
transform 1 0 27232 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_296
timestamp 1623621585
transform 1 0 28336 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_308
timestamp 1623621585
transform 1 0 29440 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1623621585
transform 1 0 29992 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_315
timestamp 1623621585
transform 1 0 30084 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_327
timestamp 1623621585
transform 1 0 31188 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_339
timestamp 1623621585
transform 1 0 32292 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_351
timestamp 1623621585
transform 1 0 33396 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1623621585
transform 1 0 35236 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_103_363
timestamp 1623621585
transform 1 0 34500 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_372
timestamp 1623621585
transform 1 0 35328 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0450_
timestamp 1623621585
transform 1 0 36524 0 1 58208
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_103_384
timestamp 1623621585
transform 1 0 36432 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_392
timestamp 1623621585
transform 1 0 37168 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0442_
timestamp 1623621585
transform 1 0 37536 0 1 58208
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1623621585
transform -1 0 38824 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_403
timestamp 1623621585
transform 1 0 38180 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1623621585
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input424
timestamp 1623621585
transform 1 0 1380 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_6
timestamp 1623621585
transform 1 0 1656 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_18
timestamp 1623621585
transform 1 0 2760 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_30
timestamp 1623621585
transform 1 0 3864 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1623621585
transform 1 0 6348 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_42
timestamp 1623621585
transform 1 0 4968 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_54
timestamp 1623621585
transform 1 0 6072 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_58
timestamp 1623621585
transform 1 0 6440 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_70
timestamp 1623621585
transform 1 0 7544 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_82
timestamp 1623621585
transform 1 0 8648 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0421_
timestamp 1623621585
transform 1 0 10120 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_94
timestamp 1623621585
transform 1 0 9752 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_102
timestamp 1623621585
transform 1 0 10488 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _0448_
timestamp 1623621585
transform 1 0 12052 0 -1 59296
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1623621585
transform 1 0 11592 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_115
timestamp 1623621585
transform 1 0 11684 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_104_124
timestamp 1623621585
transform 1 0 12512 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_136
timestamp 1623621585
transform 1 0 13616 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_148
timestamp 1623621585
transform 1 0 14720 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_160
timestamp 1623621585
transform 1 0 15824 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1623621585
transform 1 0 16836 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_168
timestamp 1623621585
transform 1 0 16560 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_104_172
timestamp 1623621585
transform 1 0 16928 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_184
timestamp 1623621585
transform 1 0 18032 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_196
timestamp 1623621585
transform 1 0 19136 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_208
timestamp 1623621585
transform 1 0 20240 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1623621585
transform 1 0 22080 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_220
timestamp 1623621585
transform 1 0 21344 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_229
timestamp 1623621585
transform 1 0 22172 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_241
timestamp 1623621585
transform 1 0 23276 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_253
timestamp 1623621585
transform 1 0 24380 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_265
timestamp 1623621585
transform 1 0 25484 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1623621585
transform 1 0 27324 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_277
timestamp 1623621585
transform 1 0 26588 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_286
timestamp 1623621585
transform 1 0 27416 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_298
timestamp 1623621585
transform 1 0 28520 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_310
timestamp 1623621585
transform 1 0 29624 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_322
timestamp 1623621585
transform 1 0 30728 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1623621585
transform 1 0 32568 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_334
timestamp 1623621585
transform 1 0 31832 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_104_343
timestamp 1623621585
transform 1 0 32660 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_355
timestamp 1623621585
transform 1 0 33764 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_367
timestamp 1623621585
transform 1 0 34868 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input232
timestamp 1623621585
transform 1 0 37076 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input233
timestamp 1623621585
transform 1 0 36432 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_379
timestamp 1623621585
transform 1 0 35972 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_383
timestamp 1623621585
transform 1 0 36340 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_387
timestamp 1623621585
transform 1 0 36708 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_395
timestamp 1623621585
transform 1 0 37444 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1623621585
transform -1 0 38824 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1623621585
transform 1 0 37812 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_400
timestamp 1623621585
transform 1 0 37904 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_406
timestamp 1623621585
transform 1 0 38456 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1623621585
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1623621585
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input425
timestamp 1623621585
transform 1 0 1380 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1623621585
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1623621585
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_6
timestamp 1623621585
transform 1 0 1656 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_18
timestamp 1623621585
transform 1 0 2760 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1623621585
transform 1 0 3772 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_27
timestamp 1623621585
transform 1 0 3588 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_30
timestamp 1623621585
transform 1 0 3864 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_30
timestamp 1623621585
transform 1 0 3864 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1623621585
transform 1 0 6348 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_42
timestamp 1623621585
transform 1 0 4968 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_54
timestamp 1623621585
transform 1 0 6072 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_42
timestamp 1623621585
transform 1 0 4968 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_54
timestamp 1623621585
transform 1 0 6072 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_58
timestamp 1623621585
transform 1 0 6440 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_66
timestamp 1623621585
transform 1 0 7176 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_78
timestamp 1623621585
transform 1 0 8280 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_70
timestamp 1623621585
transform 1 0 7544 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_82
timestamp 1623621585
transform 1 0 8648 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1623621585
transform 1 0 9016 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_87
timestamp 1623621585
transform 1 0 9108 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_99
timestamp 1623621585
transform 1 0 10212 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_94
timestamp 1623621585
transform 1 0 9752 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1623621585
transform 1 0 11592 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_111
timestamp 1623621585
transform 1 0 11316 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_123
timestamp 1623621585
transform 1 0 12420 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_106
timestamp 1623621585
transform 1 0 10856 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_115
timestamp 1623621585
transform 1 0 11684 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1623621585
transform 1 0 14260 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_135
timestamp 1623621585
transform 1 0 13524 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_144
timestamp 1623621585
transform 1 0 14352 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_127
timestamp 1623621585
transform 1 0 12788 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_139
timestamp 1623621585
transform 1 0 13892 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_156
timestamp 1623621585
transform 1 0 15456 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_151
timestamp 1623621585
transform 1 0 14996 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_163
timestamp 1623621585
transform 1 0 16100 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1623621585
transform 1 0 16836 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_168
timestamp 1623621585
transform 1 0 16560 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_180
timestamp 1623621585
transform 1 0 17664 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_172
timestamp 1623621585
transform 1 0 16928 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_184
timestamp 1623621585
transform 1 0 18032 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1623621585
transform 1 0 19504 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_192
timestamp 1623621585
transform 1 0 18768 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_201
timestamp 1623621585
transform 1 0 19596 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_196
timestamp 1623621585
transform 1 0 19136 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_208
timestamp 1623621585
transform 1 0 20240 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1623621585
transform 1 0 22080 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_213
timestamp 1623621585
transform 1 0 20700 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_225
timestamp 1623621585
transform 1 0 21804 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_220
timestamp 1623621585
transform 1 0 21344 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_229
timestamp 1623621585
transform 1 0 22172 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_237
timestamp 1623621585
transform 1 0 22908 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_249
timestamp 1623621585
transform 1 0 24012 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_241
timestamp 1623621585
transform 1 0 23276 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1623621585
transform 1 0 24748 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_258
timestamp 1623621585
transform 1 0 24840 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_270
timestamp 1623621585
transform 1 0 25944 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_106_253
timestamp 1623621585
transform 1 0 24380 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_265
timestamp 1623621585
transform 1 0 25484 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_2  _0818_
timestamp 1623621585
transform 1 0 26220 0 1 59296
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1623621585
transform 1 0 27324 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_283
timestamp 1623621585
transform 1 0 27140 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_277
timestamp 1623621585
transform 1 0 26588 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_286
timestamp 1623621585
transform 1 0 27416 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_295
timestamp 1623621585
transform 1 0 28244 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_307
timestamp 1623621585
transform 1 0 29348 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_106_298
timestamp 1623621585
transform 1 0 28520 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_310
timestamp 1623621585
transform 1 0 29624 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1623621585
transform 1 0 29992 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_105_313
timestamp 1623621585
transform 1 0 29900 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_315
timestamp 1623621585
transform 1 0 30084 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_327
timestamp 1623621585
transform 1 0 31188 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_322
timestamp 1623621585
transform 1 0 30728 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1623621585
transform 1 0 32568 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_339
timestamp 1623621585
transform 1 0 32292 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_351
timestamp 1623621585
transform 1 0 33396 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_334
timestamp 1623621585
transform 1 0 31832 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_106_343
timestamp 1623621585
transform 1 0 32660 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1623621585
transform 1 0 35236 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_363
timestamp 1623621585
transform 1 0 34500 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_105_372
timestamp 1623621585
transform 1 0 35328 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_355
timestamp 1623621585
transform 1 0 33764 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_367
timestamp 1623621585
transform 1 0 34868 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input205
timestamp 1623621585
transform 1 0 37168 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input234
timestamp 1623621585
transform 1 0 36892 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_384
timestamp 1623621585
transform 1 0 36432 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_388
timestamp 1623621585
transform 1 0 36800 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_392
timestamp 1623621585
transform 1 0 37168 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_379
timestamp 1623621585
transform 1 0 35972 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_391
timestamp 1623621585
transform 1 0 37076 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_395
timestamp 1623621585
transform 1 0 37444 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0428_
timestamp 1623621585
transform 1 0 37536 0 1 59296
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1623621585
transform -1 0 38824 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1623621585
transform -1 0 38824 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1623621585
transform 1 0 37812 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_105_403
timestamp 1623621585
transform 1 0 38180 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_400
timestamp 1623621585
transform 1 0 37904 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_406
timestamp 1623621585
transform 1 0 38456 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1623621585
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input426
timestamp 1623621585
transform 1 0 1380 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_6
timestamp 1623621585
transform 1 0 1656 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_18
timestamp 1623621585
transform 1 0 2760 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1623621585
transform 1 0 3772 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_107_26
timestamp 1623621585
transform 1 0 3496 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_30
timestamp 1623621585
transform 1 0 3864 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_42
timestamp 1623621585
transform 1 0 4968 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_54
timestamp 1623621585
transform 1 0 6072 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_66
timestamp 1623621585
transform 1 0 7176 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_78
timestamp 1623621585
transform 1 0 8280 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1623621585
transform 1 0 9016 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_87
timestamp 1623621585
transform 1 0 9108 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_99
timestamp 1623621585
transform 1 0 10212 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_111
timestamp 1623621585
transform 1 0 11316 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_123
timestamp 1623621585
transform 1 0 12420 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1623621585
transform 1 0 14260 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_135
timestamp 1623621585
transform 1 0 13524 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_144
timestamp 1623621585
transform 1 0 14352 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_156
timestamp 1623621585
transform 1 0 15456 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_168
timestamp 1623621585
transform 1 0 16560 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_180
timestamp 1623621585
transform 1 0 17664 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1623621585
transform 1 0 19504 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_192
timestamp 1623621585
transform 1 0 18768 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_201
timestamp 1623621585
transform 1 0 19596 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_213
timestamp 1623621585
transform 1 0 20700 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_225
timestamp 1623621585
transform 1 0 21804 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_237
timestamp 1623621585
transform 1 0 22908 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_249
timestamp 1623621585
transform 1 0 24012 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_2  _0816_
timestamp 1623621585
transform 1 0 25852 0 1 60384
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1623621585
transform 1 0 24748 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_258
timestamp 1623621585
transform 1 0 24840 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_266
timestamp 1623621585
transform 1 0 25576 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_279
timestamp 1623621585
transform 1 0 26772 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_291
timestamp 1623621585
transform 1 0 27876 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_303
timestamp 1623621585
transform 1 0 28980 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_311
timestamp 1623621585
transform 1 0 29716 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1623621585
transform 1 0 29992 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_315
timestamp 1623621585
transform 1 0 30084 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_327
timestamp 1623621585
transform 1 0 31188 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_339
timestamp 1623621585
transform 1 0 32292 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_351
timestamp 1623621585
transform 1 0 33396 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0956_
timestamp 1623621585
transform 1 0 34224 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1623621585
transform 1 0 35236 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_107_359
timestamp 1623621585
transform 1 0 34132 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_364
timestamp 1623621585
transform 1 0 34592 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_370
timestamp 1623621585
transform 1 0 35144 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_372
timestamp 1623621585
transform 1 0 35328 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input206
timestamp 1623621585
transform 1 0 37260 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_107_384
timestamp 1623621585
transform 1 0 36432 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_392
timestamp 1623621585
transform 1 0 37168 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1623621585
transform -1 0 38824 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input204
timestamp 1623621585
transform 1 0 37904 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_396
timestamp 1623621585
transform 1 0 37536 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_403
timestamp 1623621585
transform 1 0 38180 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1623621585
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1623621585
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1623621585
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_27
timestamp 1623621585
transform 1 0 3588 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_39
timestamp 1623621585
transform 1 0 4692 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1623621585
transform 1 0 6348 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_51
timestamp 1623621585
transform 1 0 5796 0 -1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_108_58
timestamp 1623621585
transform 1 0 6440 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_70
timestamp 1623621585
transform 1 0 7544 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_82
timestamp 1623621585
transform 1 0 8648 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_94
timestamp 1623621585
transform 1 0 9752 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1623621585
transform 1 0 11592 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_106
timestamp 1623621585
transform 1 0 10856 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_115
timestamp 1623621585
transform 1 0 11684 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_127
timestamp 1623621585
transform 1 0 12788 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_139
timestamp 1623621585
transform 1 0 13892 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_151
timestamp 1623621585
transform 1 0 14996 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_163
timestamp 1623621585
transform 1 0 16100 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1623621585
transform 1 0 16836 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_172
timestamp 1623621585
transform 1 0 16928 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_184
timestamp 1623621585
transform 1 0 18032 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_196
timestamp 1623621585
transform 1 0 19136 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_208
timestamp 1623621585
transform 1 0 20240 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1623621585
transform 1 0 22080 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_220
timestamp 1623621585
transform 1 0 21344 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_229
timestamp 1623621585
transform 1 0 22172 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_241
timestamp 1623621585
transform 1 0 23276 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_253
timestamp 1623621585
transform 1 0 24380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_265
timestamp 1623621585
transform 1 0 25484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1623621585
transform 1 0 27324 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_277
timestamp 1623621585
transform 1 0 26588 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_286
timestamp 1623621585
transform 1 0 27416 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_298
timestamp 1623621585
transform 1 0 28520 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_310
timestamp 1623621585
transform 1 0 29624 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_322
timestamp 1623621585
transform 1 0 30728 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1623621585
transform 1 0 32568 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_334
timestamp 1623621585
transform 1 0 31832 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_108_343
timestamp 1623621585
transform 1 0 32660 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_355
timestamp 1623621585
transform 1 0 33764 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_367
timestamp 1623621585
transform 1 0 34868 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input208
timestamp 1623621585
transform 1 0 37168 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_379
timestamp 1623621585
transform 1 0 35972 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_391
timestamp 1623621585
transform 1 0 37076 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_395
timestamp 1623621585
transform 1 0 37444 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1623621585
transform -1 0 38824 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1623621585
transform 1 0 37812 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_400
timestamp 1623621585
transform 1 0 37904 0 -1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_406
timestamp 1623621585
transform 1 0 38456 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1623621585
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input396
timestamp 1623621585
transform 1 0 1380 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_6
timestamp 1623621585
transform 1 0 1656 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_18
timestamp 1623621585
transform 1 0 2760 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1623621585
transform 1 0 3772 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_109_26
timestamp 1623621585
transform 1 0 3496 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_30
timestamp 1623621585
transform 1 0 3864 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_42
timestamp 1623621585
transform 1 0 4968 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_54
timestamp 1623621585
transform 1 0 6072 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_66
timestamp 1623621585
transform 1 0 7176 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_78
timestamp 1623621585
transform 1 0 8280 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1623621585
transform 1 0 9016 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_87
timestamp 1623621585
transform 1 0 9108 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_99
timestamp 1623621585
transform 1 0 10212 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_111
timestamp 1623621585
transform 1 0 11316 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_123
timestamp 1623621585
transform 1 0 12420 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1623621585
transform 1 0 14260 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_135
timestamp 1623621585
transform 1 0 13524 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_144
timestamp 1623621585
transform 1 0 14352 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_156
timestamp 1623621585
transform 1 0 15456 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_168
timestamp 1623621585
transform 1 0 16560 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_180
timestamp 1623621585
transform 1 0 17664 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1623621585
transform 1 0 19504 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_192
timestamp 1623621585
transform 1 0 18768 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_201
timestamp 1623621585
transform 1 0 19596 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_213
timestamp 1623621585
transform 1 0 20700 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_225
timestamp 1623621585
transform 1 0 21804 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_237
timestamp 1623621585
transform 1 0 22908 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_249
timestamp 1623621585
transform 1 0 24012 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1623621585
transform 1 0 24748 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_258
timestamp 1623621585
transform 1 0 24840 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_270
timestamp 1623621585
transform 1 0 25944 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_282
timestamp 1623621585
transform 1 0 27048 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_294
timestamp 1623621585
transform 1 0 28152 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_306
timestamp 1623621585
transform 1 0 29256 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1623621585
transform 1 0 29992 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_315
timestamp 1623621585
transform 1 0 30084 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_327
timestamp 1623621585
transform 1 0 31188 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_339
timestamp 1623621585
transform 1 0 32292 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_351
timestamp 1623621585
transform 1 0 33396 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1623621585
transform 1 0 35236 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_363
timestamp 1623621585
transform 1 0 34500 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_372
timestamp 1623621585
transform 1 0 35328 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input209
timestamp 1623621585
transform 1 0 37260 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_109_384
timestamp 1623621585
transform 1 0 36432 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_392
timestamp 1623621585
transform 1 0 37168 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1623621585
transform -1 0 38824 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input207
timestamp 1623621585
transform 1 0 37904 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_396
timestamp 1623621585
transform 1 0 37536 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_403
timestamp 1623621585
transform 1 0 38180 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1623621585
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input397
timestamp 1623621585
transform 1 0 1380 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_6
timestamp 1623621585
transform 1 0 1656 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_18
timestamp 1623621585
transform 1 0 2760 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_30
timestamp 1623621585
transform 1 0 3864 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1623621585
transform 1 0 6348 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_42
timestamp 1623621585
transform 1 0 4968 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_110_54
timestamp 1623621585
transform 1 0 6072 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_58
timestamp 1623621585
transform 1 0 6440 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_70
timestamp 1623621585
transform 1 0 7544 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_82
timestamp 1623621585
transform 1 0 8648 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_94
timestamp 1623621585
transform 1 0 9752 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1623621585
transform 1 0 11592 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_106
timestamp 1623621585
transform 1 0 10856 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_115
timestamp 1623621585
transform 1 0 11684 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_127
timestamp 1623621585
transform 1 0 12788 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_139
timestamp 1623621585
transform 1 0 13892 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_151
timestamp 1623621585
transform 1 0 14996 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_163
timestamp 1623621585
transform 1 0 16100 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1623621585
transform 1 0 16836 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_172
timestamp 1623621585
transform 1 0 16928 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_184
timestamp 1623621585
transform 1 0 18032 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_196
timestamp 1623621585
transform 1 0 19136 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_208
timestamp 1623621585
transform 1 0 20240 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1623621585
transform 1 0 22080 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_220
timestamp 1623621585
transform 1 0 21344 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_229
timestamp 1623621585
transform 1 0 22172 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_241
timestamp 1623621585
transform 1 0 23276 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_253
timestamp 1623621585
transform 1 0 24380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_265
timestamp 1623621585
transform 1 0 25484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1623621585
transform 1 0 27324 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_277
timestamp 1623621585
transform 1 0 26588 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_110_286
timestamp 1623621585
transform 1 0 27416 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0802_
timestamp 1623621585
transform 1 0 29808 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_298
timestamp 1623621585
transform 1 0 28520 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_110_310
timestamp 1623621585
transform 1 0 29624 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1623621585
transform 1 0 30636 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_316
timestamp 1623621585
transform 1 0 30176 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_320
timestamp 1623621585
transform 1 0 30544 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_325
timestamp 1623621585
transform 1 0 31004 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0807_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 33488 0 -1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1623621585
transform 1 0 32568 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_337
timestamp 1623621585
transform 1 0 32108 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_341
timestamp 1623621585
transform 1 0 32476 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_343
timestamp 1623621585
transform 1 0 32660 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_351
timestamp 1623621585
transform 1 0 33396 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0813_
timestamp 1623621585
transform 1 0 34776 0 -1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_110_359
timestamp 1623621585
transform 1 0 34132 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_365
timestamp 1623621585
transform 1 0 34684 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_373
timestamp 1623621585
transform 1 0 35420 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_385
timestamp 1623621585
transform 1 0 36524 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1623621585
transform -1 0 38824 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1623621585
transform 1 0 37812 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_110_397
timestamp 1623621585
transform 1 0 37628 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_110_400
timestamp 1623621585
transform 1 0 37904 0 -1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_406
timestamp 1623621585
transform 1 0 38456 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1623621585
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1623621585
transform 1 0 1380 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1623621585
transform 1 0 2484 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1623621585
transform 1 0 3772 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_111_27
timestamp 1623621585
transform 1 0 3588 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_30
timestamp 1623621585
transform 1 0 3864 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_42
timestamp 1623621585
transform 1 0 4968 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_54
timestamp 1623621585
transform 1 0 6072 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_66
timestamp 1623621585
transform 1 0 7176 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_78
timestamp 1623621585
transform 1 0 8280 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1623621585
transform 1 0 9016 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_87
timestamp 1623621585
transform 1 0 9108 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_99
timestamp 1623621585
transform 1 0 10212 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_111
timestamp 1623621585
transform 1 0 11316 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_123
timestamp 1623621585
transform 1 0 12420 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1623621585
transform 1 0 14260 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_135
timestamp 1623621585
transform 1 0 13524 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_144
timestamp 1623621585
transform 1 0 14352 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_156
timestamp 1623621585
transform 1 0 15456 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_168
timestamp 1623621585
transform 1 0 16560 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_180
timestamp 1623621585
transform 1 0 17664 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1623621585
transform 1 0 19504 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_192
timestamp 1623621585
transform 1 0 18768 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_201
timestamp 1623621585
transform 1 0 19596 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_213
timestamp 1623621585
transform 1 0 20700 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_225
timestamp 1623621585
transform 1 0 21804 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_237
timestamp 1623621585
transform 1 0 22908 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_249
timestamp 1623621585
transform 1 0 24012 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1623621585
transform 1 0 24748 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_258
timestamp 1623621585
transform 1 0 24840 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_270
timestamp 1623621585
transform 1 0 25944 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_282
timestamp 1623621585
transform 1 0 27048 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_294
timestamp 1623621585
transform 1 0 28152 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_306
timestamp 1623621585
transform 1 0 29256 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1623621585
transform 1 0 29992 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_315
timestamp 1623621585
transform 1 0 30084 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_327
timestamp 1623621585
transform 1 0 31188 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0803_
timestamp 1623621585
transform 1 0 32752 0 1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_111_339
timestamp 1623621585
transform 1 0 32292 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_343
timestamp 1623621585
transform 1 0 32660 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_351
timestamp 1623621585
transform 1 0 33396 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0804_
timestamp 1623621585
transform 1 0 33764 0 1 62560
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1623621585
transform 1 0 35236 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_111_362
timestamp 1623621585
transform 1 0 34408 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_370
timestamp 1623621585
transform 1 0 35144 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_372
timestamp 1623621585
transform 1 0 35328 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input211
timestamp 1623621585
transform 1 0 37260 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_384
timestamp 1623621585
transform 1 0 36432 0 1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_392
timestamp 1623621585
transform 1 0 37168 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1623621585
transform -1 0 38824 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input210
timestamp 1623621585
transform 1 0 37904 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_396
timestamp 1623621585
transform 1 0 37536 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_403
timestamp 1623621585
transform 1 0 38180 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1623621585
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1623621585
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input398
timestamp 1623621585
transform 1 0 1380 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input399
timestamp 1623621585
transform 1 0 1380 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_6
timestamp 1623621585
transform 1 0 1656 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_18
timestamp 1623621585
transform 1 0 2760 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_6
timestamp 1623621585
transform 1 0 1656 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_18
timestamp 1623621585
transform 1 0 2760 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1623621585
transform 1 0 3772 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_30
timestamp 1623621585
transform 1 0 3864 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_113_26
timestamp 1623621585
transform 1 0 3496 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_30
timestamp 1623621585
transform 1 0 3864 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1623621585
transform 1 0 6348 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_42
timestamp 1623621585
transform 1 0 4968 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_54
timestamp 1623621585
transform 1 0 6072 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_58
timestamp 1623621585
transform 1 0 6440 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_42
timestamp 1623621585
transform 1 0 4968 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_54
timestamp 1623621585
transform 1 0 6072 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_70
timestamp 1623621585
transform 1 0 7544 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_82
timestamp 1623621585
transform 1 0 8648 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_66
timestamp 1623621585
transform 1 0 7176 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_78
timestamp 1623621585
transform 1 0 8280 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1623621585
transform 1 0 9016 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_94
timestamp 1623621585
transform 1 0 9752 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_87
timestamp 1623621585
transform 1 0 9108 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_99
timestamp 1623621585
transform 1 0 10212 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1623621585
transform 1 0 11592 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_106
timestamp 1623621585
transform 1 0 10856 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_115
timestamp 1623621585
transform 1 0 11684 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_111
timestamp 1623621585
transform 1 0 11316 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_123
timestamp 1623621585
transform 1 0 12420 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1623621585
transform 1 0 14260 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_127
timestamp 1623621585
transform 1 0 12788 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_139
timestamp 1623621585
transform 1 0 13892 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_135
timestamp 1623621585
transform 1 0 13524 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_113_144
timestamp 1623621585
transform 1 0 14352 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0958_
timestamp 1623621585
transform 1 0 15088 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_112_151
timestamp 1623621585
transform 1 0 14996 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_163
timestamp 1623621585
transform 1 0 16100 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_158
timestamp 1623621585
transform 1 0 15640 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1623621585
transform 1 0 16836 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_172
timestamp 1623621585
transform 1 0 16928 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_184
timestamp 1623621585
transform 1 0 18032 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_170
timestamp 1623621585
transform 1 0 16744 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_182
timestamp 1623621585
transform 1 0 17848 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1623621585
transform 1 0 19504 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_196
timestamp 1623621585
transform 1 0 19136 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_208
timestamp 1623621585
transform 1 0 20240 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_194
timestamp 1623621585
transform 1 0 18952 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_113_201
timestamp 1623621585
transform 1 0 19596 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1623621585
transform 1 0 22080 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_220
timestamp 1623621585
transform 1 0 21344 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_229
timestamp 1623621585
transform 1 0 22172 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_213
timestamp 1623621585
transform 1 0 20700 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_225
timestamp 1623621585
transform 1 0 21804 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_241
timestamp 1623621585
transform 1 0 23276 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_237
timestamp 1623621585
transform 1 0 22908 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_249
timestamp 1623621585
transform 1 0 24012 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1623621585
transform 1 0 24748 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_253
timestamp 1623621585
transform 1 0 24380 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_265
timestamp 1623621585
transform 1 0 25484 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_258
timestamp 1623621585
transform 1 0 24840 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_270
timestamp 1623621585
transform 1 0 25944 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1623621585
transform 1 0 27324 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_277
timestamp 1623621585
transform 1 0 26588 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_112_286
timestamp 1623621585
transform 1 0 27416 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_282
timestamp 1623621585
transform 1 0 27048 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_298
timestamp 1623621585
transform 1 0 28520 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_310
timestamp 1623621585
transform 1 0 29624 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_294
timestamp 1623621585
transform 1 0 28152 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_306
timestamp 1623621585
transform 1 0 29256 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1623621585
transform 1 0 29992 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_322
timestamp 1623621585
transform 1 0 30728 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_315
timestamp 1623621585
transform 1 0 30084 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_327
timestamp 1623621585
transform 1 0 31188 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0805_
timestamp 1623621585
transform 1 0 33120 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1623621585
transform 1 0 32568 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_334
timestamp 1623621585
transform 1 0 31832 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_112_343
timestamp 1623621585
transform 1 0 32660 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_347
timestamp 1623621585
transform 1 0 33028 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_339
timestamp 1623621585
transform 1 0 32292 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_351
timestamp 1623621585
transform 1 0 33396 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0806_
timestamp 1623621585
transform 1 0 34132 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0809_
timestamp 1623621585
transform 1 0 33948 0 1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0810_
timestamp 1623621585
transform 1 0 35144 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1623621585
transform 1 0 35236 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_355
timestamp 1623621585
transform 1 0 33764 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_366
timestamp 1623621585
transform 1 0 34776 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_113_364
timestamp 1623621585
transform 1 0 34592 0 1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_370
timestamp 1623621585
transform 1 0 35144 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_372
timestamp 1623621585
transform 1 0 35328 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0812_
timestamp 1623621585
transform 1 0 36156 0 -1 63648
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input213
timestamp 1623621585
transform 1 0 37168 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input215
timestamp 1623621585
transform 1 0 37260 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_377
timestamp 1623621585
transform 1 0 35788 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_388
timestamp 1623621585
transform 1 0 36800 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_395
timestamp 1623621585
transform 1 0 37444 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_113_384
timestamp 1623621585
transform 1 0 36432 0 1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_113_392
timestamp 1623621585
transform 1 0 37168 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1623621585
transform -1 0 38824 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1623621585
transform -1 0 38824 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1623621585
transform 1 0 37812 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input212
timestamp 1623621585
transform 1 0 37904 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_112_400
timestamp 1623621585
transform 1 0 37904 0 -1 63648
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_406
timestamp 1623621585
transform 1 0 38456 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_113_396
timestamp 1623621585
transform 1 0 37536 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_403
timestamp 1623621585
transform 1 0 38180 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1623621585
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1623621585
transform 1 0 1380 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1623621585
transform 1 0 2484 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_27
timestamp 1623621585
transform 1 0 3588 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_39
timestamp 1623621585
transform 1 0 4692 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1623621585
transform 1 0 6348 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_51
timestamp 1623621585
transform 1 0 5796 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_114_58
timestamp 1623621585
transform 1 0 6440 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_70
timestamp 1623621585
transform 1 0 7544 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_82
timestamp 1623621585
transform 1 0 8648 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_94
timestamp 1623621585
transform 1 0 9752 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1623621585
transform 1 0 11592 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_106
timestamp 1623621585
transform 1 0 10856 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_115
timestamp 1623621585
transform 1 0 11684 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_127
timestamp 1623621585
transform 1 0 12788 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_139
timestamp 1623621585
transform 1 0 13892 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_151
timestamp 1623621585
transform 1 0 14996 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_163
timestamp 1623621585
transform 1 0 16100 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1623621585
transform 1 0 16836 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_172
timestamp 1623621585
transform 1 0 16928 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_184
timestamp 1623621585
transform 1 0 18032 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_196
timestamp 1623621585
transform 1 0 19136 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_208
timestamp 1623621585
transform 1 0 20240 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1623621585
transform 1 0 22080 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_220
timestamp 1623621585
transform 1 0 21344 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_229
timestamp 1623621585
transform 1 0 22172 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_241
timestamp 1623621585
transform 1 0 23276 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_253
timestamp 1623621585
transform 1 0 24380 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_265
timestamp 1623621585
transform 1 0 25484 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1623621585
transform 1 0 27324 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_277
timestamp 1623621585
transform 1 0 26588 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_286
timestamp 1623621585
transform 1 0 27416 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_298
timestamp 1623621585
transform 1 0 28520 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_310
timestamp 1623621585
transform 1 0 29624 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_322
timestamp 1623621585
transform 1 0 30728 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1623621585
transform 1 0 32568 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_334
timestamp 1623621585
transform 1 0 31832 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_114_343
timestamp 1623621585
transform 1 0 32660 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0811_
timestamp 1623621585
transform 1 0 34316 0 -1 64736
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_114_355
timestamp 1623621585
transform 1 0 33764 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_114_368
timestamp 1623621585
transform 1 0 34960 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_380
timestamp 1623621585
transform 1 0 36064 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_392
timestamp 1623621585
transform 1 0 37168 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1623621585
transform -1 0 38824 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1623621585
transform 1 0 37812 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_114_398
timestamp 1623621585
transform 1 0 37720 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_114_400
timestamp 1623621585
transform 1 0 37904 0 -1 64736
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_406
timestamp 1623621585
transform 1 0 38456 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1623621585
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input400
timestamp 1623621585
transform 1 0 1380 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_6
timestamp 1623621585
transform 1 0 1656 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_18
timestamp 1623621585
transform 1 0 2760 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1623621585
transform 1 0 3772 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_115_26
timestamp 1623621585
transform 1 0 3496 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_30
timestamp 1623621585
transform 1 0 3864 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_42
timestamp 1623621585
transform 1 0 4968 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_54
timestamp 1623621585
transform 1 0 6072 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_66
timestamp 1623621585
transform 1 0 7176 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_78
timestamp 1623621585
transform 1 0 8280 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1623621585
transform 1 0 9016 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_87
timestamp 1623621585
transform 1 0 9108 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_99
timestamp 1623621585
transform 1 0 10212 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_111
timestamp 1623621585
transform 1 0 11316 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_123
timestamp 1623621585
transform 1 0 12420 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1623621585
transform 1 0 14260 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_135
timestamp 1623621585
transform 1 0 13524 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_144
timestamp 1623621585
transform 1 0 14352 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_156
timestamp 1623621585
transform 1 0 15456 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_168
timestamp 1623621585
transform 1 0 16560 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_180
timestamp 1623621585
transform 1 0 17664 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1623621585
transform 1 0 19504 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_192
timestamp 1623621585
transform 1 0 18768 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_201
timestamp 1623621585
transform 1 0 19596 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_213
timestamp 1623621585
transform 1 0 20700 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_225
timestamp 1623621585
transform 1 0 21804 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_237
timestamp 1623621585
transform 1 0 22908 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_249
timestamp 1623621585
transform 1 0 24012 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1623621585
transform 1 0 24748 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_258
timestamp 1623621585
transform 1 0 24840 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_270
timestamp 1623621585
transform 1 0 25944 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_282
timestamp 1623621585
transform 1 0 27048 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_294
timestamp 1623621585
transform 1 0 28152 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_306
timestamp 1623621585
transform 1 0 29256 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1623621585
transform 1 0 29992 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_315
timestamp 1623621585
transform 1 0 30084 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_327
timestamp 1623621585
transform 1 0 31188 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_339
timestamp 1623621585
transform 1 0 32292 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_351
timestamp 1623621585
transform 1 0 33396 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1623621585
transform 1 0 35236 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_363
timestamp 1623621585
transform 1 0 34500 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_115_372
timestamp 1623621585
transform 1 0 35328 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input217
timestamp 1623621585
transform 1 0 37260 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_115_384
timestamp 1623621585
transform 1 0 36432 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_115_392
timestamp 1623621585
transform 1 0 37168 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1623621585
transform -1 0 38824 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input216
timestamp 1623621585
transform 1 0 37904 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_396
timestamp 1623621585
transform 1 0 37536 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_403
timestamp 1623621585
transform 1 0 38180 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1623621585
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input401
timestamp 1623621585
transform 1 0 1380 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_6
timestamp 1623621585
transform 1 0 1656 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_18
timestamp 1623621585
transform 1 0 2760 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_30
timestamp 1623621585
transform 1 0 3864 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1623621585
transform 1 0 6348 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_42
timestamp 1623621585
transform 1 0 4968 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_54
timestamp 1623621585
transform 1 0 6072 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_58
timestamp 1623621585
transform 1 0 6440 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_70
timestamp 1623621585
transform 1 0 7544 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_82
timestamp 1623621585
transform 1 0 8648 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_94
timestamp 1623621585
transform 1 0 9752 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1623621585
transform 1 0 11592 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_106
timestamp 1623621585
transform 1 0 10856 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_115
timestamp 1623621585
transform 1 0 11684 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_127
timestamp 1623621585
transform 1 0 12788 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_139
timestamp 1623621585
transform 1 0 13892 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_151
timestamp 1623621585
transform 1 0 14996 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_163
timestamp 1623621585
transform 1 0 16100 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1623621585
transform 1 0 16836 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_172
timestamp 1623621585
transform 1 0 16928 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_184
timestamp 1623621585
transform 1 0 18032 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_196
timestamp 1623621585
transform 1 0 19136 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_208
timestamp 1623621585
transform 1 0 20240 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1623621585
transform 1 0 22080 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_220
timestamp 1623621585
transform 1 0 21344 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_229
timestamp 1623621585
transform 1 0 22172 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_241
timestamp 1623621585
transform 1 0 23276 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_253
timestamp 1623621585
transform 1 0 24380 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_265
timestamp 1623621585
transform 1 0 25484 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1623621585
transform 1 0 27324 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_277
timestamp 1623621585
transform 1 0 26588 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_286
timestamp 1623621585
transform 1 0 27416 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_298
timestamp 1623621585
transform 1 0 28520 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_310
timestamp 1623621585
transform 1 0 29624 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_322
timestamp 1623621585
transform 1 0 30728 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1623621585
transform 1 0 32568 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_334
timestamp 1623621585
transform 1 0 31832 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_116_343
timestamp 1623621585
transform 1 0 32660 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_355
timestamp 1623621585
transform 1 0 33764 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_367
timestamp 1623621585
transform 1 0 34868 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input219
timestamp 1623621585
transform 1 0 37168 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_379
timestamp 1623621585
transform 1 0 35972 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_391
timestamp 1623621585
transform 1 0 37076 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_116_395
timestamp 1623621585
transform 1 0 37444 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1623621585
transform -1 0 38824 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1623621585
transform 1 0 37812 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_400
timestamp 1623621585
transform 1 0 37904 0 -1 65824
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_406
timestamp 1623621585
transform 1 0 38456 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1623621585
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_3
timestamp 1623621585
transform 1 0 1380 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_15
timestamp 1623621585
transform 1 0 2484 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1623621585
transform 1 0 3772 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_117_27
timestamp 1623621585
transform 1 0 3588 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_117_30
timestamp 1623621585
transform 1 0 3864 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_42
timestamp 1623621585
transform 1 0 4968 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_54
timestamp 1623621585
transform 1 0 6072 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_66
timestamp 1623621585
transform 1 0 7176 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_78
timestamp 1623621585
transform 1 0 8280 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1623621585
transform 1 0 9016 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_87
timestamp 1623621585
transform 1 0 9108 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_99
timestamp 1623621585
transform 1 0 10212 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_111
timestamp 1623621585
transform 1 0 11316 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_123
timestamp 1623621585
transform 1 0 12420 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1623621585
transform 1 0 14260 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_135
timestamp 1623621585
transform 1 0 13524 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_144
timestamp 1623621585
transform 1 0 14352 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_156
timestamp 1623621585
transform 1 0 15456 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_168
timestamp 1623621585
transform 1 0 16560 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_180
timestamp 1623621585
transform 1 0 17664 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1623621585
transform 1 0 19504 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_192
timestamp 1623621585
transform 1 0 18768 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_201
timestamp 1623621585
transform 1 0 19596 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_213
timestamp 1623621585
transform 1 0 20700 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1623621585
transform 1 0 21804 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_237
timestamp 1623621585
transform 1 0 22908 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_249
timestamp 1623621585
transform 1 0 24012 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1623621585
transform 1 0 24748 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_258
timestamp 1623621585
transform 1 0 24840 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_270
timestamp 1623621585
transform 1 0 25944 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_282
timestamp 1623621585
transform 1 0 27048 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_294
timestamp 1623621585
transform 1 0 28152 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_306
timestamp 1623621585
transform 1 0 29256 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1623621585
transform 1 0 29992 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_315
timestamp 1623621585
transform 1 0 30084 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_327
timestamp 1623621585
transform 1 0 31188 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_339
timestamp 1623621585
transform 1 0 32292 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_351
timestamp 1623621585
transform 1 0 33396 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1623621585
transform 1 0 35236 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_363
timestamp 1623621585
transform 1 0 34500 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_372
timestamp 1623621585
transform 1 0 35328 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input220
timestamp 1623621585
transform 1 0 37260 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_117_384
timestamp 1623621585
transform 1 0 36432 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_392
timestamp 1623621585
transform 1 0 37168 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1623621585
transform -1 0 38824 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input218
timestamp 1623621585
transform 1 0 37904 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_396
timestamp 1623621585
transform 1 0 37536 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_117_403
timestamp 1623621585
transform 1 0 38180 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1623621585
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1623621585
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input402
timestamp 1623621585
transform 1 0 1380 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input403
timestamp 1623621585
transform 1 0 1380 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_6
timestamp 1623621585
transform 1 0 1656 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_18
timestamp 1623621585
transform 1 0 2760 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_6
timestamp 1623621585
transform 1 0 1656 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_18
timestamp 1623621585
transform 1 0 2760 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1623621585
transform 1 0 3772 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_30
timestamp 1623621585
transform 1 0 3864 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_26
timestamp 1623621585
transform 1 0 3496 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_30
timestamp 1623621585
transform 1 0 3864 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1623621585
transform 1 0 6348 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_42
timestamp 1623621585
transform 1 0 4968 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_118_54
timestamp 1623621585
transform 1 0 6072 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_58
timestamp 1623621585
transform 1 0 6440 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_42
timestamp 1623621585
transform 1 0 4968 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_54
timestamp 1623621585
transform 1 0 6072 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_70
timestamp 1623621585
transform 1 0 7544 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_82
timestamp 1623621585
transform 1 0 8648 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_66
timestamp 1623621585
transform 1 0 7176 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_78
timestamp 1623621585
transform 1 0 8280 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1623621585
transform 1 0 9016 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_94
timestamp 1623621585
transform 1 0 9752 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_87
timestamp 1623621585
transform 1 0 9108 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_99
timestamp 1623621585
transform 1 0 10212 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1623621585
transform 1 0 11592 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_106
timestamp 1623621585
transform 1 0 10856 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_115
timestamp 1623621585
transform 1 0 11684 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_111
timestamp 1623621585
transform 1 0 11316 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_123
timestamp 1623621585
transform 1 0 12420 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1623621585
transform 1 0 14260 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_127
timestamp 1623621585
transform 1 0 12788 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_139
timestamp 1623621585
transform 1 0 13892 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_135
timestamp 1623621585
transform 1 0 13524 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_144
timestamp 1623621585
transform 1 0 14352 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_151
timestamp 1623621585
transform 1 0 14996 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_163
timestamp 1623621585
transform 1 0 16100 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_156
timestamp 1623621585
transform 1 0 15456 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1623621585
transform 1 0 16836 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_172
timestamp 1623621585
transform 1 0 16928 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_184
timestamp 1623621585
transform 1 0 18032 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_168
timestamp 1623621585
transform 1 0 16560 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_180
timestamp 1623621585
transform 1 0 17664 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1623621585
transform 1 0 19504 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_196
timestamp 1623621585
transform 1 0 19136 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_208
timestamp 1623621585
transform 1 0 20240 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_192
timestamp 1623621585
transform 1 0 18768 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_201
timestamp 1623621585
transform 1 0 19596 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1623621585
transform 1 0 22080 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_220
timestamp 1623621585
transform 1 0 21344 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_229
timestamp 1623621585
transform 1 0 22172 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_213
timestamp 1623621585
transform 1 0 20700 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_225
timestamp 1623621585
transform 1 0 21804 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_241
timestamp 1623621585
transform 1 0 23276 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_237
timestamp 1623621585
transform 1 0 22908 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_249
timestamp 1623621585
transform 1 0 24012 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1623621585
transform 1 0 24748 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_253
timestamp 1623621585
transform 1 0 24380 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_265
timestamp 1623621585
transform 1 0 25484 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_258
timestamp 1623621585
transform 1 0 24840 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_270
timestamp 1623621585
transform 1 0 25944 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1623621585
transform 1 0 27324 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_277
timestamp 1623621585
transform 1 0 26588 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_286
timestamp 1623621585
transform 1 0 27416 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_282
timestamp 1623621585
transform 1 0 27048 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_298
timestamp 1623621585
transform 1 0 28520 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_310
timestamp 1623621585
transform 1 0 29624 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_294
timestamp 1623621585
transform 1 0 28152 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_306
timestamp 1623621585
transform 1 0 29256 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1623621585
transform 1 0 29992 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_322
timestamp 1623621585
transform 1 0 30728 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_315
timestamp 1623621585
transform 1 0 30084 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_327
timestamp 1623621585
transform 1 0 31188 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1623621585
transform 1 0 32568 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_334
timestamp 1623621585
transform 1 0 31832 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_343
timestamp 1623621585
transform 1 0 32660 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_339
timestamp 1623621585
transform 1 0 32292 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_351
timestamp 1623621585
transform 1 0 33396 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1623621585
transform 1 0 35236 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_355
timestamp 1623621585
transform 1 0 33764 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_367
timestamp 1623621585
transform 1 0 34868 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_363
timestamp 1623621585
transform 1 0 34500 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_372
timestamp 1623621585
transform 1 0 35328 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input222
timestamp 1623621585
transform 1 0 37260 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_379
timestamp 1623621585
transform 1 0 35972 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_391
timestamp 1623621585
transform 1 0 37076 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_119_384
timestamp 1623621585
transform 1 0 36432 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_119_392
timestamp 1623621585
transform 1 0 37168 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1623621585
transform -1 0 38824 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1623621585
transform -1 0 38824 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1623621585
transform 1 0 37812 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input221
timestamp 1623621585
transform 1 0 37904 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_118_400
timestamp 1623621585
transform 1 0 37904 0 -1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_406
timestamp 1623621585
transform 1 0 38456 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_119_396
timestamp 1623621585
transform 1 0 37536 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_403
timestamp 1623621585
transform 1 0 38180 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1623621585
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1623621585
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1623621585
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_27
timestamp 1623621585
transform 1 0 3588 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_39
timestamp 1623621585
transform 1 0 4692 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1623621585
transform 1 0 6348 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_51
timestamp 1623621585
transform 1 0 5796 0 -1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_120_58
timestamp 1623621585
transform 1 0 6440 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_70
timestamp 1623621585
transform 1 0 7544 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_82
timestamp 1623621585
transform 1 0 8648 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_94
timestamp 1623621585
transform 1 0 9752 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1623621585
transform 1 0 11592 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_106
timestamp 1623621585
transform 1 0 10856 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_115
timestamp 1623621585
transform 1 0 11684 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_127
timestamp 1623621585
transform 1 0 12788 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_139
timestamp 1623621585
transform 1 0 13892 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_151
timestamp 1623621585
transform 1 0 14996 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_163
timestamp 1623621585
transform 1 0 16100 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1623621585
transform 1 0 16836 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_172
timestamp 1623621585
transform 1 0 16928 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_184
timestamp 1623621585
transform 1 0 18032 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_196
timestamp 1623621585
transform 1 0 19136 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_208
timestamp 1623621585
transform 1 0 20240 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1623621585
transform 1 0 22080 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_220
timestamp 1623621585
transform 1 0 21344 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_229
timestamp 1623621585
transform 1 0 22172 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_241
timestamp 1623621585
transform 1 0 23276 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_253
timestamp 1623621585
transform 1 0 24380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_265
timestamp 1623621585
transform 1 0 25484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1623621585
transform 1 0 27324 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_277
timestamp 1623621585
transform 1 0 26588 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_286
timestamp 1623621585
transform 1 0 27416 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_298
timestamp 1623621585
transform 1 0 28520 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_310
timestamp 1623621585
transform 1 0 29624 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_322
timestamp 1623621585
transform 1 0 30728 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1623621585
transform 1 0 32568 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_334
timestamp 1623621585
transform 1 0 31832 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_120_343
timestamp 1623621585
transform 1 0 32660 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_355
timestamp 1623621585
transform 1 0 33764 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_367
timestamp 1623621585
transform 1 0 34868 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input224
timestamp 1623621585
transform 1 0 37168 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_379
timestamp 1623621585
transform 1 0 35972 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_391
timestamp 1623621585
transform 1 0 37076 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_395
timestamp 1623621585
transform 1 0 37444 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1623621585
transform -1 0 38824 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1623621585
transform 1 0 37812 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_400
timestamp 1623621585
transform 1 0 37904 0 -1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_406
timestamp 1623621585
transform 1 0 38456 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1623621585
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input404
timestamp 1623621585
transform 1 0 1748 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_121_3
timestamp 1623621585
transform 1 0 1380 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_11
timestamp 1623621585
transform 1 0 2116 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1623621585
transform 1 0 3772 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_121_23
timestamp 1623621585
transform 1 0 3220 0 1 68000
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_121_30
timestamp 1623621585
transform 1 0 3864 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_42
timestamp 1623621585
transform 1 0 4968 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_54
timestamp 1623621585
transform 1 0 6072 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_66
timestamp 1623621585
transform 1 0 7176 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_78
timestamp 1623621585
transform 1 0 8280 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1623621585
transform 1 0 9016 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_87
timestamp 1623621585
transform 1 0 9108 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_99
timestamp 1623621585
transform 1 0 10212 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_111
timestamp 1623621585
transform 1 0 11316 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_123
timestamp 1623621585
transform 1 0 12420 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1623621585
transform 1 0 14260 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_135
timestamp 1623621585
transform 1 0 13524 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_144
timestamp 1623621585
transform 1 0 14352 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_156
timestamp 1623621585
transform 1 0 15456 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_168
timestamp 1623621585
transform 1 0 16560 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_180
timestamp 1623621585
transform 1 0 17664 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1623621585
transform 1 0 19504 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_192
timestamp 1623621585
transform 1 0 18768 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_201
timestamp 1623621585
transform 1 0 19596 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_213
timestamp 1623621585
transform 1 0 20700 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_225
timestamp 1623621585
transform 1 0 21804 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_237
timestamp 1623621585
transform 1 0 22908 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_249
timestamp 1623621585
transform 1 0 24012 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1623621585
transform 1 0 24748 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_258
timestamp 1623621585
transform 1 0 24840 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_270
timestamp 1623621585
transform 1 0 25944 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_282
timestamp 1623621585
transform 1 0 27048 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_294
timestamp 1623621585
transform 1 0 28152 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_121_306
timestamp 1623621585
transform 1 0 29256 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1623621585
transform 1 0 29992 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_315
timestamp 1623621585
transform 1 0 30084 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_327
timestamp 1623621585
transform 1 0 31188 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_339
timestamp 1623621585
transform 1 0 32292 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_351
timestamp 1623621585
transform 1 0 33396 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1623621585
transform 1 0 35236 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_363
timestamp 1623621585
transform 1 0 34500 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_372
timestamp 1623621585
transform 1 0 35328 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input226
timestamp 1623621585
transform 1 0 37260 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_121_384
timestamp 1623621585
transform 1 0 36432 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_121_392
timestamp 1623621585
transform 1 0 37168 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1623621585
transform -1 0 38824 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input223
timestamp 1623621585
transform 1 0 37904 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_396
timestamp 1623621585
transform 1 0 37536 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_121_403
timestamp 1623621585
transform 1 0 38180 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1623621585
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input405
timestamp 1623621585
transform 1 0 1748 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_122_3
timestamp 1623621585
transform 1 0 1380 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_11
timestamp 1623621585
transform 1 0 2116 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_23
timestamp 1623621585
transform 1 0 3220 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_35
timestamp 1623621585
transform 1 0 4324 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1623621585
transform 1 0 6348 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_47
timestamp 1623621585
transform 1 0 5428 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_55
timestamp 1623621585
transform 1 0 6164 0 -1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_122_58
timestamp 1623621585
transform 1 0 6440 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_70
timestamp 1623621585
transform 1 0 7544 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_82
timestamp 1623621585
transform 1 0 8648 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_94
timestamp 1623621585
transform 1 0 9752 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1623621585
transform 1 0 11592 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_106
timestamp 1623621585
transform 1 0 10856 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_115
timestamp 1623621585
transform 1 0 11684 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_127
timestamp 1623621585
transform 1 0 12788 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_139
timestamp 1623621585
transform 1 0 13892 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_151
timestamp 1623621585
transform 1 0 14996 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_163
timestamp 1623621585
transform 1 0 16100 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1623621585
transform 1 0 16836 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_172
timestamp 1623621585
transform 1 0 16928 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_184
timestamp 1623621585
transform 1 0 18032 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_196
timestamp 1623621585
transform 1 0 19136 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_208
timestamp 1623621585
transform 1 0 20240 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1623621585
transform 1 0 22080 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_220
timestamp 1623621585
transform 1 0 21344 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_229
timestamp 1623621585
transform 1 0 22172 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_241
timestamp 1623621585
transform 1 0 23276 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_253
timestamp 1623621585
transform 1 0 24380 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_265
timestamp 1623621585
transform 1 0 25484 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1623621585
transform 1 0 27324 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_277
timestamp 1623621585
transform 1 0 26588 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_286
timestamp 1623621585
transform 1 0 27416 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_298
timestamp 1623621585
transform 1 0 28520 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_310
timestamp 1623621585
transform 1 0 29624 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_322
timestamp 1623621585
transform 1 0 30728 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1623621585
transform 1 0 32568 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_334
timestamp 1623621585
transform 1 0 31832 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_343
timestamp 1623621585
transform 1 0 32660 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_355
timestamp 1623621585
transform 1 0 33764 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_367
timestamp 1623621585
transform 1 0 34868 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input227
timestamp 1623621585
transform 1 0 37168 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_379
timestamp 1623621585
transform 1 0 35972 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_391
timestamp 1623621585
transform 1 0 37076 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_395
timestamp 1623621585
transform 1 0 37444 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1623621585
transform -1 0 38824 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1623621585
transform 1 0 37812 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_400
timestamp 1623621585
transform 1 0 37904 0 -1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_406
timestamp 1623621585
transform 1 0 38456 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1623621585
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1623621585
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1623621585
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1623621585
transform 1 0 3772 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_123_27
timestamp 1623621585
transform 1 0 3588 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_30
timestamp 1623621585
transform 1 0 3864 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_42
timestamp 1623621585
transform 1 0 4968 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_54
timestamp 1623621585
transform 1 0 6072 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_66
timestamp 1623621585
transform 1 0 7176 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_78
timestamp 1623621585
transform 1 0 8280 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1623621585
transform 1 0 9016 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_87
timestamp 1623621585
transform 1 0 9108 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_99
timestamp 1623621585
transform 1 0 10212 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_111
timestamp 1623621585
transform 1 0 11316 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_123
timestamp 1623621585
transform 1 0 12420 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1623621585
transform 1 0 14260 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_135
timestamp 1623621585
transform 1 0 13524 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_144
timestamp 1623621585
transform 1 0 14352 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_156
timestamp 1623621585
transform 1 0 15456 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_168
timestamp 1623621585
transform 1 0 16560 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_180
timestamp 1623621585
transform 1 0 17664 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1623621585
transform 1 0 19504 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_192
timestamp 1623621585
transform 1 0 18768 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_201
timestamp 1623621585
transform 1 0 19596 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_213
timestamp 1623621585
transform 1 0 20700 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_225
timestamp 1623621585
transform 1 0 21804 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_237
timestamp 1623621585
transform 1 0 22908 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_249
timestamp 1623621585
transform 1 0 24012 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1296
timestamp 1623621585
transform 1 0 24748 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_258
timestamp 1623621585
transform 1 0 24840 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_270
timestamp 1623621585
transform 1 0 25944 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_282
timestamp 1623621585
transform 1 0 27048 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_294
timestamp 1623621585
transform 1 0 28152 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_306
timestamp 1623621585
transform 1 0 29256 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1297
timestamp 1623621585
transform 1 0 29992 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_315
timestamp 1623621585
transform 1 0 30084 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_327
timestamp 1623621585
transform 1 0 31188 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_339
timestamp 1623621585
transform 1 0 32292 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_351
timestamp 1623621585
transform 1 0 33396 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1298
timestamp 1623621585
transform 1 0 35236 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_363
timestamp 1623621585
transform 1 0 34500 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_123_372
timestamp 1623621585
transform 1 0 35328 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input246
timestamp 1623621585
transform 1 0 37076 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_123_384
timestamp 1623621585
transform 1 0 36432 0 1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_390
timestamp 1623621585
transform 1 0 36984 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_395
timestamp 1623621585
transform 1 0 37444 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1623621585
transform -1 0 38824 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1623621585
transform 1 0 37812 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_403
timestamp 1623621585
transform 1 0 38180 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1623621585
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input407
timestamp 1623621585
transform 1 0 1748 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_3
timestamp 1623621585
transform 1 0 1380 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_11
timestamp 1623621585
transform 1 0 2116 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_23
timestamp 1623621585
transform 1 0 3220 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_35
timestamp 1623621585
transform 1 0 4324 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1299
timestamp 1623621585
transform 1 0 6348 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_47
timestamp 1623621585
transform 1 0 5428 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_124_55
timestamp 1623621585
transform 1 0 6164 0 -1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_124_58
timestamp 1623621585
transform 1 0 6440 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_70
timestamp 1623621585
transform 1 0 7544 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_82
timestamp 1623621585
transform 1 0 8648 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_94
timestamp 1623621585
transform 1 0 9752 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1300
timestamp 1623621585
transform 1 0 11592 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_106
timestamp 1623621585
transform 1 0 10856 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_115
timestamp 1623621585
transform 1 0 11684 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_127
timestamp 1623621585
transform 1 0 12788 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_139
timestamp 1623621585
transform 1 0 13892 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_151
timestamp 1623621585
transform 1 0 14996 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_163
timestamp 1623621585
transform 1 0 16100 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1301
timestamp 1623621585
transform 1 0 16836 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_172
timestamp 1623621585
transform 1 0 16928 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_184
timestamp 1623621585
transform 1 0 18032 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_196
timestamp 1623621585
transform 1 0 19136 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_208
timestamp 1623621585
transform 1 0 20240 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1302
timestamp 1623621585
transform 1 0 22080 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_220
timestamp 1623621585
transform 1 0 21344 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_229
timestamp 1623621585
transform 1 0 22172 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_241
timestamp 1623621585
transform 1 0 23276 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_253
timestamp 1623621585
transform 1 0 24380 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_265
timestamp 1623621585
transform 1 0 25484 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1303
timestamp 1623621585
transform 1 0 27324 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_277
timestamp 1623621585
transform 1 0 26588 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_286
timestamp 1623621585
transform 1 0 27416 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_298
timestamp 1623621585
transform 1 0 28520 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_310
timestamp 1623621585
transform 1 0 29624 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_322
timestamp 1623621585
transform 1 0 30728 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1304
timestamp 1623621585
transform 1 0 32568 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_334
timestamp 1623621585
transform 1 0 31832 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_124_343
timestamp 1623621585
transform 1 0 32660 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_355
timestamp 1623621585
transform 1 0 33764 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_367
timestamp 1623621585
transform 1 0 34868 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input257
timestamp 1623621585
transform 1 0 37076 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_379
timestamp 1623621585
transform 1 0 35972 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_395
timestamp 1623621585
transform 1 0 37444 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1623621585
transform -1 0 38824 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1305
timestamp 1623621585
transform 1 0 37812 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_400
timestamp 1623621585
transform 1 0 37904 0 -1 70176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_406
timestamp 1623621585
transform 1 0 38456 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1623621585
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1623621585
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input408
timestamp 1623621585
transform 1 0 1748 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_3
timestamp 1623621585
transform 1 0 1380 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_15
timestamp 1623621585
transform 1 0 2484 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_3
timestamp 1623621585
transform 1 0 1380 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_11
timestamp 1623621585
transform 1 0 2116 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1306
timestamp 1623621585
transform 1 0 3772 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_125_27
timestamp 1623621585
transform 1 0 3588 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1623621585
transform 1 0 3864 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_23
timestamp 1623621585
transform 1 0 3220 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_35
timestamp 1623621585
transform 1 0 4324 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1313
timestamp 1623621585
transform 1 0 6348 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1623621585
transform 1 0 4968 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_54
timestamp 1623621585
transform 1 0 6072 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_47
timestamp 1623621585
transform 1 0 5428 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_55
timestamp 1623621585
transform 1 0 6164 0 -1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_126_58
timestamp 1623621585
transform 1 0 6440 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_66
timestamp 1623621585
transform 1 0 7176 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_78
timestamp 1623621585
transform 1 0 8280 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_70
timestamp 1623621585
transform 1 0 7544 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_82
timestamp 1623621585
transform 1 0 8648 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1307
timestamp 1623621585
transform 1 0 9016 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_87
timestamp 1623621585
transform 1 0 9108 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_99
timestamp 1623621585
transform 1 0 10212 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_94
timestamp 1623621585
transform 1 0 9752 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1314
timestamp 1623621585
transform 1 0 11592 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_111
timestamp 1623621585
transform 1 0 11316 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_123
timestamp 1623621585
transform 1 0 12420 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_106
timestamp 1623621585
transform 1 0 10856 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_115
timestamp 1623621585
transform 1 0 11684 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1308
timestamp 1623621585
transform 1 0 14260 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_135
timestamp 1623621585
transform 1 0 13524 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_144
timestamp 1623621585
transform 1 0 14352 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_127
timestamp 1623621585
transform 1 0 12788 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_139
timestamp 1623621585
transform 1 0 13892 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_156
timestamp 1623621585
transform 1 0 15456 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_151
timestamp 1623621585
transform 1 0 14996 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_163
timestamp 1623621585
transform 1 0 16100 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1315
timestamp 1623621585
transform 1 0 16836 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_168
timestamp 1623621585
transform 1 0 16560 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_180
timestamp 1623621585
transform 1 0 17664 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_172
timestamp 1623621585
transform 1 0 16928 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_184
timestamp 1623621585
transform 1 0 18032 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1309
timestamp 1623621585
transform 1 0 19504 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_192
timestamp 1623621585
transform 1 0 18768 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_201
timestamp 1623621585
transform 1 0 19596 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_196
timestamp 1623621585
transform 1 0 19136 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_208
timestamp 1623621585
transform 1 0 20240 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1316
timestamp 1623621585
transform 1 0 22080 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_213
timestamp 1623621585
transform 1 0 20700 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_225
timestamp 1623621585
transform 1 0 21804 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_220
timestamp 1623621585
transform 1 0 21344 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_229
timestamp 1623621585
transform 1 0 22172 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_237
timestamp 1623621585
transform 1 0 22908 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_249
timestamp 1623621585
transform 1 0 24012 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_241
timestamp 1623621585
transform 1 0 23276 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1310
timestamp 1623621585
transform 1 0 24748 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_258
timestamp 1623621585
transform 1 0 24840 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_270
timestamp 1623621585
transform 1 0 25944 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_253
timestamp 1623621585
transform 1 0 24380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_265
timestamp 1623621585
transform 1 0 25484 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1317
timestamp 1623621585
transform 1 0 27324 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_282
timestamp 1623621585
transform 1 0 27048 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_277
timestamp 1623621585
transform 1 0 26588 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_286
timestamp 1623621585
transform 1 0 27416 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_294
timestamp 1623621585
transform 1 0 28152 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_306
timestamp 1623621585
transform 1 0 29256 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_298
timestamp 1623621585
transform 1 0 28520 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_310
timestamp 1623621585
transform 1 0 29624 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1311
timestamp 1623621585
transform 1 0 29992 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_315
timestamp 1623621585
transform 1 0 30084 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_327
timestamp 1623621585
transform 1 0 31188 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_322
timestamp 1623621585
transform 1 0 30728 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1318
timestamp 1623621585
transform 1 0 32568 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_339
timestamp 1623621585
transform 1 0 32292 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_351
timestamp 1623621585
transform 1 0 33396 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_334
timestamp 1623621585
transform 1 0 31832 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_126_343
timestamp 1623621585
transform 1 0 32660 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1312
timestamp 1623621585
transform 1 0 35236 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_363
timestamp 1623621585
transform 1 0 34500 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_125_372
timestamp 1623621585
transform 1 0 35328 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_355
timestamp 1623621585
transform 1 0 33764 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_367
timestamp 1623621585
transform 1 0 34868 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input261
timestamp 1623621585
transform 1 0 37076 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_384
timestamp 1623621585
transform 1 0 36432 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_379
timestamp 1623621585
transform 1 0 35972 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_395
timestamp 1623621585
transform 1 0 37444 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1623621585
transform -1 0 38824 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1623621585
transform -1 0 38824 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1319
timestamp 1623621585
transform 1 0 37812 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input260
timestamp 1623621585
transform 1 0 37812 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_125_396
timestamp 1623621585
transform 1 0 37536 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_403
timestamp 1623621585
transform 1 0 38180 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_400
timestamp 1623621585
transform 1 0 37904 0 -1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_406
timestamp 1623621585
transform 1 0 38456 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1623621585
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input409
timestamp 1623621585
transform 1 0 1748 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_127_3
timestamp 1623621585
transform 1 0 1380 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_127_11
timestamp 1623621585
transform 1 0 2116 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1320
timestamp 1623621585
transform 1 0 3772 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_127_23
timestamp 1623621585
transform 1 0 3220 0 1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_127_30
timestamp 1623621585
transform 1 0 3864 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_42
timestamp 1623621585
transform 1 0 4968 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_54
timestamp 1623621585
transform 1 0 6072 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_66
timestamp 1623621585
transform 1 0 7176 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_78
timestamp 1623621585
transform 1 0 8280 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1321
timestamp 1623621585
transform 1 0 9016 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_87
timestamp 1623621585
transform 1 0 9108 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_99
timestamp 1623621585
transform 1 0 10212 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_111
timestamp 1623621585
transform 1 0 11316 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_123
timestamp 1623621585
transform 1 0 12420 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1322
timestamp 1623621585
transform 1 0 14260 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_135
timestamp 1623621585
transform 1 0 13524 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_127_144
timestamp 1623621585
transform 1 0 14352 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_156
timestamp 1623621585
transform 1 0 15456 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_168
timestamp 1623621585
transform 1 0 16560 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_180
timestamp 1623621585
transform 1 0 17664 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1323
timestamp 1623621585
transform 1 0 19504 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_192
timestamp 1623621585
transform 1 0 18768 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_127_201
timestamp 1623621585
transform 1 0 19596 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_213
timestamp 1623621585
transform 1 0 20700 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_225
timestamp 1623621585
transform 1 0 21804 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_237
timestamp 1623621585
transform 1 0 22908 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_249
timestamp 1623621585
transform 1 0 24012 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1324
timestamp 1623621585
transform 1 0 24748 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_258
timestamp 1623621585
transform 1 0 24840 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_270
timestamp 1623621585
transform 1 0 25944 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_282
timestamp 1623621585
transform 1 0 27048 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_294
timestamp 1623621585
transform 1 0 28152 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_306
timestamp 1623621585
transform 1 0 29256 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1325
timestamp 1623621585
transform 1 0 29992 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_315
timestamp 1623621585
transform 1 0 30084 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_327
timestamp 1623621585
transform 1 0 31188 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_339
timestamp 1623621585
transform 1 0 32292 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_351
timestamp 1623621585
transform 1 0 33396 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0955_
timestamp 1623621585
transform 1 0 33764 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1326
timestamp 1623621585
transform 1 0 35236 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_359
timestamp 1623621585
transform 1 0 34132 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_372
timestamp 1623621585
transform 1 0 35328 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input263
timestamp 1623621585
transform 1 0 37076 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_127_384
timestamp 1623621585
transform 1 0 36432 0 1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_390
timestamp 1623621585
transform 1 0 36984 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_127_395
timestamp 1623621585
transform 1 0 37444 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1623621585
transform -1 0 38824 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input262
timestamp 1623621585
transform 1 0 37812 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_127_403
timestamp 1623621585
transform 1 0 38180 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1623621585
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1623621585
transform 1 0 1380 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1623621585
transform 1 0 2484 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_27
timestamp 1623621585
transform 1 0 3588 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_39
timestamp 1623621585
transform 1 0 4692 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1327
timestamp 1623621585
transform 1 0 6348 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_51
timestamp 1623621585
transform 1 0 5796 0 -1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_128_58
timestamp 1623621585
transform 1 0 6440 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_70
timestamp 1623621585
transform 1 0 7544 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_82
timestamp 1623621585
transform 1 0 8648 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_94
timestamp 1623621585
transform 1 0 9752 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1328
timestamp 1623621585
transform 1 0 11592 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_106
timestamp 1623621585
transform 1 0 10856 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_115
timestamp 1623621585
transform 1 0 11684 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_127
timestamp 1623621585
transform 1 0 12788 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_139
timestamp 1623621585
transform 1 0 13892 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_151
timestamp 1623621585
transform 1 0 14996 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_163
timestamp 1623621585
transform 1 0 16100 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1329
timestamp 1623621585
transform 1 0 16836 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_172
timestamp 1623621585
transform 1 0 16928 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_184
timestamp 1623621585
transform 1 0 18032 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_196
timestamp 1623621585
transform 1 0 19136 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_208
timestamp 1623621585
transform 1 0 20240 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1330
timestamp 1623621585
transform 1 0 22080 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_220
timestamp 1623621585
transform 1 0 21344 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_229
timestamp 1623621585
transform 1 0 22172 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_241
timestamp 1623621585
transform 1 0 23276 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_253
timestamp 1623621585
transform 1 0 24380 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_265
timestamp 1623621585
transform 1 0 25484 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1331
timestamp 1623621585
transform 1 0 27324 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_277
timestamp 1623621585
transform 1 0 26588 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_286
timestamp 1623621585
transform 1 0 27416 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_298
timestamp 1623621585
transform 1 0 28520 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_310
timestamp 1623621585
transform 1 0 29624 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_322
timestamp 1623621585
transform 1 0 30728 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1332
timestamp 1623621585
transform 1 0 32568 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_334
timestamp 1623621585
transform 1 0 31832 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_128_343
timestamp 1623621585
transform 1 0 32660 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_355
timestamp 1623621585
transform 1 0 33764 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_367
timestamp 1623621585
transform 1 0 34868 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input264
timestamp 1623621585
transform 1 0 37076 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_128_379
timestamp 1623621585
transform 1 0 35972 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_128_395
timestamp 1623621585
transform 1 0 37444 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1623621585
transform -1 0 38824 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1333
timestamp 1623621585
transform 1 0 37812 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_128_400
timestamp 1623621585
transform 1 0 37904 0 -1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_406
timestamp 1623621585
transform 1 0 38456 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1623621585
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input410
timestamp 1623621585
transform 1 0 1748 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_3
timestamp 1623621585
transform 1 0 1380 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_129_11
timestamp 1623621585
transform 1 0 2116 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1334
timestamp 1623621585
transform 1 0 3772 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_129_23
timestamp 1623621585
transform 1 0 3220 0 1 72352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_129_30
timestamp 1623621585
transform 1 0 3864 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_42
timestamp 1623621585
transform 1 0 4968 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_54
timestamp 1623621585
transform 1 0 6072 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_66
timestamp 1623621585
transform 1 0 7176 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_78
timestamp 1623621585
transform 1 0 8280 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1335
timestamp 1623621585
transform 1 0 9016 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_87
timestamp 1623621585
transform 1 0 9108 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_99
timestamp 1623621585
transform 1 0 10212 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_111
timestamp 1623621585
transform 1 0 11316 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_123
timestamp 1623621585
transform 1 0 12420 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1336
timestamp 1623621585
transform 1 0 14260 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_135
timestamp 1623621585
transform 1 0 13524 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_144
timestamp 1623621585
transform 1 0 14352 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_156
timestamp 1623621585
transform 1 0 15456 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_168
timestamp 1623621585
transform 1 0 16560 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_180
timestamp 1623621585
transform 1 0 17664 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1337
timestamp 1623621585
transform 1 0 19504 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_192
timestamp 1623621585
transform 1 0 18768 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_201
timestamp 1623621585
transform 1 0 19596 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_213
timestamp 1623621585
transform 1 0 20700 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_225
timestamp 1623621585
transform 1 0 21804 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_237
timestamp 1623621585
transform 1 0 22908 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_249
timestamp 1623621585
transform 1 0 24012 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1338
timestamp 1623621585
transform 1 0 24748 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_258
timestamp 1623621585
transform 1 0 24840 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_270
timestamp 1623621585
transform 1 0 25944 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_282
timestamp 1623621585
transform 1 0 27048 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_294
timestamp 1623621585
transform 1 0 28152 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_306
timestamp 1623621585
transform 1 0 29256 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1339
timestamp 1623621585
transform 1 0 29992 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_315
timestamp 1623621585
transform 1 0 30084 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_327
timestamp 1623621585
transform 1 0 31188 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_339
timestamp 1623621585
transform 1 0 32292 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_351
timestamp 1623621585
transform 1 0 33396 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1340
timestamp 1623621585
transform 1 0 35236 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_363
timestamp 1623621585
transform 1 0 34500 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_129_372
timestamp 1623621585
transform 1 0 35328 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_384
timestamp 1623621585
transform 1 0 36432 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1623621585
transform -1 0 38824 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input265
timestamp 1623621585
transform 1 0 37812 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_129_396
timestamp 1623621585
transform 1 0 37536 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_403
timestamp 1623621585
transform 1 0 38180 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1623621585
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input411
timestamp 1623621585
transform 1 0 1748 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_130_3
timestamp 1623621585
transform 1 0 1380 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_11
timestamp 1623621585
transform 1 0 2116 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_23
timestamp 1623621585
transform 1 0 3220 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_35
timestamp 1623621585
transform 1 0 4324 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1341
timestamp 1623621585
transform 1 0 6348 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_47
timestamp 1623621585
transform 1 0 5428 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_130_55
timestamp 1623621585
transform 1 0 6164 0 -1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_130_58
timestamp 1623621585
transform 1 0 6440 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_70
timestamp 1623621585
transform 1 0 7544 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_82
timestamp 1623621585
transform 1 0 8648 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_94
timestamp 1623621585
transform 1 0 9752 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1342
timestamp 1623621585
transform 1 0 11592 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_106
timestamp 1623621585
transform 1 0 10856 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_115
timestamp 1623621585
transform 1 0 11684 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_127
timestamp 1623621585
transform 1 0 12788 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_139
timestamp 1623621585
transform 1 0 13892 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_151
timestamp 1623621585
transform 1 0 14996 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_163
timestamp 1623621585
transform 1 0 16100 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1343
timestamp 1623621585
transform 1 0 16836 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_172
timestamp 1623621585
transform 1 0 16928 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_184
timestamp 1623621585
transform 1 0 18032 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_196
timestamp 1623621585
transform 1 0 19136 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_208
timestamp 1623621585
transform 1 0 20240 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1344
timestamp 1623621585
transform 1 0 22080 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_220
timestamp 1623621585
transform 1 0 21344 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_229
timestamp 1623621585
transform 1 0 22172 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_241
timestamp 1623621585
transform 1 0 23276 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_253
timestamp 1623621585
transform 1 0 24380 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_265
timestamp 1623621585
transform 1 0 25484 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1345
timestamp 1623621585
transform 1 0 27324 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_277
timestamp 1623621585
transform 1 0 26588 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_286
timestamp 1623621585
transform 1 0 27416 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_298
timestamp 1623621585
transform 1 0 28520 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_310
timestamp 1623621585
transform 1 0 29624 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_322
timestamp 1623621585
transform 1 0 30728 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1346
timestamp 1623621585
transform 1 0 32568 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_334
timestamp 1623621585
transform 1 0 31832 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_130_343
timestamp 1623621585
transform 1 0 32660 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_355
timestamp 1623621585
transform 1 0 33764 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_367
timestamp 1623621585
transform 1 0 34868 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input266
timestamp 1623621585
transform 1 0 37076 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_379
timestamp 1623621585
transform 1 0 35972 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_130_395
timestamp 1623621585
transform 1 0 37444 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1623621585
transform -1 0 38824 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1347
timestamp 1623621585
transform 1 0 37812 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_400
timestamp 1623621585
transform 1 0 37904 0 -1 73440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_406
timestamp 1623621585
transform 1 0 38456 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1623621585
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1623621585
transform 1 0 1380 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1623621585
transform 1 0 2484 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1348
timestamp 1623621585
transform 1 0 3772 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_131_27
timestamp 1623621585
transform 1 0 3588 0 1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_30
timestamp 1623621585
transform 1 0 3864 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_42
timestamp 1623621585
transform 1 0 4968 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_54
timestamp 1623621585
transform 1 0 6072 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_66
timestamp 1623621585
transform 1 0 7176 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_78
timestamp 1623621585
transform 1 0 8280 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1349
timestamp 1623621585
transform 1 0 9016 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_87
timestamp 1623621585
transform 1 0 9108 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_99
timestamp 1623621585
transform 1 0 10212 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_111
timestamp 1623621585
transform 1 0 11316 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_123
timestamp 1623621585
transform 1 0 12420 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1350
timestamp 1623621585
transform 1 0 14260 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_135
timestamp 1623621585
transform 1 0 13524 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_144
timestamp 1623621585
transform 1 0 14352 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_156
timestamp 1623621585
transform 1 0 15456 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_168
timestamp 1623621585
transform 1 0 16560 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_180
timestamp 1623621585
transform 1 0 17664 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1351
timestamp 1623621585
transform 1 0 19504 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_192
timestamp 1623621585
transform 1 0 18768 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_201
timestamp 1623621585
transform 1 0 19596 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_213
timestamp 1623621585
transform 1 0 20700 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_225
timestamp 1623621585
transform 1 0 21804 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_237
timestamp 1623621585
transform 1 0 22908 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_131_249
timestamp 1623621585
transform 1 0 24012 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1352
timestamp 1623621585
transform 1 0 24748 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_258
timestamp 1623621585
transform 1 0 24840 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_270
timestamp 1623621585
transform 1 0 25944 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_282
timestamp 1623621585
transform 1 0 27048 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0431_
timestamp 1623621585
transform 1 0 29164 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_131_294
timestamp 1623621585
transform 1 0 28152 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_131_302
timestamp 1623621585
transform 1 0 28888 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_309
timestamp 1623621585
transform 1 0 29532 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1353
timestamp 1623621585
transform 1 0 29992 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_131_313
timestamp 1623621585
transform 1 0 29900 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_315
timestamp 1623621585
transform 1 0 30084 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_327
timestamp 1623621585
transform 1 0 31188 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_339
timestamp 1623621585
transform 1 0 32292 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_351
timestamp 1623621585
transform 1 0 33396 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1354
timestamp 1623621585
transform 1 0 35236 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_363
timestamp 1623621585
transform 1 0 34500 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_372
timestamp 1623621585
transform 1 0 35328 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1623621585
transform 1 0 37076 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_131_384
timestamp 1623621585
transform 1 0 36432 0 1 73440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_390
timestamp 1623621585
transform 1 0 36984 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_395
timestamp 1623621585
transform 1 0 37444 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1623621585
transform -1 0 38824 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1623621585
transform 1 0 37812 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_403
timestamp 1623621585
transform 1 0 38180 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1623621585
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1623621585
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input412
timestamp 1623621585
transform 1 0 1748 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input413
timestamp 1623621585
transform 1 0 1748 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_132_3
timestamp 1623621585
transform 1 0 1380 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_11
timestamp 1623621585
transform 1 0 2116 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_3
timestamp 1623621585
transform 1 0 1380 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_11
timestamp 1623621585
transform 1 0 2116 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1362
timestamp 1623621585
transform 1 0 3772 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_23
timestamp 1623621585
transform 1 0 3220 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_35
timestamp 1623621585
transform 1 0 4324 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_23
timestamp 1623621585
transform 1 0 3220 0 1 74528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_30
timestamp 1623621585
transform 1 0 3864 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1355
timestamp 1623621585
transform 1 0 6348 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_47
timestamp 1623621585
transform 1 0 5428 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_132_55
timestamp 1623621585
transform 1 0 6164 0 -1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_132_58
timestamp 1623621585
transform 1 0 6440 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_42
timestamp 1623621585
transform 1 0 4968 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_54
timestamp 1623621585
transform 1 0 6072 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_70
timestamp 1623621585
transform 1 0 7544 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_82
timestamp 1623621585
transform 1 0 8648 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_66
timestamp 1623621585
transform 1 0 7176 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_78
timestamp 1623621585
transform 1 0 8280 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1363
timestamp 1623621585
transform 1 0 9016 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_94
timestamp 1623621585
transform 1 0 9752 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_87
timestamp 1623621585
transform 1 0 9108 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_99
timestamp 1623621585
transform 1 0 10212 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1356
timestamp 1623621585
transform 1 0 11592 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_106
timestamp 1623621585
transform 1 0 10856 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_115
timestamp 1623621585
transform 1 0 11684 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_111
timestamp 1623621585
transform 1 0 11316 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_123
timestamp 1623621585
transform 1 0 12420 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1364
timestamp 1623621585
transform 1 0 14260 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_127
timestamp 1623621585
transform 1 0 12788 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_139
timestamp 1623621585
transform 1 0 13892 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_135
timestamp 1623621585
transform 1 0 13524 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_144
timestamp 1623621585
transform 1 0 14352 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_151
timestamp 1623621585
transform 1 0 14996 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_163
timestamp 1623621585
transform 1 0 16100 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_156
timestamp 1623621585
transform 1 0 15456 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1357
timestamp 1623621585
transform 1 0 16836 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_172
timestamp 1623621585
transform 1 0 16928 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_184
timestamp 1623621585
transform 1 0 18032 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_168
timestamp 1623621585
transform 1 0 16560 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_180
timestamp 1623621585
transform 1 0 17664 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1365
timestamp 1623621585
transform 1 0 19504 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_196
timestamp 1623621585
transform 1 0 19136 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_208
timestamp 1623621585
transform 1 0 20240 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_192
timestamp 1623621585
transform 1 0 18768 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_201
timestamp 1623621585
transform 1 0 19596 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1358
timestamp 1623621585
transform 1 0 22080 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_220
timestamp 1623621585
transform 1 0 21344 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_229
timestamp 1623621585
transform 1 0 22172 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_213
timestamp 1623621585
transform 1 0 20700 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_225
timestamp 1623621585
transform 1 0 21804 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_241
timestamp 1623621585
transform 1 0 23276 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_237
timestamp 1623621585
transform 1 0 22908 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_249
timestamp 1623621585
transform 1 0 24012 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1366
timestamp 1623621585
transform 1 0 24748 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_253
timestamp 1623621585
transform 1 0 24380 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_265
timestamp 1623621585
transform 1 0 25484 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_258
timestamp 1623621585
transform 1 0 24840 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_270
timestamp 1623621585
transform 1 0 25944 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1359
timestamp 1623621585
transform 1 0 27324 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_277
timestamp 1623621585
transform 1 0 26588 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_286
timestamp 1623621585
transform 1 0 27416 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_282
timestamp 1623621585
transform 1 0 27048 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_298
timestamp 1623621585
transform 1 0 28520 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_310
timestamp 1623621585
transform 1 0 29624 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_294
timestamp 1623621585
transform 1 0 28152 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_306
timestamp 1623621585
transform 1 0 29256 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1367
timestamp 1623621585
transform 1 0 29992 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_322
timestamp 1623621585
transform 1 0 30728 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_315
timestamp 1623621585
transform 1 0 30084 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_327
timestamp 1623621585
transform 1 0 31188 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1360
timestamp 1623621585
transform 1 0 32568 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_334
timestamp 1623621585
transform 1 0 31832 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_343
timestamp 1623621585
transform 1 0 32660 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_339
timestamp 1623621585
transform 1 0 32292 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_351
timestamp 1623621585
transform 1 0 33396 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1368
timestamp 1623621585
transform 1 0 35236 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_355
timestamp 1623621585
transform 1 0 33764 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_367
timestamp 1623621585
transform 1 0 34868 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_363
timestamp 1623621585
transform 1 0 34500 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_372
timestamp 1623621585
transform 1 0 35328 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1623621585
transform 1 0 37076 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_379
timestamp 1623621585
transform 1 0 35972 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_132_395
timestamp 1623621585
transform 1 0 37444 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_133_384
timestamp 1623621585
transform 1 0 36432 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1623621585
transform -1 0 38824 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1623621585
transform -1 0 38824 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1361
timestamp 1623621585
transform 1 0 37812 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1623621585
transform 1 0 37812 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_132_400
timestamp 1623621585
transform 1 0 37904 0 -1 74528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_406
timestamp 1623621585
transform 1 0 38456 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_133_396
timestamp 1623621585
transform 1 0 37536 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_133_403
timestamp 1623621585
transform 1 0 38180 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1623621585
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1623621585
transform 1 0 1380 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1623621585
transform 1 0 2484 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_27
timestamp 1623621585
transform 1 0 3588 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_39
timestamp 1623621585
transform 1 0 4692 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1369
timestamp 1623621585
transform 1 0 6348 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_51
timestamp 1623621585
transform 1 0 5796 0 -1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_134_58
timestamp 1623621585
transform 1 0 6440 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_70
timestamp 1623621585
transform 1 0 7544 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_82
timestamp 1623621585
transform 1 0 8648 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_94
timestamp 1623621585
transform 1 0 9752 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1370
timestamp 1623621585
transform 1 0 11592 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_106
timestamp 1623621585
transform 1 0 10856 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_115
timestamp 1623621585
transform 1 0 11684 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_127
timestamp 1623621585
transform 1 0 12788 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_139
timestamp 1623621585
transform 1 0 13892 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_151
timestamp 1623621585
transform 1 0 14996 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_163
timestamp 1623621585
transform 1 0 16100 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1371
timestamp 1623621585
transform 1 0 16836 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_172
timestamp 1623621585
transform 1 0 16928 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_184
timestamp 1623621585
transform 1 0 18032 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_196
timestamp 1623621585
transform 1 0 19136 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_208
timestamp 1623621585
transform 1 0 20240 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1372
timestamp 1623621585
transform 1 0 22080 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_220
timestamp 1623621585
transform 1 0 21344 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_229
timestamp 1623621585
transform 1 0 22172 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_241
timestamp 1623621585
transform 1 0 23276 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_253
timestamp 1623621585
transform 1 0 24380 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_265
timestamp 1623621585
transform 1 0 25484 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1373
timestamp 1623621585
transform 1 0 27324 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_277
timestamp 1623621585
transform 1 0 26588 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_286
timestamp 1623621585
transform 1 0 27416 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_298
timestamp 1623621585
transform 1 0 28520 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_310
timestamp 1623621585
transform 1 0 29624 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_322
timestamp 1623621585
transform 1 0 30728 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1374
timestamp 1623621585
transform 1 0 32568 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_334
timestamp 1623621585
transform 1 0 31832 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_134_343
timestamp 1623621585
transform 1 0 32660 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_355
timestamp 1623621585
transform 1 0 33764 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_367
timestamp 1623621585
transform 1 0 34868 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1623621585
transform 1 0 37076 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_379
timestamp 1623621585
transform 1 0 35972 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_395
timestamp 1623621585
transform 1 0 37444 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1623621585
transform -1 0 38824 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1375
timestamp 1623621585
transform 1 0 37812 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_400
timestamp 1623621585
transform 1 0 37904 0 -1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_406
timestamp 1623621585
transform 1 0 38456 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1623621585
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input414
timestamp 1623621585
transform 1 0 1748 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_135_3
timestamp 1623621585
transform 1 0 1380 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_11
timestamp 1623621585
transform 1 0 2116 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1376
timestamp 1623621585
transform 1 0 3772 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_135_23
timestamp 1623621585
transform 1 0 3220 0 1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_135_30
timestamp 1623621585
transform 1 0 3864 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_42
timestamp 1623621585
transform 1 0 4968 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_54
timestamp 1623621585
transform 1 0 6072 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_66
timestamp 1623621585
transform 1 0 7176 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_78
timestamp 1623621585
transform 1 0 8280 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1377
timestamp 1623621585
transform 1 0 9016 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_87
timestamp 1623621585
transform 1 0 9108 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_99
timestamp 1623621585
transform 1 0 10212 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_111
timestamp 1623621585
transform 1 0 11316 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_123
timestamp 1623621585
transform 1 0 12420 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1378
timestamp 1623621585
transform 1 0 14260 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_135
timestamp 1623621585
transform 1 0 13524 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_135_144
timestamp 1623621585
transform 1 0 14352 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_156
timestamp 1623621585
transform 1 0 15456 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_168
timestamp 1623621585
transform 1 0 16560 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_180
timestamp 1623621585
transform 1 0 17664 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1379
timestamp 1623621585
transform 1 0 19504 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_192
timestamp 1623621585
transform 1 0 18768 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_135_201
timestamp 1623621585
transform 1 0 19596 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_213
timestamp 1623621585
transform 1 0 20700 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_225
timestamp 1623621585
transform 1 0 21804 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_237
timestamp 1623621585
transform 1 0 22908 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_249
timestamp 1623621585
transform 1 0 24012 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0735_
timestamp 1623621585
transform 1 0 25208 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1380
timestamp 1623621585
transform 1 0 24748 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_135_258
timestamp 1623621585
transform 1 0 24840 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_266
timestamp 1623621585
transform 1 0 25576 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_278
timestamp 1623621585
transform 1 0 26680 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_290
timestamp 1623621585
transform 1 0 27784 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_302
timestamp 1623621585
transform 1 0 28888 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1381
timestamp 1623621585
transform 1 0 29992 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_315
timestamp 1623621585
transform 1 0 30084 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_327
timestamp 1623621585
transform 1 0 31188 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_339
timestamp 1623621585
transform 1 0 32292 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_351
timestamp 1623621585
transform 1 0 33396 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1382
timestamp 1623621585
transform 1 0 35236 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_363
timestamp 1623621585
transform 1 0 34500 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_135_372
timestamp 1623621585
transform 1 0 35328 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input242
timestamp 1623621585
transform 1 0 37076 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_135_384
timestamp 1623621585
transform 1 0 36432 0 1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_390
timestamp 1623621585
transform 1 0 36984 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_135_395
timestamp 1623621585
transform 1 0 37444 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1623621585
transform -1 0 38824 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input241
timestamp 1623621585
transform 1 0 37812 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_135_403
timestamp 1623621585
transform 1 0 38180 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1623621585
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input415
timestamp 1623621585
transform 1 0 1380 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_6
timestamp 1623621585
transform 1 0 1656 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_18
timestamp 1623621585
transform 1 0 2760 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_30
timestamp 1623621585
transform 1 0 3864 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1383
timestamp 1623621585
transform 1 0 6348 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_42
timestamp 1623621585
transform 1 0 4968 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_136_54
timestamp 1623621585
transform 1 0 6072 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_58
timestamp 1623621585
transform 1 0 6440 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_70
timestamp 1623621585
transform 1 0 7544 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_82
timestamp 1623621585
transform 1 0 8648 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_94
timestamp 1623621585
transform 1 0 9752 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1384
timestamp 1623621585
transform 1 0 11592 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_106
timestamp 1623621585
transform 1 0 10856 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_115
timestamp 1623621585
transform 1 0 11684 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_127
timestamp 1623621585
transform 1 0 12788 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_139
timestamp 1623621585
transform 1 0 13892 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_151
timestamp 1623621585
transform 1 0 14996 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_163
timestamp 1623621585
transform 1 0 16100 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1385
timestamp 1623621585
transform 1 0 16836 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_172
timestamp 1623621585
transform 1 0 16928 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_184
timestamp 1623621585
transform 1 0 18032 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_196
timestamp 1623621585
transform 1 0 19136 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_208
timestamp 1623621585
transform 1 0 20240 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1386
timestamp 1623621585
transform 1 0 22080 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_220
timestamp 1623621585
transform 1 0 21344 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_229
timestamp 1623621585
transform 1 0 22172 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_241
timestamp 1623621585
transform 1 0 23276 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1623621585
transform 1 0 24748 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_253
timestamp 1623621585
transform 1 0 24380 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_136_261
timestamp 1623621585
transform 1 0 25116 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1387
timestamp 1623621585
transform 1 0 27324 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_273
timestamp 1623621585
transform 1 0 26220 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_286
timestamp 1623621585
transform 1 0 27416 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_298
timestamp 1623621585
transform 1 0 28520 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_310
timestamp 1623621585
transform 1 0 29624 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_322
timestamp 1623621585
transform 1 0 30728 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1388
timestamp 1623621585
transform 1 0 32568 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_334
timestamp 1623621585
transform 1 0 31832 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_136_343
timestamp 1623621585
transform 1 0 32660 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_355
timestamp 1623621585
transform 1 0 33764 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_367
timestamp 1623621585
transform 1 0 34868 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input243
timestamp 1623621585
transform 1 0 37076 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_136_379
timestamp 1623621585
transform 1 0 35972 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_395
timestamp 1623621585
transform 1 0 37444 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1623621585
transform -1 0 38824 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1389
timestamp 1623621585
transform 1 0 37812 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_136_400
timestamp 1623621585
transform 1 0 37904 0 -1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_406
timestamp 1623621585
transform 1 0 38456 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1623621585
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1623621585
transform 1 0 1380 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1623621585
transform 1 0 2484 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1390
timestamp 1623621585
transform 1 0 3772 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_137_27
timestamp 1623621585
transform 1 0 3588 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_30
timestamp 1623621585
transform 1 0 3864 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_42
timestamp 1623621585
transform 1 0 4968 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_54
timestamp 1623621585
transform 1 0 6072 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_66
timestamp 1623621585
transform 1 0 7176 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_78
timestamp 1623621585
transform 1 0 8280 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1391
timestamp 1623621585
transform 1 0 9016 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_87
timestamp 1623621585
transform 1 0 9108 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_99
timestamp 1623621585
transform 1 0 10212 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_111
timestamp 1623621585
transform 1 0 11316 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_123
timestamp 1623621585
transform 1 0 12420 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1392
timestamp 1623621585
transform 1 0 14260 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_135
timestamp 1623621585
transform 1 0 13524 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_144
timestamp 1623621585
transform 1 0 14352 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_156
timestamp 1623621585
transform 1 0 15456 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_168
timestamp 1623621585
transform 1 0 16560 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_180
timestamp 1623621585
transform 1 0 17664 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1393
timestamp 1623621585
transform 1 0 19504 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_192
timestamp 1623621585
transform 1 0 18768 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_201
timestamp 1623621585
transform 1 0 19596 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_213
timestamp 1623621585
transform 1 0 20700 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_225
timestamp 1623621585
transform 1 0 21804 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_237
timestamp 1623621585
transform 1 0 22908 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_249
timestamp 1623621585
transform 1 0 24012 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0410_
timestamp 1623621585
transform 1 0 25208 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1394
timestamp 1623621585
transform 1 0 24748 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_258
timestamp 1623621585
transform 1 0 24840 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_266
timestamp 1623621585
transform 1 0 25576 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_278
timestamp 1623621585
transform 1 0 26680 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_290
timestamp 1623621585
transform 1 0 27784 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0706_
timestamp 1623621585
transform 1 0 28980 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_302
timestamp 1623621585
transform 1 0 28888 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_137_307
timestamp 1623621585
transform 1 0 29348 0 1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1395
timestamp 1623621585
transform 1 0 29992 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_137_313
timestamp 1623621585
transform 1 0 29900 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_315
timestamp 1623621585
transform 1 0 30084 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_327
timestamp 1623621585
transform 1 0 31188 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_339
timestamp 1623621585
transform 1 0 32292 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_351
timestamp 1623621585
transform 1 0 33396 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1396
timestamp 1623621585
transform 1 0 35236 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_363
timestamp 1623621585
transform 1 0 34500 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_137_372
timestamp 1623621585
transform 1 0 35328 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_384
timestamp 1623621585
transform 1 0 36432 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1623621585
transform -1 0 38824 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input244
timestamp 1623621585
transform 1 0 37812 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_137_396
timestamp 1623621585
transform 1 0 37536 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_403
timestamp 1623621585
transform 1 0 38180 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1623621585
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_278
timestamp 1623621585
transform 1 0 1104 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input416
timestamp 1623621585
transform 1 0 1380 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input418
timestamp 1623621585
transform 1 0 1748 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_6
timestamp 1623621585
transform 1 0 1656 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_18
timestamp 1623621585
transform 1 0 2760 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_3
timestamp 1623621585
transform 1 0 1380 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_139_11
timestamp 1623621585
transform 1 0 2116 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1404
timestamp 1623621585
transform 1 0 3772 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_30
timestamp 1623621585
transform 1 0 3864 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_23
timestamp 1623621585
transform 1 0 3220 0 1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_139_30
timestamp 1623621585
transform 1 0 3864 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1397
timestamp 1623621585
transform 1 0 6348 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_42
timestamp 1623621585
transform 1 0 4968 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_54
timestamp 1623621585
transform 1 0 6072 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_58
timestamp 1623621585
transform 1 0 6440 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_42
timestamp 1623621585
transform 1 0 4968 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_54
timestamp 1623621585
transform 1 0 6072 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_70
timestamp 1623621585
transform 1 0 7544 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_82
timestamp 1623621585
transform 1 0 8648 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_66
timestamp 1623621585
transform 1 0 7176 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_78
timestamp 1623621585
transform 1 0 8280 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1405
timestamp 1623621585
transform 1 0 9016 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_94
timestamp 1623621585
transform 1 0 9752 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_87
timestamp 1623621585
transform 1 0 9108 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_99
timestamp 1623621585
transform 1 0 10212 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1398
timestamp 1623621585
transform 1 0 11592 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_106
timestamp 1623621585
transform 1 0 10856 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_115
timestamp 1623621585
transform 1 0 11684 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_111
timestamp 1623621585
transform 1 0 11316 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_123
timestamp 1623621585
transform 1 0 12420 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1406
timestamp 1623621585
transform 1 0 14260 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_127
timestamp 1623621585
transform 1 0 12788 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_139
timestamp 1623621585
transform 1 0 13892 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_135
timestamp 1623621585
transform 1 0 13524 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_144
timestamp 1623621585
transform 1 0 14352 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_151
timestamp 1623621585
transform 1 0 14996 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_163
timestamp 1623621585
transform 1 0 16100 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_156
timestamp 1623621585
transform 1 0 15456 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1399
timestamp 1623621585
transform 1 0 16836 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_172
timestamp 1623621585
transform 1 0 16928 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_184
timestamp 1623621585
transform 1 0 18032 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_168
timestamp 1623621585
transform 1 0 16560 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_180
timestamp 1623621585
transform 1 0 17664 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1407
timestamp 1623621585
transform 1 0 19504 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_196
timestamp 1623621585
transform 1 0 19136 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_208
timestamp 1623621585
transform 1 0 20240 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_192
timestamp 1623621585
transform 1 0 18768 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_201
timestamp 1623621585
transform 1 0 19596 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1400
timestamp 1623621585
transform 1 0 22080 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_220
timestamp 1623621585
transform 1 0 21344 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_229
timestamp 1623621585
transform 1 0 22172 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_213
timestamp 1623621585
transform 1 0 20700 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_225
timestamp 1623621585
transform 1 0 21804 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_241
timestamp 1623621585
transform 1 0 23276 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_237
timestamp 1623621585
transform 1 0 22908 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_249
timestamp 1623621585
transform 1 0 24012 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1408
timestamp 1623621585
transform 1 0 24748 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_253
timestamp 1623621585
transform 1 0 24380 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_265
timestamp 1623621585
transform 1 0 25484 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_258
timestamp 1623621585
transform 1 0 24840 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_270
timestamp 1623621585
transform 1 0 25944 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1401
timestamp 1623621585
transform 1 0 27324 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_277
timestamp 1623621585
transform 1 0 26588 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_286
timestamp 1623621585
transform 1 0 27416 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_282
timestamp 1623621585
transform 1 0 27048 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_139_290
timestamp 1623621585
transform 1 0 27784 0 1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  _0411_
timestamp 1623621585
transform 1 0 27968 0 1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0485_
timestamp 1623621585
transform 1 0 29164 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_298
timestamp 1623621585
transform 1 0 28520 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_310
timestamp 1623621585
transform 1 0 29624 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_298
timestamp 1623621585
transform 1 0 28520 0 1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_304
timestamp 1623621585
transform 1 0 29072 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_139_309
timestamp 1623621585
transform 1 0 29532 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1409
timestamp 1623621585
transform 1 0 29992 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_322
timestamp 1623621585
transform 1 0 30728 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_139_313
timestamp 1623621585
transform 1 0 29900 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_139_315
timestamp 1623621585
transform 1 0 30084 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_327
timestamp 1623621585
transform 1 0 31188 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1402
timestamp 1623621585
transform 1 0 32568 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_334
timestamp 1623621585
transform 1 0 31832 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_138_343
timestamp 1623621585
transform 1 0 32660 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_339
timestamp 1623621585
transform 1 0 32292 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_139_351
timestamp 1623621585
transform 1 0 33396 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1410
timestamp 1623621585
transform 1 0 35236 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_355
timestamp 1623621585
transform 1 0 33764 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_367
timestamp 1623621585
transform 1 0 34868 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_363
timestamp 1623621585
transform 1 0 34500 0 1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_139_372
timestamp 1623621585
transform 1 0 35328 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input245
timestamp 1623621585
transform 1 0 37076 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input248
timestamp 1623621585
transform 1 0 37076 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_379
timestamp 1623621585
transform 1 0 35972 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_395
timestamp 1623621585
transform 1 0 37444 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_139_384
timestamp 1623621585
transform 1 0 36432 0 1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_390
timestamp 1623621585
transform 1 0 36984 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_139_395
timestamp 1623621585
transform 1 0 37444 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1623621585
transform -1 0 38824 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_279
timestamp 1623621585
transform -1 0 38824 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1403
timestamp 1623621585
transform 1 0 37812 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input247
timestamp 1623621585
transform 1 0 37812 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_138_400
timestamp 1623621585
transform 1 0 37904 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_406
timestamp 1623621585
transform 1 0 38456 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_139_403
timestamp 1623621585
transform 1 0 38180 0 1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_280
timestamp 1623621585
transform 1 0 1104 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_140_3
timestamp 1623621585
transform 1 0 1380 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_15
timestamp 1623621585
transform 1 0 2484 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_27
timestamp 1623621585
transform 1 0 3588 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_39
timestamp 1623621585
transform 1 0 4692 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1411
timestamp 1623621585
transform 1 0 6348 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_140_51
timestamp 1623621585
transform 1 0 5796 0 -1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_140_58
timestamp 1623621585
transform 1 0 6440 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_70
timestamp 1623621585
transform 1 0 7544 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_82
timestamp 1623621585
transform 1 0 8648 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_94
timestamp 1623621585
transform 1 0 9752 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1412
timestamp 1623621585
transform 1 0 11592 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_106
timestamp 1623621585
transform 1 0 10856 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_140_115
timestamp 1623621585
transform 1 0 11684 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_127
timestamp 1623621585
transform 1 0 12788 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_139
timestamp 1623621585
transform 1 0 13892 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_151
timestamp 1623621585
transform 1 0 14996 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_163
timestamp 1623621585
transform 1 0 16100 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1413
timestamp 1623621585
transform 1 0 16836 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_172
timestamp 1623621585
transform 1 0 16928 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_184
timestamp 1623621585
transform 1 0 18032 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_196
timestamp 1623621585
transform 1 0 19136 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_208
timestamp 1623621585
transform 1 0 20240 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1414
timestamp 1623621585
transform 1 0 22080 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_220
timestamp 1623621585
transform 1 0 21344 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_140_229
timestamp 1623621585
transform 1 0 22172 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_241
timestamp 1623621585
transform 1 0 23276 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_253
timestamp 1623621585
transform 1 0 24380 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_265
timestamp 1623621585
transform 1 0 25484 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0769_
timestamp 1623621585
transform 1 0 27784 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1415
timestamp 1623621585
transform 1 0 27324 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_140_277
timestamp 1623621585
transform 1 0 26588 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_140_286
timestamp 1623621585
transform 1 0 27416 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0652_
timestamp 1623621585
transform 1 0 29164 0 -1 78880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_140_298
timestamp 1623621585
transform 1 0 28520 0 -1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_304
timestamp 1623621585
transform 1 0 29072 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_140_315
timestamp 1623621585
transform 1 0 30084 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_327
timestamp 1623621585
transform 1 0 31188 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1416
timestamp 1623621585
transform 1 0 32568 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_140_339
timestamp 1623621585
transform 1 0 32292 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_140_343
timestamp 1623621585
transform 1 0 32660 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_355
timestamp 1623621585
transform 1 0 33764 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_140_367
timestamp 1623621585
transform 1 0 34868 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input249
timestamp 1623621585
transform 1 0 37076 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_140_379
timestamp 1623621585
transform 1 0 35972 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_140_395
timestamp 1623621585
transform 1 0 37444 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_281
timestamp 1623621585
transform -1 0 38824 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1417
timestamp 1623621585
transform 1 0 37812 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_140_400
timestamp 1623621585
transform 1 0 37904 0 -1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_406
timestamp 1623621585
transform 1 0 38456 0 -1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_282
timestamp 1623621585
transform 1 0 1104 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input419
timestamp 1623621585
transform 1 0 1748 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_141_3
timestamp 1623621585
transform 1 0 1380 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_141_11
timestamp 1623621585
transform 1 0 2116 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1418
timestamp 1623621585
transform 1 0 3772 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_141_23
timestamp 1623621585
transform 1 0 3220 0 1 78880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_141_30
timestamp 1623621585
transform 1 0 3864 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_42
timestamp 1623621585
transform 1 0 4968 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_54
timestamp 1623621585
transform 1 0 6072 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_66
timestamp 1623621585
transform 1 0 7176 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_78
timestamp 1623621585
transform 1 0 8280 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1419
timestamp 1623621585
transform 1 0 9016 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_87
timestamp 1623621585
transform 1 0 9108 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_99
timestamp 1623621585
transform 1 0 10212 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_111
timestamp 1623621585
transform 1 0 11316 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_123
timestamp 1623621585
transform 1 0 12420 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1420
timestamp 1623621585
transform 1 0 14260 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_135
timestamp 1623621585
transform 1 0 13524 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_144
timestamp 1623621585
transform 1 0 14352 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_156
timestamp 1623621585
transform 1 0 15456 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_168
timestamp 1623621585
transform 1 0 16560 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_180
timestamp 1623621585
transform 1 0 17664 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1421
timestamp 1623621585
transform 1 0 19504 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_192
timestamp 1623621585
transform 1 0 18768 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_201
timestamp 1623621585
transform 1 0 19596 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_213
timestamp 1623621585
transform 1 0 20700 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_225
timestamp 1623621585
transform 1 0 21804 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_237
timestamp 1623621585
transform 1 0 22908 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_141_249
timestamp 1623621585
transform 1 0 24012 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1422
timestamp 1623621585
transform 1 0 24748 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_258
timestamp 1623621585
transform 1 0 24840 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_270
timestamp 1623621585
transform 1 0 25944 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0745_
timestamp 1623621585
transform 1 0 27048 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_141_290
timestamp 1623621585
transform 1 0 27784 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0598_
timestamp 1623621585
transform 1 0 29256 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0761_
timestamp 1623621585
transform 1 0 28152 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_141_302
timestamp 1623621585
transform 1 0 28888 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_141_310
timestamp 1623621585
transform 1 0 29624 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1423
timestamp 1623621585
transform 1 0 29992 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_141_315
timestamp 1623621585
transform 1 0 30084 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_327
timestamp 1623621585
transform 1 0 31188 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_339
timestamp 1623621585
transform 1 0 32292 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_351
timestamp 1623621585
transform 1 0 33396 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1424
timestamp 1623621585
transform 1 0 35236 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_141_363
timestamp 1623621585
transform 1 0 34500 0 1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_141_372
timestamp 1623621585
transform 1 0 35328 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_141_384
timestamp 1623621585
transform 1 0 36432 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_283
timestamp 1623621585
transform -1 0 38824 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input250
timestamp 1623621585
transform 1 0 37904 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_141_396
timestamp 1623621585
transform 1 0 37536 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_141_403
timestamp 1623621585
transform 1 0 38180 0 1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_284
timestamp 1623621585
transform 1 0 1104 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input427
timestamp 1623621585
transform 1 0 1380 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_6
timestamp 1623621585
transform 1 0 1656 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_18
timestamp 1623621585
transform 1 0 2760 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_30
timestamp 1623621585
transform 1 0 3864 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1425
timestamp 1623621585
transform 1 0 6348 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_42
timestamp 1623621585
transform 1 0 4968 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_142_54
timestamp 1623621585
transform 1 0 6072 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_58
timestamp 1623621585
transform 1 0 6440 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_70
timestamp 1623621585
transform 1 0 7544 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_82
timestamp 1623621585
transform 1 0 8648 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_94
timestamp 1623621585
transform 1 0 9752 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1426
timestamp 1623621585
transform 1 0 11592 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_106
timestamp 1623621585
transform 1 0 10856 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_115
timestamp 1623621585
transform 1 0 11684 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_127
timestamp 1623621585
transform 1 0 12788 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_139
timestamp 1623621585
transform 1 0 13892 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_151
timestamp 1623621585
transform 1 0 14996 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_163
timestamp 1623621585
transform 1 0 16100 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1427
timestamp 1623621585
transform 1 0 16836 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_172
timestamp 1623621585
transform 1 0 16928 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_184
timestamp 1623621585
transform 1 0 18032 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_196
timestamp 1623621585
transform 1 0 19136 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_208
timestamp 1623621585
transform 1 0 20240 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1428
timestamp 1623621585
transform 1 0 22080 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_142_220
timestamp 1623621585
transform 1 0 21344 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_142_229
timestamp 1623621585
transform 1 0 22172 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_241
timestamp 1623621585
transform 1 0 23276 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_253
timestamp 1623621585
transform 1 0 24380 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_265
timestamp 1623621585
transform 1 0 25484 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0737_
timestamp 1623621585
transform 1 0 27784 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0753_
timestamp 1623621585
transform 1 0 26220 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1429
timestamp 1623621585
transform 1 0 27324 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_281
timestamp 1623621585
transform 1 0 26956 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_142_286
timestamp 1623621585
transform 1 0 27416 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 29532 0 -1 79968
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_142_298
timestamp 1623621585
transform 1 0 28520 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_142_306
timestamp 1623621585
transform 1 0 29256 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_323
timestamp 1623621585
transform 1 0 30820 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1430
timestamp 1623621585
transform 1 0 32568 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_142_335
timestamp 1623621585
transform 1 0 31924 0 -1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_341
timestamp 1623621585
transform 1 0 32476 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_142_343
timestamp 1623621585
transform 1 0 32660 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_355
timestamp 1623621585
transform 1 0 33764 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_142_367
timestamp 1623621585
transform 1 0 34868 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input252
timestamp 1623621585
transform 1 0 37168 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_142_379
timestamp 1623621585
transform 1 0 35972 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_391
timestamp 1623621585
transform 1 0 37076 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_142_395
timestamp 1623621585
transform 1 0 37444 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_285
timestamp 1623621585
transform -1 0 38824 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1431
timestamp 1623621585
transform 1 0 37812 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_142_400
timestamp 1623621585
transform 1 0 37904 0 -1 79968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_406
timestamp 1623621585
transform 1 0 38456 0 -1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_286
timestamp 1623621585
transform 1 0 1104 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_143_3
timestamp 1623621585
transform 1 0 1380 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_15
timestamp 1623621585
transform 1 0 2484 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1432
timestamp 1623621585
transform 1 0 3772 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_143_27
timestamp 1623621585
transform 1 0 3588 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_143_30
timestamp 1623621585
transform 1 0 3864 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_42
timestamp 1623621585
transform 1 0 4968 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_54
timestamp 1623621585
transform 1 0 6072 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_66
timestamp 1623621585
transform 1 0 7176 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_78
timestamp 1623621585
transform 1 0 8280 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1433
timestamp 1623621585
transform 1 0 9016 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_87
timestamp 1623621585
transform 1 0 9108 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_99
timestamp 1623621585
transform 1 0 10212 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_111
timestamp 1623621585
transform 1 0 11316 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_123
timestamp 1623621585
transform 1 0 12420 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1434
timestamp 1623621585
transform 1 0 14260 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_135
timestamp 1623621585
transform 1 0 13524 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_143_144
timestamp 1623621585
transform 1 0 14352 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_156
timestamp 1623621585
transform 1 0 15456 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_168
timestamp 1623621585
transform 1 0 16560 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_180
timestamp 1623621585
transform 1 0 17664 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1435
timestamp 1623621585
transform 1 0 19504 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_192
timestamp 1623621585
transform 1 0 18768 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_143_201
timestamp 1623621585
transform 1 0 19596 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_213
timestamp 1623621585
transform 1 0 20700 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_225
timestamp 1623621585
transform 1 0 21804 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_237
timestamp 1623621585
transform 1 0 22908 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_143_249
timestamp 1623621585
transform 1 0 24012 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1436
timestamp 1623621585
transform 1 0 24748 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_258
timestamp 1623621585
transform 1 0 24840 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_270
timestamp 1623621585
transform 1 0 25944 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0720_
timestamp 1623621585
transform 1 0 27140 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_143_282
timestamp 1623621585
transform 1 0 27048 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_143_291
timestamp 1623621585
transform 1 0 27876 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0728_
timestamp 1623621585
transform 1 0 28244 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_143_303
timestamp 1623621585
transform 1 0 28980 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_143_311
timestamp 1623621585
transform 1 0 29716 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _0446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 31004 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1437
timestamp 1623621585
transform 1 0 29992 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_143_315
timestamp 1623621585
transform 1 0 30084 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_143_323
timestamp 1623621585
transform 1 0 30820 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_143_333
timestamp 1623621585
transform 1 0 31740 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_143_345
timestamp 1623621585
transform 1 0 32844 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1438
timestamp 1623621585
transform 1 0 35236 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_143_357
timestamp 1623621585
transform 1 0 33948 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_369
timestamp 1623621585
transform 1 0 35052 0 1 79968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_143_372
timestamp 1623621585
transform 1 0 35328 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input253
timestamp 1623621585
transform 1 0 37260 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_143_384
timestamp 1623621585
transform 1 0 36432 0 1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_143_392
timestamp 1623621585
transform 1 0 37168 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_287
timestamp 1623621585
transform -1 0 38824 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input251
timestamp 1623621585
transform 1 0 37904 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_143_396
timestamp 1623621585
transform 1 0 37536 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_143_403
timestamp 1623621585
transform 1 0 38180 0 1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_288
timestamp 1623621585
transform 1 0 1104 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input438
timestamp 1623621585
transform 1 0 1380 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_6
timestamp 1623621585
transform 1 0 1656 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_18
timestamp 1623621585
transform 1 0 2760 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_30
timestamp 1623621585
transform 1 0 3864 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1439
timestamp 1623621585
transform 1 0 6348 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_42
timestamp 1623621585
transform 1 0 4968 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_144_54
timestamp 1623621585
transform 1 0 6072 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_144_58
timestamp 1623621585
transform 1 0 6440 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_70
timestamp 1623621585
transform 1 0 7544 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_82
timestamp 1623621585
transform 1 0 8648 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_94
timestamp 1623621585
transform 1 0 9752 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1440
timestamp 1623621585
transform 1 0 11592 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_106
timestamp 1623621585
transform 1 0 10856 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_144_115
timestamp 1623621585
transform 1 0 11684 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_127
timestamp 1623621585
transform 1 0 12788 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_139
timestamp 1623621585
transform 1 0 13892 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_151
timestamp 1623621585
transform 1 0 14996 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_163
timestamp 1623621585
transform 1 0 16100 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1441
timestamp 1623621585
transform 1 0 16836 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_172
timestamp 1623621585
transform 1 0 16928 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_184
timestamp 1623621585
transform 1 0 18032 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_196
timestamp 1623621585
transform 1 0 19136 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_208
timestamp 1623621585
transform 1 0 20240 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1442
timestamp 1623621585
transform 1 0 22080 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_220
timestamp 1623621585
transform 1 0 21344 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_144_229
timestamp 1623621585
transform 1 0 22172 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_241
timestamp 1623621585
transform 1 0 23276 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_253
timestamp 1623621585
transform 1 0 24380 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_265
timestamp 1623621585
transform 1 0 25484 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0711_
timestamp 1623621585
transform 1 0 27784 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1443
timestamp 1623621585
transform 1 0 27324 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_144_277
timestamp 1623621585
transform 1 0 26588 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_144_286
timestamp 1623621585
transform 1 0 27416 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0738_
timestamp 1623621585
transform 1 0 29532 0 -1 81056
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_144_298
timestamp 1623621585
transform 1 0 28520 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_144_306
timestamp 1623621585
transform 1 0 29256 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _0437_
timestamp 1623621585
transform 1 0 31188 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_144_323
timestamp 1623621585
transform 1 0 30820 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1444
timestamp 1623621585
transform 1 0 32568 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_144_335
timestamp 1623621585
transform 1 0 31924 0 -1 81056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_341
timestamp 1623621585
transform 1 0 32476 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_144_343
timestamp 1623621585
transform 1 0 32660 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_355
timestamp 1623621585
transform 1 0 33764 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_367
timestamp 1623621585
transform 1 0 34868 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_144_379
timestamp 1623621585
transform 1 0 35972 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_391
timestamp 1623621585
transform 1 0 37076 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_289
timestamp 1623621585
transform -1 0 38824 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1445
timestamp 1623621585
transform 1 0 37812 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_144_400
timestamp 1623621585
transform 1 0 37904 0 -1 81056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_406
timestamp 1623621585
transform 1 0 38456 0 -1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_290
timestamp 1623621585
transform 1 0 1104 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_292
timestamp 1623621585
transform 1 0 1104 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input449
timestamp 1623621585
transform 1 0 1748 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_145_3
timestamp 1623621585
transform 1 0 1380 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_145_11
timestamp 1623621585
transform 1 0 2116 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_3
timestamp 1623621585
transform 1 0 1380 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_15
timestamp 1623621585
transform 1 0 2484 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1446
timestamp 1623621585
transform 1 0 3772 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_145_23
timestamp 1623621585
transform 1 0 3220 0 1 81056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_145_30
timestamp 1623621585
transform 1 0 3864 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_27
timestamp 1623621585
transform 1 0 3588 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_39
timestamp 1623621585
transform 1 0 4692 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1453
timestamp 1623621585
transform 1 0 6348 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_42
timestamp 1623621585
transform 1 0 4968 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_54
timestamp 1623621585
transform 1 0 6072 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_51
timestamp 1623621585
transform 1 0 5796 0 -1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_146_58
timestamp 1623621585
transform 1 0 6440 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_66
timestamp 1623621585
transform 1 0 7176 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_78
timestamp 1623621585
transform 1 0 8280 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_70
timestamp 1623621585
transform 1 0 7544 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_82
timestamp 1623621585
transform 1 0 8648 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1447
timestamp 1623621585
transform 1 0 9016 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_87
timestamp 1623621585
transform 1 0 9108 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_99
timestamp 1623621585
transform 1 0 10212 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_94
timestamp 1623621585
transform 1 0 9752 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1454
timestamp 1623621585
transform 1 0 11592 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_111
timestamp 1623621585
transform 1 0 11316 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_123
timestamp 1623621585
transform 1 0 12420 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_106
timestamp 1623621585
transform 1 0 10856 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_115
timestamp 1623621585
transform 1 0 11684 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1448
timestamp 1623621585
transform 1 0 14260 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_145_135
timestamp 1623621585
transform 1 0 13524 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_144
timestamp 1623621585
transform 1 0 14352 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_127
timestamp 1623621585
transform 1 0 12788 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_139
timestamp 1623621585
transform 1 0 13892 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_156
timestamp 1623621585
transform 1 0 15456 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_151
timestamp 1623621585
transform 1 0 14996 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_163
timestamp 1623621585
transform 1 0 16100 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1455
timestamp 1623621585
transform 1 0 16836 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_168
timestamp 1623621585
transform 1 0 16560 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_180
timestamp 1623621585
transform 1 0 17664 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_172
timestamp 1623621585
transform 1 0 16928 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_184
timestamp 1623621585
transform 1 0 18032 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1449
timestamp 1623621585
transform 1 0 19504 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_145_192
timestamp 1623621585
transform 1 0 18768 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_201
timestamp 1623621585
transform 1 0 19596 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_196
timestamp 1623621585
transform 1 0 19136 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_208
timestamp 1623621585
transform 1 0 20240 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1456
timestamp 1623621585
transform 1 0 22080 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_213
timestamp 1623621585
transform 1 0 20700 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_225
timestamp 1623621585
transform 1 0 21804 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_220
timestamp 1623621585
transform 1 0 21344 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_229
timestamp 1623621585
transform 1 0 22172 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_237
timestamp 1623621585
transform 1 0 22908 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_145_249
timestamp 1623621585
transform 1 0 24012 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_146_241
timestamp 1623621585
transform 1 0 23276 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1450
timestamp 1623621585
transform 1 0 24748 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_258
timestamp 1623621585
transform 1 0 24840 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_145_270
timestamp 1623621585
transform 1 0 25944 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_253
timestamp 1623621585
transform 1 0 24380 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_265
timestamp 1623621585
transform 1 0 25484 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1457
timestamp 1623621585
transform 1 0 27324 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_282
timestamp 1623621585
transform 1 0 27048 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_277
timestamp 1623621585
transform 1 0 26588 0 -1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_146_286
timestamp 1623621585
transform 1 0 27416 0 -1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _0712_
timestamp 1623621585
transform 1 0 29716 0 -1 82144
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0746_
timestamp 1623621585
transform 1 0 28336 0 1 81056
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0762_
timestamp 1623621585
transform 1 0 28060 0 -1 82144
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_145_294
timestamp 1623621585
transform 1 0 28152 0 1 81056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_145_310
timestamp 1623621585
transform 1 0 29624 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_292
timestamp 1623621585
transform 1 0 27968 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_307
timestamp 1623621585
transform 1 0 29348 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0729_
timestamp 1623621585
transform 1 0 30452 0 1 81056
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1451
timestamp 1623621585
transform 1 0 29992 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_145_315
timestamp 1623621585
transform 1 0 30084 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_145_333
timestamp 1623621585
transform 1 0 31740 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_146_325
timestamp 1623621585
transform 1 0 31004 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0754_
timestamp 1623621585
transform 1 0 32108 0 1 81056
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1458
timestamp 1623621585
transform 1 0 32568 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_145_351
timestamp 1623621585
transform 1 0 33396 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_146_337
timestamp 1623621585
transform 1 0 32108 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_146_341
timestamp 1623621585
transform 1 0 32476 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_343
timestamp 1623621585
transform 1 0 32660 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1452
timestamp 1623621585
transform 1 0 35236 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_145_363
timestamp 1623621585
transform 1 0 34500 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_145_372
timestamp 1623621585
transform 1 0 35328 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_355
timestamp 1623621585
transform 1 0 33764 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_146_367
timestamp 1623621585
transform 1 0 34868 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input255
timestamp 1623621585
transform 1 0 37260 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input258
timestamp 1623621585
transform 1 0 37168 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_145_384
timestamp 1623621585
transform 1 0 36432 0 1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_145_392
timestamp 1623621585
transform 1 0 37168 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_146_379
timestamp 1623621585
transform 1 0 35972 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_391
timestamp 1623621585
transform 1 0 37076 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_146_395
timestamp 1623621585
transform 1 0 37444 0 -1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_291
timestamp 1623621585
transform -1 0 38824 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_293
timestamp 1623621585
transform -1 0 38824 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1459
timestamp 1623621585
transform 1 0 37812 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input254
timestamp 1623621585
transform 1 0 37904 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_145_396
timestamp 1623621585
transform 1 0 37536 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_145_403
timestamp 1623621585
transform 1 0 38180 0 1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_146_400
timestamp 1623621585
transform 1 0 37904 0 -1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_406
timestamp 1623621585
transform 1 0 38456 0 -1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_294
timestamp 1623621585
transform 1 0 1104 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input452
timestamp 1623621585
transform 1 0 1748 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_147_3
timestamp 1623621585
transform 1 0 1380 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_147_11
timestamp 1623621585
transform 1 0 2116 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1460
timestamp 1623621585
transform 1 0 3772 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_147_23
timestamp 1623621585
transform 1 0 3220 0 1 82144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_147_30
timestamp 1623621585
transform 1 0 3864 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_42
timestamp 1623621585
transform 1 0 4968 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_54
timestamp 1623621585
transform 1 0 6072 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_66
timestamp 1623621585
transform 1 0 7176 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_78
timestamp 1623621585
transform 1 0 8280 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1461
timestamp 1623621585
transform 1 0 9016 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_87
timestamp 1623621585
transform 1 0 9108 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_99
timestamp 1623621585
transform 1 0 10212 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_111
timestamp 1623621585
transform 1 0 11316 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_123
timestamp 1623621585
transform 1 0 12420 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1462
timestamp 1623621585
transform 1 0 14260 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_135
timestamp 1623621585
transform 1 0 13524 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_147_144
timestamp 1623621585
transform 1 0 14352 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_156
timestamp 1623621585
transform 1 0 15456 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_168
timestamp 1623621585
transform 1 0 16560 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_180
timestamp 1623621585
transform 1 0 17664 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1463
timestamp 1623621585
transform 1 0 19504 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_147_192
timestamp 1623621585
transform 1 0 18768 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_147_201
timestamp 1623621585
transform 1 0 19596 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_213
timestamp 1623621585
transform 1 0 20700 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_225
timestamp 1623621585
transform 1 0 21804 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_237
timestamp 1623621585
transform 1 0 22908 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_147_249
timestamp 1623621585
transform 1 0 24012 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1464
timestamp 1623621585
transform 1 0 24748 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_258
timestamp 1623621585
transform 1 0 24840 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_270
timestamp 1623621585
transform 1 0 25944 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0683_
timestamp 1623621585
transform 1 0 27324 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_147_282
timestamp 1623621585
transform 1 0 27048 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0691_
timestamp 1623621585
transform 1 0 28428 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_147_293
timestamp 1623621585
transform 1 0 28060 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_147_305
timestamp 1623621585
transform 1 0 29164 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0721_
timestamp 1623621585
transform 1 0 30452 0 1 82144
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1465
timestamp 1623621585
transform 1 0 29992 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_147_313
timestamp 1623621585
transform 1 0 29900 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_147_315
timestamp 1623621585
transform 1 0 30084 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_147_333
timestamp 1623621585
transform 1 0 31740 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_147_345
timestamp 1623621585
transform 1 0 32844 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1466
timestamp 1623621585
transform 1 0 35236 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_147_357
timestamp 1623621585
transform 1 0 33948 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_369
timestamp 1623621585
transform 1 0 35052 0 1 82144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_147_372
timestamp 1623621585
transform 1 0 35328 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input259
timestamp 1623621585
transform 1 0 37260 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_147_384
timestamp 1623621585
transform 1 0 36432 0 1 82144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_147_392
timestamp 1623621585
transform 1 0 37168 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_295
timestamp 1623621585
transform -1 0 38824 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input256
timestamp 1623621585
transform 1 0 37904 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_147_396
timestamp 1623621585
transform 1 0 37536 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_147_403
timestamp 1623621585
transform 1 0 38180 0 1 82144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_296
timestamp 1623621585
transform 1 0 1104 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input453
timestamp 1623621585
transform 1 0 1380 0 -1 83232
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_148_13
timestamp 1623621585
transform 1 0 2300 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_25
timestamp 1623621585
transform 1 0 3404 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_37
timestamp 1623621585
transform 1 0 4508 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1467
timestamp 1623621585
transform 1 0 6348 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_49
timestamp 1623621585
transform 1 0 5612 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_58
timestamp 1623621585
transform 1 0 6440 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_70
timestamp 1623621585
transform 1 0 7544 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_82
timestamp 1623621585
transform 1 0 8648 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_94
timestamp 1623621585
transform 1 0 9752 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1468
timestamp 1623621585
transform 1 0 11592 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_106
timestamp 1623621585
transform 1 0 10856 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_115
timestamp 1623621585
transform 1 0 11684 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_127
timestamp 1623621585
transform 1 0 12788 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_139
timestamp 1623621585
transform 1 0 13892 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_151
timestamp 1623621585
transform 1 0 14996 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_163
timestamp 1623621585
transform 1 0 16100 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1469
timestamp 1623621585
transform 1 0 16836 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_148_172
timestamp 1623621585
transform 1 0 16928 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_184
timestamp 1623621585
transform 1 0 18032 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_196
timestamp 1623621585
transform 1 0 19136 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_208
timestamp 1623621585
transform 1 0 20240 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1470
timestamp 1623621585
transform 1 0 22080 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_220
timestamp 1623621585
transform 1 0 21344 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_148_229
timestamp 1623621585
transform 1 0 22172 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_241
timestamp 1623621585
transform 1 0 23276 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_253
timestamp 1623621585
transform 1 0 24380 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_265
timestamp 1623621585
transform 1 0 25484 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0674_
timestamp 1623621585
transform 1 0 27784 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1471
timestamp 1623621585
transform 1 0 27324 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_148_277
timestamp 1623621585
transform 1 0 26588 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_148_286
timestamp 1623621585
transform 1 0 27416 0 -1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_148_298
timestamp 1623621585
transform 1 0 28520 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_148_310
timestamp 1623621585
transform 1 0 29624 0 -1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0692_
timestamp 1623621585
transform 1 0 29992 0 -1 83232
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_148_328
timestamp 1623621585
transform 1 0 31280 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1472
timestamp 1623621585
transform 1 0 32568 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_148_340
timestamp 1623621585
transform 1 0 32384 0 -1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_148_343
timestamp 1623621585
transform 1 0 32660 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_355
timestamp 1623621585
transform 1 0 33764 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_367
timestamp 1623621585
transform 1 0 34868 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_148_379
timestamp 1623621585
transform 1 0 35972 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_391
timestamp 1623621585
transform 1 0 37076 0 -1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_297
timestamp 1623621585
transform -1 0 38824 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1473
timestamp 1623621585
transform 1 0 37812 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_148_400
timestamp 1623621585
transform 1 0 37904 0 -1 83232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_406
timestamp 1623621585
transform 1 0 38456 0 -1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_298
timestamp 1623621585
transform 1 0 1104 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_149_3
timestamp 1623621585
transform 1 0 1380 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_15
timestamp 1623621585
transform 1 0 2484 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1474
timestamp 1623621585
transform 1 0 3772 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_149_27
timestamp 1623621585
transform 1 0 3588 0 1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_149_30
timestamp 1623621585
transform 1 0 3864 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_42
timestamp 1623621585
transform 1 0 4968 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_54
timestamp 1623621585
transform 1 0 6072 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_66
timestamp 1623621585
transform 1 0 7176 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_78
timestamp 1623621585
transform 1 0 8280 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1475
timestamp 1623621585
transform 1 0 9016 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_87
timestamp 1623621585
transform 1 0 9108 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_99
timestamp 1623621585
transform 1 0 10212 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_111
timestamp 1623621585
transform 1 0 11316 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_123
timestamp 1623621585
transform 1 0 12420 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1476
timestamp 1623621585
transform 1 0 14260 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_135
timestamp 1623621585
transform 1 0 13524 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_144
timestamp 1623621585
transform 1 0 14352 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_156
timestamp 1623621585
transform 1 0 15456 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_168
timestamp 1623621585
transform 1 0 16560 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_180
timestamp 1623621585
transform 1 0 17664 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1477
timestamp 1623621585
transform 1 0 19504 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_149_192
timestamp 1623621585
transform 1 0 18768 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_149_201
timestamp 1623621585
transform 1 0 19596 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_213
timestamp 1623621585
transform 1 0 20700 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_225
timestamp 1623621585
transform 1 0 21804 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_237
timestamp 1623621585
transform 1 0 22908 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_149_249
timestamp 1623621585
transform 1 0 24012 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1478
timestamp 1623621585
transform 1 0 24748 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_258
timestamp 1623621585
transform 1 0 24840 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_270
timestamp 1623621585
transform 1 0 25944 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0657_
timestamp 1623621585
transform 1 0 27508 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_149_282
timestamp 1623621585
transform 1 0 27048 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_286
timestamp 1623621585
transform 1 0 27416 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0627_
timestamp 1623621585
transform 1 0 29256 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_149_295
timestamp 1623621585
transform 1 0 28244 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_149_303
timestamp 1623621585
transform 1 0 28980 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_149_310
timestamp 1623621585
transform 1 0 29624 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0684_
timestamp 1623621585
transform 1 0 30452 0 1 83232
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1479
timestamp 1623621585
transform 1 0 29992 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_149_315
timestamp 1623621585
transform 1 0 30084 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_149_333
timestamp 1623621585
transform 1 0 31740 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_149_345
timestamp 1623621585
transform 1 0 32844 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1480
timestamp 1623621585
transform 1 0 35236 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_149_357
timestamp 1623621585
transform 1 0 33948 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_369
timestamp 1623621585
transform 1 0 35052 0 1 83232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_149_372
timestamp 1623621585
transform 1 0 35328 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input278
timestamp 1623621585
transform 1 0 37260 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_149_384
timestamp 1623621585
transform 1 0 36432 0 1 83232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_149_392
timestamp 1623621585
transform 1 0 37168 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_299
timestamp 1623621585
transform -1 0 38824 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input267
timestamp 1623621585
transform 1 0 37904 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_149_396
timestamp 1623621585
transform 1 0 37536 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_149_403
timestamp 1623621585
transform 1 0 38180 0 1 83232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_300
timestamp 1623621585
transform 1 0 1104 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input454
timestamp 1623621585
transform 1 0 1748 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_150_3
timestamp 1623621585
transform 1 0 1380 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_150_11
timestamp 1623621585
transform 1 0 2116 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_23
timestamp 1623621585
transform 1 0 3220 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_35
timestamp 1623621585
transform 1 0 4324 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1481
timestamp 1623621585
transform 1 0 6348 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_47
timestamp 1623621585
transform 1 0 5428 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_150_55
timestamp 1623621585
transform 1 0 6164 0 -1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_150_58
timestamp 1623621585
transform 1 0 6440 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_70
timestamp 1623621585
transform 1 0 7544 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_82
timestamp 1623621585
transform 1 0 8648 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_94
timestamp 1623621585
transform 1 0 9752 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1482
timestamp 1623621585
transform 1 0 11592 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_106
timestamp 1623621585
transform 1 0 10856 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_150_115
timestamp 1623621585
transform 1 0 11684 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_127
timestamp 1623621585
transform 1 0 12788 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_139
timestamp 1623621585
transform 1 0 13892 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_151
timestamp 1623621585
transform 1 0 14996 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_163
timestamp 1623621585
transform 1 0 16100 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1483
timestamp 1623621585
transform 1 0 16836 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_150_172
timestamp 1623621585
transform 1 0 16928 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_184
timestamp 1623621585
transform 1 0 18032 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_196
timestamp 1623621585
transform 1 0 19136 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_208
timestamp 1623621585
transform 1 0 20240 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1484
timestamp 1623621585
transform 1 0 22080 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_220
timestamp 1623621585
transform 1 0 21344 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_150_229
timestamp 1623621585
transform 1 0 22172 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_241
timestamp 1623621585
transform 1 0 23276 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_253
timestamp 1623621585
transform 1 0 24380 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_265
timestamp 1623621585
transform 1 0 25484 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0666_
timestamp 1623621585
transform 1 0 27784 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1485
timestamp 1623621585
transform 1 0 27324 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_150_277
timestamp 1623621585
transform 1 0 26588 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_150_286
timestamp 1623621585
transform 1 0 27416 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0544_
timestamp 1623621585
transform 1 0 28888 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0573_
timestamp 1623621585
transform 1 0 29624 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_150_298
timestamp 1623621585
transform 1 0 28520 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_150_305
timestamp 1623621585
transform 1 0 29164 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_150_309
timestamp 1623621585
transform 1 0 29532 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0667_
timestamp 1623621585
transform 1 0 30360 0 -1 84320
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_150_314
timestamp 1623621585
transform 1 0 29992 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_150_332
timestamp 1623621585
transform 1 0 31648 0 -1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1486
timestamp 1623621585
transform 1 0 32568 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_150_340
timestamp 1623621585
transform 1 0 32384 0 -1 84320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_150_343
timestamp 1623621585
transform 1 0 32660 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_355
timestamp 1623621585
transform 1 0 33764 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_150_367
timestamp 1623621585
transform 1 0 34868 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input292
timestamp 1623621585
transform 1 0 37168 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_150_379
timestamp 1623621585
transform 1 0 35972 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_391
timestamp 1623621585
transform 1 0 37076 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_150_395
timestamp 1623621585
transform 1 0 37444 0 -1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_301
timestamp 1623621585
transform -1 0 38824 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1487
timestamp 1623621585
transform 1 0 37812 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_150_400
timestamp 1623621585
transform 1 0 37904 0 -1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_406
timestamp 1623621585
transform 1 0 38456 0 -1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_302
timestamp 1623621585
transform 1 0 1104 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_304
timestamp 1623621585
transform 1 0 1104 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input455
timestamp 1623621585
transform 1 0 1748 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_3
timestamp 1623621585
transform 1 0 1380 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_151_11
timestamp 1623621585
transform 1 0 2116 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_3
timestamp 1623621585
transform 1 0 1380 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_15
timestamp 1623621585
transform 1 0 2484 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1488
timestamp 1623621585
transform 1 0 3772 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_23
timestamp 1623621585
transform 1 0 3220 0 1 84320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_151_30
timestamp 1623621585
transform 1 0 3864 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_27
timestamp 1623621585
transform 1 0 3588 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_39
timestamp 1623621585
transform 1 0 4692 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1495
timestamp 1623621585
transform 1 0 6348 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_42
timestamp 1623621585
transform 1 0 4968 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_54
timestamp 1623621585
transform 1 0 6072 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_51
timestamp 1623621585
transform 1 0 5796 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_152_58
timestamp 1623621585
transform 1 0 6440 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_66
timestamp 1623621585
transform 1 0 7176 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_78
timestamp 1623621585
transform 1 0 8280 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_70
timestamp 1623621585
transform 1 0 7544 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_82
timestamp 1623621585
transform 1 0 8648 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1489
timestamp 1623621585
transform 1 0 9016 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_87
timestamp 1623621585
transform 1 0 9108 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_99
timestamp 1623621585
transform 1 0 10212 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_94
timestamp 1623621585
transform 1 0 9752 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1496
timestamp 1623621585
transform 1 0 11592 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_111
timestamp 1623621585
transform 1 0 11316 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_123
timestamp 1623621585
transform 1 0 12420 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_106
timestamp 1623621585
transform 1 0 10856 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_152_115
timestamp 1623621585
transform 1 0 11684 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1490
timestamp 1623621585
transform 1 0 14260 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_135
timestamp 1623621585
transform 1 0 13524 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_144
timestamp 1623621585
transform 1 0 14352 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_127
timestamp 1623621585
transform 1 0 12788 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_139
timestamp 1623621585
transform 1 0 13892 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_156
timestamp 1623621585
transform 1 0 15456 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_151
timestamp 1623621585
transform 1 0 14996 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_163
timestamp 1623621585
transform 1 0 16100 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1497
timestamp 1623621585
transform 1 0 16836 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_168
timestamp 1623621585
transform 1 0 16560 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_180
timestamp 1623621585
transform 1 0 17664 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_172
timestamp 1623621585
transform 1 0 16928 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_184
timestamp 1623621585
transform 1 0 18032 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1491
timestamp 1623621585
transform 1 0 19504 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_192
timestamp 1623621585
transform 1 0 18768 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_201
timestamp 1623621585
transform 1 0 19596 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_196
timestamp 1623621585
transform 1 0 19136 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_208
timestamp 1623621585
transform 1 0 20240 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1498
timestamp 1623621585
transform 1 0 22080 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_213
timestamp 1623621585
transform 1 0 20700 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_225
timestamp 1623621585
transform 1 0 21804 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_220
timestamp 1623621585
transform 1 0 21344 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_152_229
timestamp 1623621585
transform 1 0 22172 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0707_
timestamp 1623621585
transform 1 0 23092 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_151_237
timestamp 1623621585
transform 1 0 22908 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_249
timestamp 1623621585
transform 1 0 24012 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_152_237
timestamp 1623621585
transform 1 0 22908 0 -1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_152_243
timestamp 1623621585
transform 1 0 23460 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1492
timestamp 1623621585
transform 1 0 24748 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_258
timestamp 1623621585
transform 1 0 24840 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_151_270
timestamp 1623621585
transform 1 0 25944 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_255
timestamp 1623621585
transform 1 0 24564 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_267
timestamp 1623621585
transform 1 0 25668 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0436_
timestamp 1623621585
transform 1 0 27784 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0545_
timestamp 1623621585
transform 1 0 26588 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0629_
timestamp 1623621585
transform 1 0 27784 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1499
timestamp 1623621585
transform 1 0 27324 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_282
timestamp 1623621585
transform 1 0 27048 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_152_275
timestamp 1623621585
transform 1 0 26404 0 -1 85408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_152_281
timestamp 1623621585
transform 1 0 26956 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_152_286
timestamp 1623621585
transform 1 0 27416 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0486_
timestamp 1623621585
transform 1 0 28888 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0637_
timestamp 1623621585
transform 1 0 28888 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_151_298
timestamp 1623621585
transform 1 0 28520 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_151_306
timestamp 1623621585
transform 1 0 29256 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_152_298
timestamp 1623621585
transform 1 0 28520 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_152_310
timestamp 1623621585
transform 1 0 29624 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0452_
timestamp 1623621585
transform 1 0 29992 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0638_
timestamp 1623621585
transform 1 0 30728 0 -1 85408
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0658_
timestamp 1623621585
transform 1 0 30452 0 1 84320
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1493
timestamp 1623621585
transform 1 0 29992 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_151_315
timestamp 1623621585
transform 1 0 30084 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_333
timestamp 1623621585
transform 1 0 31740 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_152_318
timestamp 1623621585
transform 1 0 30360 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0675_
timestamp 1623621585
transform 1 0 32108 0 1 84320
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1623621585
transform 1 0 33304 0 -1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1500
timestamp 1623621585
transform 1 0 32568 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_151_351
timestamp 1623621585
transform 1 0 33396 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_336
timestamp 1623621585
transform 1 0 32016 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_152_343
timestamp 1623621585
transform 1 0 32660 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_349
timestamp 1623621585
transform 1 0 33212 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_354
timestamp 1623621585
transform 1 0 33672 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1494
timestamp 1623621585
transform 1 0 35236 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_151_363
timestamp 1623621585
transform 1 0 34500 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_151_372
timestamp 1623621585
transform 1 0 35328 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_152_366
timestamp 1623621585
transform 1 0 34776 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input293
timestamp 1623621585
transform 1 0 37260 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_151_384
timestamp 1623621585
transform 1 0 36432 0 1 84320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_392
timestamp 1623621585
transform 1 0 37168 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_152_378
timestamp 1623621585
transform 1 0 35880 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_390
timestamp 1623621585
transform 1 0 36984 0 -1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_303
timestamp 1623621585
transform -1 0 38824 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_305
timestamp 1623621585
transform -1 0 38824 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1501
timestamp 1623621585
transform 1 0 37812 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input289
timestamp 1623621585
transform 1 0 37904 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_151_396
timestamp 1623621585
transform 1 0 37536 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_151_403
timestamp 1623621585
transform 1 0 38180 0 1 84320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_152_398
timestamp 1623621585
transform 1 0 37720 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_152_400
timestamp 1623621585
transform 1 0 37904 0 -1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_406
timestamp 1623621585
transform 1 0 38456 0 -1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_306
timestamp 1623621585
transform 1 0 1104 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input456
timestamp 1623621585
transform 1 0 1748 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_153_3
timestamp 1623621585
transform 1 0 1380 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_153_11
timestamp 1623621585
transform 1 0 2116 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1502
timestamp 1623621585
transform 1 0 3772 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_153_23
timestamp 1623621585
transform 1 0 3220 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_153_30
timestamp 1623621585
transform 1 0 3864 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_42
timestamp 1623621585
transform 1 0 4968 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_54
timestamp 1623621585
transform 1 0 6072 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_66
timestamp 1623621585
transform 1 0 7176 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_78
timestamp 1623621585
transform 1 0 8280 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1503
timestamp 1623621585
transform 1 0 9016 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_87
timestamp 1623621585
transform 1 0 9108 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_99
timestamp 1623621585
transform 1 0 10212 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_111
timestamp 1623621585
transform 1 0 11316 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_123
timestamp 1623621585
transform 1 0 12420 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1504
timestamp 1623621585
transform 1 0 14260 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_153_135
timestamp 1623621585
transform 1 0 13524 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_153_144
timestamp 1623621585
transform 1 0 14352 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_156
timestamp 1623621585
transform 1 0 15456 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_168
timestamp 1623621585
transform 1 0 16560 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_180
timestamp 1623621585
transform 1 0 17664 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1505
timestamp 1623621585
transform 1 0 19504 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_153_192
timestamp 1623621585
transform 1 0 18768 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_153_201
timestamp 1623621585
transform 1 0 19596 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_213
timestamp 1623621585
transform 1 0 20700 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_225
timestamp 1623621585
transform 1 0 21804 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_237
timestamp 1623621585
transform 1 0 22908 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_153_249
timestamp 1623621585
transform 1 0 24012 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1506
timestamp 1623621585
transform 1 0 24748 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_258
timestamp 1623621585
transform 1 0 24840 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_153_270
timestamp 1623621585
transform 1 0 25944 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0445_
timestamp 1623621585
transform 1 0 27784 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_153_282
timestamp 1623621585
transform 1 0 27048 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0620_
timestamp 1623621585
transform 1 0 28888 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_153_298
timestamp 1623621585
transform 1 0 28520 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_153_310
timestamp 1623621585
transform 1 0 29624 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0630_
timestamp 1623621585
transform 1 0 30728 0 1 85408
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1507
timestamp 1623621585
transform 1 0 29992 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_153_315
timestamp 1623621585
transform 1 0 30084 0 1 85408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_321
timestamp 1623621585
transform 1 0 30636 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0430_
timestamp 1623621585
transform 1 0 33488 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _0463_
timestamp 1623621585
transform 1 0 32384 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_153_336
timestamp 1623621585
transform 1 0 32016 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_153_348
timestamp 1623621585
transform 1 0 33120 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1508
timestamp 1623621585
transform 1 0 35236 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_153_356
timestamp 1623621585
transform 1 0 33856 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_153_368
timestamp 1623621585
transform 1 0 34960 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_153_372
timestamp 1623621585
transform 1 0 35328 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input295
timestamp 1623621585
transform 1 0 37260 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_153_384
timestamp 1623621585
transform 1 0 36432 0 1 85408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_153_392
timestamp 1623621585
transform 1 0 37168 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_307
timestamp 1623621585
transform -1 0 38824 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input294
timestamp 1623621585
transform 1 0 37904 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_153_396
timestamp 1623621585
transform 1 0 37536 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_153_403
timestamp 1623621585
transform 1 0 38180 0 1 85408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_308
timestamp 1623621585
transform 1 0 1104 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input457
timestamp 1623621585
transform 1 0 1748 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_154_3
timestamp 1623621585
transform 1 0 1380 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_154_11
timestamp 1623621585
transform 1 0 2116 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_23
timestamp 1623621585
transform 1 0 3220 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_35
timestamp 1623621585
transform 1 0 4324 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1509
timestamp 1623621585
transform 1 0 6348 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_47
timestamp 1623621585
transform 1 0 5428 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_55
timestamp 1623621585
transform 1 0 6164 0 -1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_154_58
timestamp 1623621585
transform 1 0 6440 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_70
timestamp 1623621585
transform 1 0 7544 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_82
timestamp 1623621585
transform 1 0 8648 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_94
timestamp 1623621585
transform 1 0 9752 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1510
timestamp 1623621585
transform 1 0 11592 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_106
timestamp 1623621585
transform 1 0 10856 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_154_115
timestamp 1623621585
transform 1 0 11684 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_127
timestamp 1623621585
transform 1 0 12788 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_139
timestamp 1623621585
transform 1 0 13892 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_151
timestamp 1623621585
transform 1 0 14996 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_163
timestamp 1623621585
transform 1 0 16100 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1511
timestamp 1623621585
transform 1 0 16836 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_172
timestamp 1623621585
transform 1 0 16928 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_184
timestamp 1623621585
transform 1 0 18032 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1623621585
transform 1 0 19872 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_196
timestamp 1623621585
transform 1 0 19136 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_154_207
timestamp 1623621585
transform 1 0 20148 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1512
timestamp 1623621585
transform 1 0 22080 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_219
timestamp 1623621585
transform 1 0 21252 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_227
timestamp 1623621585
transform 1 0 21988 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_229
timestamp 1623621585
transform 1 0 22172 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0432_
timestamp 1623621585
transform 1 0 23368 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_154_241
timestamp 1623621585
transform 1 0 23276 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_154_246
timestamp 1623621585
transform 1 0 23736 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_258
timestamp 1623621585
transform 1 0 24840 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_270
timestamp 1623621585
transform 1 0 25944 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0488_
timestamp 1623621585
transform 1 0 26588 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1513
timestamp 1623621585
transform 1 0 27324 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_154_276
timestamp 1623621585
transform 1 0 26496 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_154_281
timestamp 1623621585
transform 1 0 26956 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_154_286
timestamp 1623621585
transform 1 0 27416 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0583_
timestamp 1623621585
transform 1 0 27968 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0603_
timestamp 1623621585
transform 1 0 29072 0 -1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_154_300
timestamp 1623621585
transform 1 0 28704 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_154_312
timestamp 1623621585
transform 1 0 29808 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0519_
timestamp 1623621585
transform 1 0 30176 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0613_
timestamp 1623621585
transform 1 0 30912 0 -1 86496
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_154_320
timestamp 1623621585
transform 1 0 30544 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0543_
timestamp 1623621585
transform 1 0 33028 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1514
timestamp 1623621585
transform 1 0 32568 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_154_338
timestamp 1623621585
transform 1 0 32200 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_154_343
timestamp 1623621585
transform 1 0 32660 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_154_351
timestamp 1623621585
transform 1 0 33396 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_363
timestamp 1623621585
transform 1 0 34500 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_154_375
timestamp 1623621585
transform 1 0 35604 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input297
timestamp 1623621585
transform 1 0 37168 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_154_387
timestamp 1623621585
transform 1 0 36708 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_154_391
timestamp 1623621585
transform 1 0 37076 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_154_395
timestamp 1623621585
transform 1 0 37444 0 -1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_309
timestamp 1623621585
transform -1 0 38824 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1515
timestamp 1623621585
transform 1 0 37812 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_154_400
timestamp 1623621585
transform 1 0 37904 0 -1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_406
timestamp 1623621585
transform 1 0 38456 0 -1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_310
timestamp 1623621585
transform 1 0 1104 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_155_3
timestamp 1623621585
transform 1 0 1380 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_15
timestamp 1623621585
transform 1 0 2484 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1516
timestamp 1623621585
transform 1 0 3772 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_155_27
timestamp 1623621585
transform 1 0 3588 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_155_30
timestamp 1623621585
transform 1 0 3864 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_42
timestamp 1623621585
transform 1 0 4968 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_54
timestamp 1623621585
transform 1 0 6072 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_66
timestamp 1623621585
transform 1 0 7176 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_78
timestamp 1623621585
transform 1 0 8280 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1517
timestamp 1623621585
transform 1 0 9016 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_87
timestamp 1623621585
transform 1 0 9108 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_99
timestamp 1623621585
transform 1 0 10212 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_111
timestamp 1623621585
transform 1 0 11316 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_123
timestamp 1623621585
transform 1 0 12420 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1518
timestamp 1623621585
transform 1 0 14260 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_155_135
timestamp 1623621585
transform 1 0 13524 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_144
timestamp 1623621585
transform 1 0 14352 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_156
timestamp 1623621585
transform 1 0 15456 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_168
timestamp 1623621585
transform 1 0 16560 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_180
timestamp 1623621585
transform 1 0 17664 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1519
timestamp 1623621585
transform 1 0 19504 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_155_192
timestamp 1623621585
transform 1 0 18768 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_201
timestamp 1623621585
transform 1 0 19596 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_213
timestamp 1623621585
transform 1 0 20700 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_225
timestamp 1623621585
transform 1 0 21804 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0487_
timestamp 1623621585
transform 1 0 23828 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_4  _0799_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22448 0 1 86496
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_155_231
timestamp 1623621585
transform 1 0 22356 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_155_243
timestamp 1623621585
transform 1 0 23460 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1520
timestamp 1623621585
transform 1 0 24748 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_155_251
timestamp 1623621585
transform 1 0 24196 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_155_258
timestamp 1623621585
transform 1 0 24840 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_155_270
timestamp 1623621585
transform 1 0 25944 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0612_
timestamp 1623621585
transform 1 0 26864 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_155_278
timestamp 1623621585
transform 1 0 26680 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_155_288
timestamp 1623621585
transform 1 0 27600 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0462_
timestamp 1623621585
transform 1 0 27968 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_155_300
timestamp 1623621585
transform 1 0 28704 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_155_312
timestamp 1623621585
transform 1 0 29808 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0604_
timestamp 1623621585
transform 1 0 31004 0 1 86496
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1521
timestamp 1623621585
transform 1 0 29992 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_155_315
timestamp 1623621585
transform 1 0 30084 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_155_323
timestamp 1623621585
transform 1 0 30820 0 1 86496
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_2  _0455_
timestamp 1623621585
transform 1 0 32660 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_155_339
timestamp 1623621585
transform 1 0 32292 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_155_351
timestamp 1623621585
transform 1 0 33396 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1623621585
transform 1 0 33764 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1522
timestamp 1623621585
transform 1 0 35236 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_155_359
timestamp 1623621585
transform 1 0 34132 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_155_372
timestamp 1623621585
transform 1 0 35328 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input298
timestamp 1623621585
transform 1 0 37260 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_155_384
timestamp 1623621585
transform 1 0 36432 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_155_392
timestamp 1623621585
transform 1 0 37168 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_311
timestamp 1623621585
transform -1 0 38824 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input296
timestamp 1623621585
transform 1 0 37904 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_155_396
timestamp 1623621585
transform 1 0 37536 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_155_403
timestamp 1623621585
transform 1 0 38180 0 1 86496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_312
timestamp 1623621585
transform 1 0 1104 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input458
timestamp 1623621585
transform 1 0 1748 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_156_3
timestamp 1623621585
transform 1 0 1380 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_156_11
timestamp 1623621585
transform 1 0 2116 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_23
timestamp 1623621585
transform 1 0 3220 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_35
timestamp 1623621585
transform 1 0 4324 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1523
timestamp 1623621585
transform 1 0 6348 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_47
timestamp 1623621585
transform 1 0 5428 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_156_55
timestamp 1623621585
transform 1 0 6164 0 -1 87584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_156_58
timestamp 1623621585
transform 1 0 6440 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_70
timestamp 1623621585
transform 1 0 7544 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_82
timestamp 1623621585
transform 1 0 8648 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_94
timestamp 1623621585
transform 1 0 9752 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1524
timestamp 1623621585
transform 1 0 11592 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_106
timestamp 1623621585
transform 1 0 10856 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_156_115
timestamp 1623621585
transform 1 0 11684 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_127
timestamp 1623621585
transform 1 0 12788 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_139
timestamp 1623621585
transform 1 0 13892 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_151
timestamp 1623621585
transform 1 0 14996 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_163
timestamp 1623621585
transform 1 0 16100 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1525
timestamp 1623621585
transform 1 0 16836 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_156_172
timestamp 1623621585
transform 1 0 16928 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_184
timestamp 1623621585
transform 1 0 18032 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_196
timestamp 1623621585
transform 1 0 19136 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_208
timestamp 1623621585
transform 1 0 20240 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1526
timestamp 1623621585
transform 1 0 22080 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_156_220
timestamp 1623621585
transform 1 0 21344 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_156_229
timestamp 1623621585
transform 1 0 22172 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0653_
timestamp 1623621585
transform 1 0 23276 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_156_245
timestamp 1623621585
transform 1 0 23644 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_257
timestamp 1623621585
transform 1 0 24748 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_269
timestamp 1623621585
transform 1 0 25852 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1527
timestamp 1623621585
transform 1 0 27324 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_156_281
timestamp 1623621585
transform 1 0 26956 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_156_286
timestamp 1623621585
transform 1 0 27416 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0454_
timestamp 1623621585
transform 1 0 27968 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0621_
timestamp 1623621585
transform 1 0 29256 0 -1 87584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_156_300
timestamp 1623621585
transform 1 0 28704 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _0584_
timestamp 1623621585
transform 1 0 30912 0 -1 87584
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_156_320
timestamp 1623621585
transform 1 0 30544 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0484_
timestamp 1623621585
transform 1 0 33028 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1528
timestamp 1623621585
transform 1 0 32568 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_156_338
timestamp 1623621585
transform 1 0 32200 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_156_343
timestamp 1623621585
transform 1 0 32660 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_156_351
timestamp 1623621585
transform 1 0 33396 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_363
timestamp 1623621585
transform 1 0 34500 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_375
timestamp 1623621585
transform 1 0 35604 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_156_387
timestamp 1623621585
transform 1 0 36708 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_313
timestamp 1623621585
transform -1 0 38824 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1529
timestamp 1623621585
transform 1 0 37812 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_156_400
timestamp 1623621585
transform 1 0 37904 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_406
timestamp 1623621585
transform 1 0 38456 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_314
timestamp 1623621585
transform 1 0 1104 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input428
timestamp 1623621585
transform 1 0 1748 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_157_3
timestamp 1623621585
transform 1 0 1380 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_157_11
timestamp 1623621585
transform 1 0 2116 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1530
timestamp 1623621585
transform 1 0 3772 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_157_23
timestamp 1623621585
transform 1 0 3220 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_157_30
timestamp 1623621585
transform 1 0 3864 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_42
timestamp 1623621585
transform 1 0 4968 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_54
timestamp 1623621585
transform 1 0 6072 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_66
timestamp 1623621585
transform 1 0 7176 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_78
timestamp 1623621585
transform 1 0 8280 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1531
timestamp 1623621585
transform 1 0 9016 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_87
timestamp 1623621585
transform 1 0 9108 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_99
timestamp 1623621585
transform 1 0 10212 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_111
timestamp 1623621585
transform 1 0 11316 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_123
timestamp 1623621585
transform 1 0 12420 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1532
timestamp 1623621585
transform 1 0 14260 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_157_135
timestamp 1623621585
transform 1 0 13524 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_157_144
timestamp 1623621585
transform 1 0 14352 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_156
timestamp 1623621585
transform 1 0 15456 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_168
timestamp 1623621585
transform 1 0 16560 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_180
timestamp 1623621585
transform 1 0 17664 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1533
timestamp 1623621585
transform 1 0 19504 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_157_192
timestamp 1623621585
transform 1 0 18768 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_157_201
timestamp 1623621585
transform 1 0 19596 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_213
timestamp 1623621585
transform 1 0 20700 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_225
timestamp 1623621585
transform 1 0 21804 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_157_237
timestamp 1623621585
transform 1 0 22908 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_249
timestamp 1623621585
transform 1 0 24012 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1534
timestamp 1623621585
transform 1 0 24748 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_258
timestamp 1623621585
transform 1 0 24840 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_157_270
timestamp 1623621585
transform 1 0 25944 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0575_
timestamp 1623621585
transform 1 0 26956 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_157_278
timestamp 1623621585
transform 1 0 26680 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_157_289
timestamp 1623621585
transform 1 0 27692 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0558_
timestamp 1623621585
transform 1 0 28060 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_157_301
timestamp 1623621585
transform 1 0 28796 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0550_
timestamp 1623621585
transform 1 0 31464 0 1 87584
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0651_
timestamp 1623621585
transform 1 0 30728 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1535
timestamp 1623621585
transform 1 0 29992 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_157_313
timestamp 1623621585
transform 1 0 29900 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_157_315
timestamp 1623621585
transform 1 0 30084 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_321
timestamp 1623621585
transform 1 0 30636 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_157_326
timestamp 1623621585
transform 1 0 31096 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0483_
timestamp 1623621585
transform 1 0 33120 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_157_344
timestamp 1623621585
transform 1 0 32752 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_157_352
timestamp 1623621585
transform 1 0 33488 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1536
timestamp 1623621585
transform 1 0 35236 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_157_364
timestamp 1623621585
transform 1 0 34592 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_370
timestamp 1623621585
transform 1 0 35144 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_157_372
timestamp 1623621585
transform 1 0 35328 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input269
timestamp 1623621585
transform 1 0 37260 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_157_384
timestamp 1623621585
transform 1 0 36432 0 1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_157_392
timestamp 1623621585
transform 1 0 37168 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_315
timestamp 1623621585
transform -1 0 38824 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input268
timestamp 1623621585
transform 1 0 37904 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_157_396
timestamp 1623621585
transform 1 0 37536 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_157_403
timestamp 1623621585
transform 1 0 38180 0 1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_316
timestamp 1623621585
transform 1 0 1104 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_318
timestamp 1623621585
transform 1 0 1104 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input429
timestamp 1623621585
transform 1 0 1748 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_158_3
timestamp 1623621585
transform 1 0 1380 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_15
timestamp 1623621585
transform 1 0 2484 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_3
timestamp 1623621585
transform 1 0 1380 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_159_11
timestamp 1623621585
transform 1 0 2116 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1544
timestamp 1623621585
transform 1 0 3772 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_27
timestamp 1623621585
transform 1 0 3588 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_39
timestamp 1623621585
transform 1 0 4692 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_23
timestamp 1623621585
transform 1 0 3220 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_159_30
timestamp 1623621585
transform 1 0 3864 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1537
timestamp 1623621585
transform 1 0 6348 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_158_51
timestamp 1623621585
transform 1 0 5796 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_158_58
timestamp 1623621585
transform 1 0 6440 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_42
timestamp 1623621585
transform 1 0 4968 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_54
timestamp 1623621585
transform 1 0 6072 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_70
timestamp 1623621585
transform 1 0 7544 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_82
timestamp 1623621585
transform 1 0 8648 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_66
timestamp 1623621585
transform 1 0 7176 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_78
timestamp 1623621585
transform 1 0 8280 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1545
timestamp 1623621585
transform 1 0 9016 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_94
timestamp 1623621585
transform 1 0 9752 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_87
timestamp 1623621585
transform 1 0 9108 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_99
timestamp 1623621585
transform 1 0 10212 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1538
timestamp 1623621585
transform 1 0 11592 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_106
timestamp 1623621585
transform 1 0 10856 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_115
timestamp 1623621585
transform 1 0 11684 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_111
timestamp 1623621585
transform 1 0 11316 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_123
timestamp 1623621585
transform 1 0 12420 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1546
timestamp 1623621585
transform 1 0 14260 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_127
timestamp 1623621585
transform 1 0 12788 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_139
timestamp 1623621585
transform 1 0 13892 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_135
timestamp 1623621585
transform 1 0 13524 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_144
timestamp 1623621585
transform 1 0 14352 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_151
timestamp 1623621585
transform 1 0 14996 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_163
timestamp 1623621585
transform 1 0 16100 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_156
timestamp 1623621585
transform 1 0 15456 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1539
timestamp 1623621585
transform 1 0 16836 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_172
timestamp 1623621585
transform 1 0 16928 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_184
timestamp 1623621585
transform 1 0 18032 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_168
timestamp 1623621585
transform 1 0 16560 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_180
timestamp 1623621585
transform 1 0 17664 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1547
timestamp 1623621585
transform 1 0 19504 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_196
timestamp 1623621585
transform 1 0 19136 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_208
timestamp 1623621585
transform 1 0 20240 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_192
timestamp 1623621585
transform 1 0 18768 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_159_201
timestamp 1623621585
transform 1 0 19596 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1540
timestamp 1623621585
transform 1 0 22080 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_220
timestamp 1623621585
transform 1 0 21344 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_158_229
timestamp 1623621585
transform 1 0 22172 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_213
timestamp 1623621585
transform 1 0 20700 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_225
timestamp 1623621585
transform 1 0 21804 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0599_
timestamp 1623621585
transform 1 0 23460 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_158_241
timestamp 1623621585
transform 1 0 23276 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_237
timestamp 1623621585
transform 1 0 22908 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_159_247
timestamp 1623621585
transform 1 0 23828 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1548
timestamp 1623621585
transform 1 0 24748 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_253
timestamp 1623621585
transform 1 0 24380 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_265
timestamp 1623621585
transform 1 0 25484 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_159_255
timestamp 1623621585
transform 1 0 24564 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_159_258
timestamp 1623621585
transform 1 0 24840 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_159_270
timestamp 1623621585
transform 1 0 25944 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1541
timestamp 1623621585
transform 1 0 27324 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_277
timestamp 1623621585
transform 1 0 26588 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_158_286
timestamp 1623621585
transform 1 0 27416 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_159_282
timestamp 1623621585
transform 1 0 27048 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0529_
timestamp 1623621585
transform 1 0 28244 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0549_
timestamp 1623621585
transform 1 0 28060 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0566_
timestamp 1623621585
transform 1 0 29164 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_158_292
timestamp 1623621585
transform 1 0 27968 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_158_301
timestamp 1623621585
transform 1 0 28796 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_294
timestamp 1623621585
transform 1 0 28152 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_159_303
timestamp 1623621585
transform 1 0 28980 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_159_311
timestamp 1623621585
transform 1 0 29716 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0559_
timestamp 1623621585
transform 1 0 30912 0 -1 88672
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1549
timestamp 1623621585
transform 1 0 29992 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_158_313
timestamp 1623621585
transform 1 0 29900 0 -1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_158_321
timestamp 1623621585
transform 1 0 30636 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_159_315
timestamp 1623621585
transform 1 0 30084 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_327
timestamp 1623621585
transform 1 0 31188 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0513_
timestamp 1623621585
transform 1 0 31924 0 1 88672
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0576_
timestamp 1623621585
transform 1 0 33028 0 -1 88672
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1542
timestamp 1623621585
transform 1 0 32568 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_158_338
timestamp 1623621585
transform 1 0 32200 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_158_343
timestamp 1623621585
transform 1 0 32660 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_159_349
timestamp 1623621585
transform 1 0 33212 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1550
timestamp 1623621585
transform 1 0 35236 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_158_361
timestamp 1623621585
transform 1 0 34316 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_158_373
timestamp 1623621585
transform 1 0 35420 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_159_361
timestamp 1623621585
transform 1 0 34316 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_159_369
timestamp 1623621585
transform 1 0 35052 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_159_372
timestamp 1623621585
transform 1 0 35328 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input271
timestamp 1623621585
transform 1 0 37168 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input272
timestamp 1623621585
transform 1 0 37260 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_158_385
timestamp 1623621585
transform 1 0 36524 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_391
timestamp 1623621585
transform 1 0 37076 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_158_395
timestamp 1623621585
transform 1 0 37444 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_159_384
timestamp 1623621585
transform 1 0 36432 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_159_392
timestamp 1623621585
transform 1 0 37168 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_317
timestamp 1623621585
transform -1 0 38824 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_319
timestamp 1623621585
transform -1 0 38824 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1543
timestamp 1623621585
transform 1 0 37812 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input270
timestamp 1623621585
transform 1 0 37904 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_158_400
timestamp 1623621585
transform 1 0 37904 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_406
timestamp 1623621585
transform 1 0 38456 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_159_396
timestamp 1623621585
transform 1 0 37536 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_159_403
timestamp 1623621585
transform 1 0 38180 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_320
timestamp 1623621585
transform 1 0 1104 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input430
timestamp 1623621585
transform 1 0 1748 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_160_3
timestamp 1623621585
transform 1 0 1380 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_160_11
timestamp 1623621585
transform 1 0 2116 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_23
timestamp 1623621585
transform 1 0 3220 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_35
timestamp 1623621585
transform 1 0 4324 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1551
timestamp 1623621585
transform 1 0 6348 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_47
timestamp 1623621585
transform 1 0 5428 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_160_55
timestamp 1623621585
transform 1 0 6164 0 -1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_160_58
timestamp 1623621585
transform 1 0 6440 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_70
timestamp 1623621585
transform 1 0 7544 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_82
timestamp 1623621585
transform 1 0 8648 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_94
timestamp 1623621585
transform 1 0 9752 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1552
timestamp 1623621585
transform 1 0 11592 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_106
timestamp 1623621585
transform 1 0 10856 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_115
timestamp 1623621585
transform 1 0 11684 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_127
timestamp 1623621585
transform 1 0 12788 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_139
timestamp 1623621585
transform 1 0 13892 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_151
timestamp 1623621585
transform 1 0 14996 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_163
timestamp 1623621585
transform 1 0 16100 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1553
timestamp 1623621585
transform 1 0 16836 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_172
timestamp 1623621585
transform 1 0 16928 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_184
timestamp 1623621585
transform 1 0 18032 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_196
timestamp 1623621585
transform 1 0 19136 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_208
timestamp 1623621585
transform 1 0 20240 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1554
timestamp 1623621585
transform 1 0 22080 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_220
timestamp 1623621585
transform 1 0 21344 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_160_229
timestamp 1623621585
transform 1 0 22172 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_241
timestamp 1623621585
transform 1 0 23276 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_253
timestamp 1623621585
transform 1 0 24380 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_265
timestamp 1623621585
transform 1 0 25484 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1555
timestamp 1623621585
transform 1 0 27324 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_160_277
timestamp 1623621585
transform 1 0 26588 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_160_286
timestamp 1623621585
transform 1 0 27416 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0521_
timestamp 1623621585
transform 1 0 28244 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_160_294
timestamp 1623621585
transform 1 0 28152 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_160_303
timestamp 1623621585
transform 1 0 28980 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0530_
timestamp 1623621585
transform 1 0 30912 0 -1 89760
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_160_315
timestamp 1623621585
transform 1 0 30084 0 -1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_160_323
timestamp 1623621585
transform 1 0 30820 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0567_
timestamp 1623621585
transform 1 0 33028 0 -1 89760
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1556
timestamp 1623621585
transform 1 0 32568 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_160_338
timestamp 1623621585
transform 1 0 32200 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_160_343
timestamp 1623621585
transform 1 0 32660 0 -1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_160_361
timestamp 1623621585
transform 1 0 34316 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_373
timestamp 1623621585
transform 1 0 35420 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_160_385
timestamp 1623621585
transform 1 0 36524 0 -1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_321
timestamp 1623621585
transform -1 0 38824 0 -1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1557
timestamp 1623621585
transform 1 0 37812 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_160_397
timestamp 1623621585
transform 1 0 37628 0 -1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_160_400
timestamp 1623621585
transform 1 0 37904 0 -1 89760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_406
timestamp 1623621585
transform 1 0 38456 0 -1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_322
timestamp 1623621585
transform 1 0 1104 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_161_3
timestamp 1623621585
transform 1 0 1380 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_15
timestamp 1623621585
transform 1 0 2484 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1558
timestamp 1623621585
transform 1 0 3772 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_161_27
timestamp 1623621585
transform 1 0 3588 0 1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_161_30
timestamp 1623621585
transform 1 0 3864 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_42
timestamp 1623621585
transform 1 0 4968 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_54
timestamp 1623621585
transform 1 0 6072 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_66
timestamp 1623621585
transform 1 0 7176 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_78
timestamp 1623621585
transform 1 0 8280 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1559
timestamp 1623621585
transform 1 0 9016 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_87
timestamp 1623621585
transform 1 0 9108 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_99
timestamp 1623621585
transform 1 0 10212 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_111
timestamp 1623621585
transform 1 0 11316 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_123
timestamp 1623621585
transform 1 0 12420 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1560
timestamp 1623621585
transform 1 0 14260 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_161_135
timestamp 1623621585
transform 1 0 13524 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_161_144
timestamp 1623621585
transform 1 0 14352 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_156
timestamp 1623621585
transform 1 0 15456 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_168
timestamp 1623621585
transform 1 0 16560 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_180
timestamp 1623621585
transform 1 0 17664 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0787_
timestamp 1623621585
transform 1 0 18584 0 1 89760
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1561
timestamp 1623621585
transform 1 0 19504 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_161_188
timestamp 1623621585
transform 1 0 18400 0 1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_161_196
timestamp 1623621585
transform 1 0 19136 0 1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_161_201
timestamp 1623621585
transform 1 0 19596 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_213
timestamp 1623621585
transform 1 0 20700 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_225
timestamp 1623621585
transform 1 0 21804 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_237
timestamp 1623621585
transform 1 0 22908 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_249
timestamp 1623621585
transform 1 0 24012 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1562
timestamp 1623621585
transform 1 0 24748 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_258
timestamp 1623621585
transform 1 0 24840 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_270
timestamp 1623621585
transform 1 0 25944 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_161_282
timestamp 1623621585
transform 1 0 27048 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0512_
timestamp 1623621585
transform 1 0 28336 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_161_294
timestamp 1623621585
transform 1 0 28152 0 1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_161_304
timestamp 1623621585
transform 1 0 29072 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_161_312
timestamp 1623621585
transform 1 0 29808 0 1 89760
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1563
timestamp 1623621585
transform 1 0 29992 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_315
timestamp 1623621585
transform 1 0 30084 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_161_327
timestamp 1623621585
transform 1 0 31188 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0495_
timestamp 1623621585
transform 1 0 32016 0 1 89760
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_161_335
timestamp 1623621585
transform 1 0 31924 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_350
timestamp 1623621585
transform 1 0 33304 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1564
timestamp 1623621585
transform 1 0 35236 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_161_362
timestamp 1623621585
transform 1 0 34408 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_161_370
timestamp 1623621585
transform 1 0 35144 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_161_372
timestamp 1623621585
transform 1 0 35328 0 1 89760
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input274
timestamp 1623621585
transform 1 0 37260 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_161_384
timestamp 1623621585
transform 1 0 36432 0 1 89760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_161_392
timestamp 1623621585
transform 1 0 37168 0 1 89760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_323
timestamp 1623621585
transform -1 0 38824 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input273
timestamp 1623621585
transform 1 0 37904 0 1 89760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_161_396
timestamp 1623621585
transform 1 0 37536 0 1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_161_403
timestamp 1623621585
transform 1 0 38180 0 1 89760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_324
timestamp 1623621585
transform 1 0 1104 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input431
timestamp 1623621585
transform 1 0 1748 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_162_3
timestamp 1623621585
transform 1 0 1380 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_162_11
timestamp 1623621585
transform 1 0 2116 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_23
timestamp 1623621585
transform 1 0 3220 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_35
timestamp 1623621585
transform 1 0 4324 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1565
timestamp 1623621585
transform 1 0 6348 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_47
timestamp 1623621585
transform 1 0 5428 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_162_55
timestamp 1623621585
transform 1 0 6164 0 -1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_162_58
timestamp 1623621585
transform 1 0 6440 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_70
timestamp 1623621585
transform 1 0 7544 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_82
timestamp 1623621585
transform 1 0 8648 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_94
timestamp 1623621585
transform 1 0 9752 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1566
timestamp 1623621585
transform 1 0 11592 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_106
timestamp 1623621585
transform 1 0 10856 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_162_115
timestamp 1623621585
transform 1 0 11684 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_127
timestamp 1623621585
transform 1 0 12788 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_139
timestamp 1623621585
transform 1 0 13892 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_151
timestamp 1623621585
transform 1 0 14996 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_163
timestamp 1623621585
transform 1 0 16100 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0789_
timestamp 1623621585
transform 1 0 18032 0 -1 90848
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1567
timestamp 1623621585
transform 1 0 16836 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_172
timestamp 1623621585
transform 1 0 16928 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_190
timestamp 1623621585
transform 1 0 18584 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_202
timestamp 1623621585
transform 1 0 19688 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1568
timestamp 1623621585
transform 1 0 22080 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_162_214
timestamp 1623621585
transform 1 0 20792 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_162_226
timestamp 1623621585
transform 1 0 21896 0 -1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_162_229
timestamp 1623621585
transform 1 0 22172 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_241
timestamp 1623621585
transform 1 0 23276 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_253
timestamp 1623621585
transform 1 0 24380 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_265
timestamp 1623621585
transform 1 0 25484 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1569
timestamp 1623621585
transform 1 0 27324 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_162_277
timestamp 1623621585
transform 1 0 26588 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_162_286
timestamp 1623621585
transform 1 0 27416 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0494_
timestamp 1623621585
transform 1 0 28336 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_162_294
timestamp 1623621585
transform 1 0 28152 0 -1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_162_304
timestamp 1623621585
transform 1 0 29072 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0522_
timestamp 1623621585
transform 1 0 30912 0 -1 90848
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_162_316
timestamp 1623621585
transform 1 0 30176 0 -1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0597_
timestamp 1623621585
transform 1 0 33028 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1570
timestamp 1623621585
transform 1 0 32568 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_162_338
timestamp 1623621585
transform 1 0 32200 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_162_343
timestamp 1623621585
transform 1 0 32660 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_162_351
timestamp 1623621585
transform 1 0 33396 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_363
timestamp 1623621585
transform 1 0 34500 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_162_375
timestamp 1623621585
transform 1 0 35604 0 -1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input276
timestamp 1623621585
transform 1 0 37168 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_162_387
timestamp 1623621585
transform 1 0 36708 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_162_391
timestamp 1623621585
transform 1 0 37076 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_162_395
timestamp 1623621585
transform 1 0 37444 0 -1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_325
timestamp 1623621585
transform -1 0 38824 0 -1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1571
timestamp 1623621585
transform 1 0 37812 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_162_400
timestamp 1623621585
transform 1 0 37904 0 -1 90848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_406
timestamp 1623621585
transform 1 0 38456 0 -1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_326
timestamp 1623621585
transform 1 0 1104 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_163_3
timestamp 1623621585
transform 1 0 1380 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_15
timestamp 1623621585
transform 1 0 2484 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1572
timestamp 1623621585
transform 1 0 3772 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_163_27
timestamp 1623621585
transform 1 0 3588 0 1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_163_30
timestamp 1623621585
transform 1 0 3864 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_42
timestamp 1623621585
transform 1 0 4968 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_54
timestamp 1623621585
transform 1 0 6072 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_66
timestamp 1623621585
transform 1 0 7176 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_78
timestamp 1623621585
transform 1 0 8280 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1573
timestamp 1623621585
transform 1 0 9016 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_87
timestamp 1623621585
transform 1 0 9108 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_99
timestamp 1623621585
transform 1 0 10212 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_111
timestamp 1623621585
transform 1 0 11316 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_123
timestamp 1623621585
transform 1 0 12420 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1574
timestamp 1623621585
transform 1 0 14260 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_135
timestamp 1623621585
transform 1 0 13524 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_163_144
timestamp 1623621585
transform 1 0 14352 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_156
timestamp 1623621585
transform 1 0 15456 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_168
timestamp 1623621585
transform 1 0 16560 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_180
timestamp 1623621585
transform 1 0 17664 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1575
timestamp 1623621585
transform 1 0 19504 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_192
timestamp 1623621585
transform 1 0 18768 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_163_201
timestamp 1623621585
transform 1 0 19596 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_213
timestamp 1623621585
transform 1 0 20700 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_225
timestamp 1623621585
transform 1 0 21804 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_237
timestamp 1623621585
transform 1 0 22908 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_249
timestamp 1623621585
transform 1 0 24012 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1576
timestamp 1623621585
transform 1 0 24748 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_258
timestamp 1623621585
transform 1 0 24840 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_270
timestamp 1623621585
transform 1 0 25944 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_163_282
timestamp 1623621585
transform 1 0 27048 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__a221o_1  _0504_
timestamp 1623621585
transform 1 0 28336 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_163_294
timestamp 1623621585
transform 1 0 28152 0 1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_163_304
timestamp 1623621585
transform 1 0 29072 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_163_312
timestamp 1623621585
transform 1 0 29808 0 1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1577
timestamp 1623621585
transform 1 0 29992 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_163_315
timestamp 1623621585
transform 1 0 30084 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_163_327
timestamp 1623621585
transform 1 0 31188 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0505_
timestamp 1623621585
transform 1 0 31924 0 1 90848
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_163_349
timestamp 1623621585
transform 1 0 33212 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1578
timestamp 1623621585
transform 1 0 35236 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_163_361
timestamp 1623621585
transform 1 0 34316 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_163_369
timestamp 1623621585
transform 1 0 35052 0 1 90848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_163_372
timestamp 1623621585
transform 1 0 35328 0 1 90848
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input277
timestamp 1623621585
transform 1 0 37260 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_163_384
timestamp 1623621585
transform 1 0 36432 0 1 90848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_163_392
timestamp 1623621585
transform 1 0 37168 0 1 90848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_327
timestamp 1623621585
transform -1 0 38824 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input275
timestamp 1623621585
transform 1 0 37904 0 1 90848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_163_396
timestamp 1623621585
transform 1 0 37536 0 1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_163_403
timestamp 1623621585
transform 1 0 38180 0 1 90848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_328
timestamp 1623621585
transform 1 0 1104 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input432
timestamp 1623621585
transform 1 0 1748 0 -1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_164_3
timestamp 1623621585
transform 1 0 1380 0 -1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_164_11
timestamp 1623621585
transform 1 0 2116 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_23
timestamp 1623621585
transform 1 0 3220 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_35
timestamp 1623621585
transform 1 0 4324 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1579
timestamp 1623621585
transform 1 0 6348 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_47
timestamp 1623621585
transform 1 0 5428 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_164_55
timestamp 1623621585
transform 1 0 6164 0 -1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_164_58
timestamp 1623621585
transform 1 0 6440 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_70
timestamp 1623621585
transform 1 0 7544 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_82
timestamp 1623621585
transform 1 0 8648 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0948_
timestamp 1623621585
transform 1 0 10672 0 -1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_164_94
timestamp 1623621585
transform 1 0 9752 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_164_102
timestamp 1623621585
transform 1 0 10488 0 -1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1580
timestamp 1623621585
transform 1 0 11592 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_164_108
timestamp 1623621585
transform 1 0 11040 0 -1 91936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_164_115
timestamp 1623621585
transform 1 0 11684 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_127
timestamp 1623621585
transform 1 0 12788 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_139
timestamp 1623621585
transform 1 0 13892 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1623621585
transform 1 0 15732 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_164_151
timestamp 1623621585
transform 1 0 14996 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_164_162
timestamp 1623621585
transform 1 0 16008 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1581
timestamp 1623621585
transform 1 0 16836 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_164_170
timestamp 1623621585
transform 1 0 16744 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_164_172
timestamp 1623621585
transform 1 0 16928 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_184
timestamp 1623621585
transform 1 0 18032 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_196
timestamp 1623621585
transform 1 0 19136 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_208
timestamp 1623621585
transform 1 0 20240 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1582
timestamp 1623621585
transform 1 0 22080 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_220
timestamp 1623621585
transform 1 0 21344 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_229
timestamp 1623621585
transform 1 0 22172 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_241
timestamp 1623621585
transform 1 0 23276 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_253
timestamp 1623621585
transform 1 0 24380 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_265
timestamp 1623621585
transform 1 0 25484 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1583
timestamp 1623621585
transform 1 0 27324 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_277
timestamp 1623621585
transform 1 0 26588 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_286
timestamp 1623621585
transform 1 0 27416 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_298
timestamp 1623621585
transform 1 0 28520 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_310
timestamp 1623621585
transform 1 0 29624 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_322
timestamp 1623621585
transform 1 0 30728 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1584
timestamp 1623621585
transform 1 0 32568 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_164_334
timestamp 1623621585
transform 1 0 31832 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_164_343
timestamp 1623621585
transform 1 0 32660 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_355
timestamp 1623621585
transform 1 0 33764 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_367
timestamp 1623621585
transform 1 0 34868 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_164_379
timestamp 1623621585
transform 1 0 35972 0 -1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_391
timestamp 1623621585
transform 1 0 37076 0 -1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_329
timestamp 1623621585
transform -1 0 38824 0 -1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1585
timestamp 1623621585
transform 1 0 37812 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_164_400
timestamp 1623621585
transform 1 0 37904 0 -1 91936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_406
timestamp 1623621585
transform 1 0 38456 0 -1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_330
timestamp 1623621585
transform 1 0 1104 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_332
timestamp 1623621585
transform 1 0 1104 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input433
timestamp 1623621585
transform 1 0 1748 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_165_3
timestamp 1623621585
transform 1 0 1380 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_165_11
timestamp 1623621585
transform 1 0 2116 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_3
timestamp 1623621585
transform 1 0 1380 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_15
timestamp 1623621585
transform 1 0 2484 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1586
timestamp 1623621585
transform 1 0 3772 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_165_23
timestamp 1623621585
transform 1 0 3220 0 1 91936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_165_30
timestamp 1623621585
transform 1 0 3864 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_27
timestamp 1623621585
transform 1 0 3588 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_39
timestamp 1623621585
transform 1 0 4692 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1593
timestamp 1623621585
transform 1 0 6348 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_42
timestamp 1623621585
transform 1 0 4968 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_54
timestamp 1623621585
transform 1 0 6072 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_51
timestamp 1623621585
transform 1 0 5796 0 -1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_166_58
timestamp 1623621585
transform 1 0 6440 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_66
timestamp 1623621585
transform 1 0 7176 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_78
timestamp 1623621585
transform 1 0 8280 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_70
timestamp 1623621585
transform 1 0 7544 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_82
timestamp 1623621585
transform 1 0 8648 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1587
timestamp 1623621585
transform 1 0 9016 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_87
timestamp 1623621585
transform 1 0 9108 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_99
timestamp 1623621585
transform 1 0 10212 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_94
timestamp 1623621585
transform 1 0 9752 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1594
timestamp 1623621585
transform 1 0 11592 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_111
timestamp 1623621585
transform 1 0 11316 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_123
timestamp 1623621585
transform 1 0 12420 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_106
timestamp 1623621585
transform 1 0 10856 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_115
timestamp 1623621585
transform 1 0 11684 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1588
timestamp 1623621585
transform 1 0 14260 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_135
timestamp 1623621585
transform 1 0 13524 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_144
timestamp 1623621585
transform 1 0 14352 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_127
timestamp 1623621585
transform 1 0 12788 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_139
timestamp 1623621585
transform 1 0 13892 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_156
timestamp 1623621585
transform 1 0 15456 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_151
timestamp 1623621585
transform 1 0 14996 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_163
timestamp 1623621585
transform 1 0 16100 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1595
timestamp 1623621585
transform 1 0 16836 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_168
timestamp 1623621585
transform 1 0 16560 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_180
timestamp 1623621585
transform 1 0 17664 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_172
timestamp 1623621585
transform 1 0 16928 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_184
timestamp 1623621585
transform 1 0 18032 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _0781_
timestamp 1623621585
transform 1 0 19964 0 1 91936
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1589
timestamp 1623621585
transform 1 0 19504 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_192
timestamp 1623621585
transform 1 0 18768 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_165_201
timestamp 1623621585
transform 1 0 19596 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_166_196
timestamp 1623621585
transform 1 0 19136 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_208
timestamp 1623621585
transform 1 0 20240 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1596
timestamp 1623621585
transform 1 0 22080 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_211
timestamp 1623621585
transform 1 0 20516 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_223
timestamp 1623621585
transform 1 0 21620 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_220
timestamp 1623621585
transform 1 0 21344 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_229
timestamp 1623621585
transform 1 0 22172 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_235
timestamp 1623621585
transform 1 0 22724 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_247
timestamp 1623621585
transform 1 0 23828 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_241
timestamp 1623621585
transform 1 0 23276 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1590
timestamp 1623621585
transform 1 0 24748 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_165_255
timestamp 1623621585
transform 1 0 24564 0 1 91936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_165_258
timestamp 1623621585
transform 1 0 24840 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_270
timestamp 1623621585
transform 1 0 25944 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_253
timestamp 1623621585
transform 1 0 24380 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_265
timestamp 1623621585
transform 1 0 25484 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1597
timestamp 1623621585
transform 1 0 27324 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_282
timestamp 1623621585
transform 1 0 27048 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_277
timestamp 1623621585
transform 1 0 26588 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_286
timestamp 1623621585
transform 1 0 27416 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_294
timestamp 1623621585
transform 1 0 28152 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_165_306
timestamp 1623621585
transform 1 0 29256 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_298
timestamp 1623621585
transform 1 0 28520 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_310
timestamp 1623621585
transform 1 0 29624 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1591
timestamp 1623621585
transform 1 0 29992 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_315
timestamp 1623621585
transform 1 0 30084 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_327
timestamp 1623621585
transform 1 0 31188 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_322
timestamp 1623621585
transform 1 0 30728 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1598
timestamp 1623621585
transform 1 0 32568 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_165_339
timestamp 1623621585
transform 1 0 32292 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_165_351
timestamp 1623621585
transform 1 0 33396 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_334
timestamp 1623621585
transform 1 0 31832 0 -1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_166_343
timestamp 1623621585
transform 1 0 32660 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1592
timestamp 1623621585
transform 1 0 35236 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_165_363
timestamp 1623621585
transform 1 0 34500 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_165_372
timestamp 1623621585
transform 1 0 35328 0 1 91936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_355
timestamp 1623621585
transform 1 0 33764 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_166_367
timestamp 1623621585
transform 1 0 34868 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input280
timestamp 1623621585
transform 1 0 37260 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input282
timestamp 1623621585
transform 1 0 37168 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_165_384
timestamp 1623621585
transform 1 0 36432 0 1 91936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_165_392
timestamp 1623621585
transform 1 0 37168 0 1 91936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_166_379
timestamp 1623621585
transform 1 0 35972 0 -1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_391
timestamp 1623621585
transform 1 0 37076 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_166_395
timestamp 1623621585
transform 1 0 37444 0 -1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_331
timestamp 1623621585
transform -1 0 38824 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_333
timestamp 1623621585
transform -1 0 38824 0 -1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1599
timestamp 1623621585
transform 1 0 37812 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input279
timestamp 1623621585
transform 1 0 37904 0 1 91936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_165_396
timestamp 1623621585
transform 1 0 37536 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_165_403
timestamp 1623621585
transform 1 0 38180 0 1 91936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_166_400
timestamp 1623621585
transform 1 0 37904 0 -1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_406
timestamp 1623621585
transform 1 0 38456 0 -1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_334
timestamp 1623621585
transform 1 0 1104 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input434
timestamp 1623621585
transform 1 0 1748 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_167_3
timestamp 1623621585
transform 1 0 1380 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_167_11
timestamp 1623621585
transform 1 0 2116 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1600
timestamp 1623621585
transform 1 0 3772 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_167_23
timestamp 1623621585
transform 1 0 3220 0 1 93024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_167_30
timestamp 1623621585
transform 1 0 3864 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_42
timestamp 1623621585
transform 1 0 4968 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_54
timestamp 1623621585
transform 1 0 6072 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_66
timestamp 1623621585
transform 1 0 7176 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_78
timestamp 1623621585
transform 1 0 8280 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1601
timestamp 1623621585
transform 1 0 9016 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_87
timestamp 1623621585
transform 1 0 9108 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_99
timestamp 1623621585
transform 1 0 10212 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_111
timestamp 1623621585
transform 1 0 11316 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_123
timestamp 1623621585
transform 1 0 12420 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1602
timestamp 1623621585
transform 1 0 14260 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_135
timestamp 1623621585
transform 1 0 13524 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_144
timestamp 1623621585
transform 1 0 14352 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_156
timestamp 1623621585
transform 1 0 15456 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_168
timestamp 1623621585
transform 1 0 16560 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_180
timestamp 1623621585
transform 1 0 17664 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1603
timestamp 1623621585
transform 1 0 19504 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_192
timestamp 1623621585
transform 1 0 18768 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_201
timestamp 1623621585
transform 1 0 19596 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_213
timestamp 1623621585
transform 1 0 20700 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_225
timestamp 1623621585
transform 1 0 21804 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_237
timestamp 1623621585
transform 1 0 22908 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_249
timestamp 1623621585
transform 1 0 24012 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1604
timestamp 1623621585
transform 1 0 24748 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_258
timestamp 1623621585
transform 1 0 24840 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_270
timestamp 1623621585
transform 1 0 25944 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_282
timestamp 1623621585
transform 1 0 27048 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_294
timestamp 1623621585
transform 1 0 28152 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_167_306
timestamp 1623621585
transform 1 0 29256 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1605
timestamp 1623621585
transform 1 0 29992 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_167_315
timestamp 1623621585
transform 1 0 30084 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_327
timestamp 1623621585
transform 1 0 31188 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_339
timestamp 1623621585
transform 1 0 32292 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_167_351
timestamp 1623621585
transform 1 0 33396 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1606
timestamp 1623621585
transform 1 0 35236 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_167_363
timestamp 1623621585
transform 1 0 34500 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_167_372
timestamp 1623621585
transform 1 0 35328 0 1 93024
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input283
timestamp 1623621585
transform 1 0 37260 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_167_384
timestamp 1623621585
transform 1 0 36432 0 1 93024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_167_392
timestamp 1623621585
transform 1 0 37168 0 1 93024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_335
timestamp 1623621585
transform -1 0 38824 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input281
timestamp 1623621585
transform 1 0 37904 0 1 93024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_167_396
timestamp 1623621585
transform 1 0 37536 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_167_403
timestamp 1623621585
transform 1 0 38180 0 1 93024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_336
timestamp 1623621585
transform 1 0 1104 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input435
timestamp 1623621585
transform 1 0 1748 0 -1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_168_3
timestamp 1623621585
transform 1 0 1380 0 -1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_168_11
timestamp 1623621585
transform 1 0 2116 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_23
timestamp 1623621585
transform 1 0 3220 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_35
timestamp 1623621585
transform 1 0 4324 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1607
timestamp 1623621585
transform 1 0 6348 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_47
timestamp 1623621585
transform 1 0 5428 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_168_55
timestamp 1623621585
transform 1 0 6164 0 -1 94112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_168_58
timestamp 1623621585
transform 1 0 6440 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_70
timestamp 1623621585
transform 1 0 7544 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_82
timestamp 1623621585
transform 1 0 8648 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_94
timestamp 1623621585
transform 1 0 9752 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1608
timestamp 1623621585
transform 1 0 11592 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_106
timestamp 1623621585
transform 1 0 10856 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_115
timestamp 1623621585
transform 1 0 11684 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_127
timestamp 1623621585
transform 1 0 12788 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_139
timestamp 1623621585
transform 1 0 13892 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_151
timestamp 1623621585
transform 1 0 14996 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_163
timestamp 1623621585
transform 1 0 16100 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1609
timestamp 1623621585
transform 1 0 16836 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_168_172
timestamp 1623621585
transform 1 0 16928 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_184
timestamp 1623621585
transform 1 0 18032 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_196
timestamp 1623621585
transform 1 0 19136 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_208
timestamp 1623621585
transform 1 0 20240 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1610
timestamp 1623621585
transform 1 0 22080 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_220
timestamp 1623621585
transform 1 0 21344 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_229
timestamp 1623621585
transform 1 0 22172 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_241
timestamp 1623621585
transform 1 0 23276 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_253
timestamp 1623621585
transform 1 0 24380 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_265
timestamp 1623621585
transform 1 0 25484 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1611
timestamp 1623621585
transform 1 0 27324 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_277
timestamp 1623621585
transform 1 0 26588 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_286
timestamp 1623621585
transform 1 0 27416 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_298
timestamp 1623621585
transform 1 0 28520 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_310
timestamp 1623621585
transform 1 0 29624 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_322
timestamp 1623621585
transform 1 0 30728 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1612
timestamp 1623621585
transform 1 0 32568 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_168_334
timestamp 1623621585
transform 1 0 31832 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_168_343
timestamp 1623621585
transform 1 0 32660 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_355
timestamp 1623621585
transform 1 0 33764 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_367
timestamp 1623621585
transform 1 0 34868 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_168_379
timestamp 1623621585
transform 1 0 35972 0 -1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_391
timestamp 1623621585
transform 1 0 37076 0 -1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_337
timestamp 1623621585
transform -1 0 38824 0 -1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1613
timestamp 1623621585
transform 1 0 37812 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_168_400
timestamp 1623621585
transform 1 0 37904 0 -1 94112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_406
timestamp 1623621585
transform 1 0 38456 0 -1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_338
timestamp 1623621585
transform 1 0 1104 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_169_3
timestamp 1623621585
transform 1 0 1380 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_15
timestamp 1623621585
transform 1 0 2484 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1614
timestamp 1623621585
transform 1 0 3772 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_169_27
timestamp 1623621585
transform 1 0 3588 0 1 94112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_169_30
timestamp 1623621585
transform 1 0 3864 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_42
timestamp 1623621585
transform 1 0 4968 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_54
timestamp 1623621585
transform 1 0 6072 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_66
timestamp 1623621585
transform 1 0 7176 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_78
timestamp 1623621585
transform 1 0 8280 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1615
timestamp 1623621585
transform 1 0 9016 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_87
timestamp 1623621585
transform 1 0 9108 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_99
timestamp 1623621585
transform 1 0 10212 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_111
timestamp 1623621585
transform 1 0 11316 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_123
timestamp 1623621585
transform 1 0 12420 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1616
timestamp 1623621585
transform 1 0 14260 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_135
timestamp 1623621585
transform 1 0 13524 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_144
timestamp 1623621585
transform 1 0 14352 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_156
timestamp 1623621585
transform 1 0 15456 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_168
timestamp 1623621585
transform 1 0 16560 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_180
timestamp 1623621585
transform 1 0 17664 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1617
timestamp 1623621585
transform 1 0 19504 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_192
timestamp 1623621585
transform 1 0 18768 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_201
timestamp 1623621585
transform 1 0 19596 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_213
timestamp 1623621585
transform 1 0 20700 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_225
timestamp 1623621585
transform 1 0 21804 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_237
timestamp 1623621585
transform 1 0 22908 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_249
timestamp 1623621585
transform 1 0 24012 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1618
timestamp 1623621585
transform 1 0 24748 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_258
timestamp 1623621585
transform 1 0 24840 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_270
timestamp 1623621585
transform 1 0 25944 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_282
timestamp 1623621585
transform 1 0 27048 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_294
timestamp 1623621585
transform 1 0 28152 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_169_306
timestamp 1623621585
transform 1 0 29256 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1619
timestamp 1623621585
transform 1 0 29992 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_169_315
timestamp 1623621585
transform 1 0 30084 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_327
timestamp 1623621585
transform 1 0 31188 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_339
timestamp 1623621585
transform 1 0 32292 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_169_351
timestamp 1623621585
transform 1 0 33396 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1620
timestamp 1623621585
transform 1 0 35236 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_169_363
timestamp 1623621585
transform 1 0 34500 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_169_372
timestamp 1623621585
transform 1 0 35328 0 1 94112
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input285
timestamp 1623621585
transform 1 0 37260 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_169_384
timestamp 1623621585
transform 1 0 36432 0 1 94112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_169_392
timestamp 1623621585
transform 1 0 37168 0 1 94112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_339
timestamp 1623621585
transform -1 0 38824 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input284
timestamp 1623621585
transform 1 0 37904 0 1 94112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_169_396
timestamp 1623621585
transform 1 0 37536 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_169_403
timestamp 1623621585
transform 1 0 38180 0 1 94112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_340
timestamp 1623621585
transform 1 0 1104 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input436
timestamp 1623621585
transform 1 0 1748 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_170_3
timestamp 1623621585
transform 1 0 1380 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_170_11
timestamp 1623621585
transform 1 0 2116 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_23
timestamp 1623621585
transform 1 0 3220 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_35
timestamp 1623621585
transform 1 0 4324 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1621
timestamp 1623621585
transform 1 0 6348 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_47
timestamp 1623621585
transform 1 0 5428 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_170_55
timestamp 1623621585
transform 1 0 6164 0 -1 95200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_170_58
timestamp 1623621585
transform 1 0 6440 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_70
timestamp 1623621585
transform 1 0 7544 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_82
timestamp 1623621585
transform 1 0 8648 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_94
timestamp 1623621585
transform 1 0 9752 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1622
timestamp 1623621585
transform 1 0 11592 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_106
timestamp 1623621585
transform 1 0 10856 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_115
timestamp 1623621585
transform 1 0 11684 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_127
timestamp 1623621585
transform 1 0 12788 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_139
timestamp 1623621585
transform 1 0 13892 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_151
timestamp 1623621585
transform 1 0 14996 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_163
timestamp 1623621585
transform 1 0 16100 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1623
timestamp 1623621585
transform 1 0 16836 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_170_172
timestamp 1623621585
transform 1 0 16928 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_184
timestamp 1623621585
transform 1 0 18032 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_196
timestamp 1623621585
transform 1 0 19136 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_208
timestamp 1623621585
transform 1 0 20240 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1624
timestamp 1623621585
transform 1 0 22080 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_220
timestamp 1623621585
transform 1 0 21344 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_229
timestamp 1623621585
transform 1 0 22172 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_241
timestamp 1623621585
transform 1 0 23276 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_253
timestamp 1623621585
transform 1 0 24380 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_265
timestamp 1623621585
transform 1 0 25484 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1625
timestamp 1623621585
transform 1 0 27324 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_277
timestamp 1623621585
transform 1 0 26588 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_286
timestamp 1623621585
transform 1 0 27416 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_298
timestamp 1623621585
transform 1 0 28520 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_310
timestamp 1623621585
transform 1 0 29624 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_322
timestamp 1623621585
transform 1 0 30728 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1626
timestamp 1623621585
transform 1 0 32568 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_170_334
timestamp 1623621585
transform 1 0 31832 0 -1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_170_343
timestamp 1623621585
transform 1 0 32660 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_355
timestamp 1623621585
transform 1 0 33764 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_170_367
timestamp 1623621585
transform 1 0 34868 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input287
timestamp 1623621585
transform 1 0 37168 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_170_379
timestamp 1623621585
transform 1 0 35972 0 -1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_391
timestamp 1623621585
transform 1 0 37076 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_170_395
timestamp 1623621585
transform 1 0 37444 0 -1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_341
timestamp 1623621585
transform -1 0 38824 0 -1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1627
timestamp 1623621585
transform 1 0 37812 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_170_400
timestamp 1623621585
transform 1 0 37904 0 -1 95200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_406
timestamp 1623621585
transform 1 0 38456 0 -1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_342
timestamp 1623621585
transform 1 0 1104 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_344
timestamp 1623621585
transform 1 0 1104 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input437
timestamp 1623621585
transform 1 0 1748 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_171_3
timestamp 1623621585
transform 1 0 1380 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_171_11
timestamp 1623621585
transform 1 0 2116 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_3
timestamp 1623621585
transform 1 0 1380 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_15
timestamp 1623621585
transform 1 0 2484 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1628
timestamp 1623621585
transform 1 0 3772 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_171_23
timestamp 1623621585
transform 1 0 3220 0 1 95200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_171_30
timestamp 1623621585
transform 1 0 3864 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_27
timestamp 1623621585
transform 1 0 3588 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_39
timestamp 1623621585
transform 1 0 4692 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1635
timestamp 1623621585
transform 1 0 6348 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_42
timestamp 1623621585
transform 1 0 4968 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_54
timestamp 1623621585
transform 1 0 6072 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_51
timestamp 1623621585
transform 1 0 5796 0 -1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_172_58
timestamp 1623621585
transform 1 0 6440 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_66
timestamp 1623621585
transform 1 0 7176 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_78
timestamp 1623621585
transform 1 0 8280 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_70
timestamp 1623621585
transform 1 0 7544 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_82
timestamp 1623621585
transform 1 0 8648 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1629
timestamp 1623621585
transform 1 0 9016 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_87
timestamp 1623621585
transform 1 0 9108 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_99
timestamp 1623621585
transform 1 0 10212 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_94
timestamp 1623621585
transform 1 0 9752 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1636
timestamp 1623621585
transform 1 0 11592 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_111
timestamp 1623621585
transform 1 0 11316 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_123
timestamp 1623621585
transform 1 0 12420 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_106
timestamp 1623621585
transform 1 0 10856 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_115
timestamp 1623621585
transform 1 0 11684 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1630
timestamp 1623621585
transform 1 0 14260 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_135
timestamp 1623621585
transform 1 0 13524 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_144
timestamp 1623621585
transform 1 0 14352 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_127
timestamp 1623621585
transform 1 0 12788 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_139
timestamp 1623621585
transform 1 0 13892 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_156
timestamp 1623621585
transform 1 0 15456 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_151
timestamp 1623621585
transform 1 0 14996 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_163
timestamp 1623621585
transform 1 0 16100 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1637
timestamp 1623621585
transform 1 0 16836 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_168
timestamp 1623621585
transform 1 0 16560 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_180
timestamp 1623621585
transform 1 0 17664 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_172
timestamp 1623621585
transform 1 0 16928 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_184
timestamp 1623621585
transform 1 0 18032 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1631
timestamp 1623621585
transform 1 0 19504 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_192
timestamp 1623621585
transform 1 0 18768 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_201
timestamp 1623621585
transform 1 0 19596 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_196
timestamp 1623621585
transform 1 0 19136 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_208
timestamp 1623621585
transform 1 0 20240 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1638
timestamp 1623621585
transform 1 0 22080 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_213
timestamp 1623621585
transform 1 0 20700 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_225
timestamp 1623621585
transform 1 0 21804 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_172_220
timestamp 1623621585
transform 1 0 21344 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_229
timestamp 1623621585
transform 1 0 22172 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _0796_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 22816 0 1 95200
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_171_233
timestamp 1623621585
transform 1 0 22540 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_249
timestamp 1623621585
transform 1 0 24012 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_241
timestamp 1623621585
transform 1 0 23276 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1632
timestamp 1623621585
transform 1 0 24748 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_258
timestamp 1623621585
transform 1 0 24840 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_270
timestamp 1623621585
transform 1 0 25944 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_253
timestamp 1623621585
transform 1 0 24380 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_265
timestamp 1623621585
transform 1 0 25484 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1639
timestamp 1623621585
transform 1 0 27324 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_282
timestamp 1623621585
transform 1 0 27048 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_277
timestamp 1623621585
transform 1 0 26588 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_286
timestamp 1623621585
transform 1 0 27416 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_294
timestamp 1623621585
transform 1 0 28152 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_171_306
timestamp 1623621585
transform 1 0 29256 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_298
timestamp 1623621585
transform 1 0 28520 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_310
timestamp 1623621585
transform 1 0 29624 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1633
timestamp 1623621585
transform 1 0 29992 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_315
timestamp 1623621585
transform 1 0 30084 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_327
timestamp 1623621585
transform 1 0 31188 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_322
timestamp 1623621585
transform 1 0 30728 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1640
timestamp 1623621585
transform 1 0 32568 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_171_339
timestamp 1623621585
transform 1 0 32292 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_171_351
timestamp 1623621585
transform 1 0 33396 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_334
timestamp 1623621585
transform 1 0 31832 0 -1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_172_343
timestamp 1623621585
transform 1 0 32660 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1634
timestamp 1623621585
transform 1 0 35236 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_171_363
timestamp 1623621585
transform 1 0 34500 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_171_372
timestamp 1623621585
transform 1 0 35328 0 1 95200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_355
timestamp 1623621585
transform 1 0 33764 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_172_367
timestamp 1623621585
transform 1 0 34868 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input288
timestamp 1623621585
transform 1 0 37260 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input290
timestamp 1623621585
transform 1 0 37168 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_171_384
timestamp 1623621585
transform 1 0 36432 0 1 95200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_171_392
timestamp 1623621585
transform 1 0 37168 0 1 95200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_172_379
timestamp 1623621585
transform 1 0 35972 0 -1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_391
timestamp 1623621585
transform 1 0 37076 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_172_395
timestamp 1623621585
transform 1 0 37444 0 -1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_343
timestamp 1623621585
transform -1 0 38824 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_345
timestamp 1623621585
transform -1 0 38824 0 -1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1641
timestamp 1623621585
transform 1 0 37812 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input286
timestamp 1623621585
transform 1 0 37904 0 1 95200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_171_396
timestamp 1623621585
transform 1 0 37536 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_171_403
timestamp 1623621585
transform 1 0 38180 0 1 95200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_172_400
timestamp 1623621585
transform 1 0 37904 0 -1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_406
timestamp 1623621585
transform 1 0 38456 0 -1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_346
timestamp 1623621585
transform 1 0 1104 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input439
timestamp 1623621585
transform 1 0 1748 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_173_3
timestamp 1623621585
transform 1 0 1380 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_173_11
timestamp 1623621585
transform 1 0 2116 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1642
timestamp 1623621585
transform 1 0 3772 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_173_23
timestamp 1623621585
transform 1 0 3220 0 1 96288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_173_30
timestamp 1623621585
transform 1 0 3864 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_42
timestamp 1623621585
transform 1 0 4968 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_54
timestamp 1623621585
transform 1 0 6072 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_66
timestamp 1623621585
transform 1 0 7176 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_78
timestamp 1623621585
transform 1 0 8280 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1643
timestamp 1623621585
transform 1 0 9016 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_87
timestamp 1623621585
transform 1 0 9108 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_99
timestamp 1623621585
transform 1 0 10212 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_111
timestamp 1623621585
transform 1 0 11316 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_123
timestamp 1623621585
transform 1 0 12420 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1644
timestamp 1623621585
transform 1 0 14260 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_135
timestamp 1623621585
transform 1 0 13524 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_144
timestamp 1623621585
transform 1 0 14352 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_156
timestamp 1623621585
transform 1 0 15456 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0792_
timestamp 1623621585
transform 1 0 18032 0 1 96288
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_173_168
timestamp 1623621585
transform 1 0 16560 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_180
timestamp 1623621585
transform 1 0 17664 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1645
timestamp 1623621585
transform 1 0 19504 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_191
timestamp 1623621585
transform 1 0 18676 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_173_199
timestamp 1623621585
transform 1 0 19412 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_201
timestamp 1623621585
transform 1 0 19596 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_213
timestamp 1623621585
transform 1 0 20700 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_225
timestamp 1623621585
transform 1 0 21804 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_237
timestamp 1623621585
transform 1 0 22908 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_249
timestamp 1623621585
transform 1 0 24012 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1646
timestamp 1623621585
transform 1 0 24748 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_258
timestamp 1623621585
transform 1 0 24840 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_270
timestamp 1623621585
transform 1 0 25944 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_282
timestamp 1623621585
transform 1 0 27048 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_294
timestamp 1623621585
transform 1 0 28152 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_173_306
timestamp 1623621585
transform 1 0 29256 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1647
timestamp 1623621585
transform 1 0 29992 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_173_315
timestamp 1623621585
transform 1 0 30084 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_327
timestamp 1623621585
transform 1 0 31188 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_339
timestamp 1623621585
transform 1 0 32292 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_173_351
timestamp 1623621585
transform 1 0 33396 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1648
timestamp 1623621585
transform 1 0 35236 0 1 96288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_173_363
timestamp 1623621585
transform 1 0 34500 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_173_372
timestamp 1623621585
transform 1 0 35328 0 1 96288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input291
timestamp 1623621585
transform 1 0 37168 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_173_384
timestamp 1623621585
transform 1 0 36432 0 1 96288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_173_395
timestamp 1623621585
transform 1 0 37444 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_347
timestamp 1623621585
transform -1 0 38824 0 1 96288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input299
timestamp 1623621585
transform 1 0 37812 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_173_403
timestamp 1623621585
transform 1 0 38180 0 1 96288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_348
timestamp 1623621585
transform 1 0 1104 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input440
timestamp 1623621585
transform 1 0 1748 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_174_3
timestamp 1623621585
transform 1 0 1380 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_174_11
timestamp 1623621585
transform 1 0 2116 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_23
timestamp 1623621585
transform 1 0 3220 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_35
timestamp 1623621585
transform 1 0 4324 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1649
timestamp 1623621585
transform 1 0 6348 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_47
timestamp 1623621585
transform 1 0 5428 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_174_55
timestamp 1623621585
transform 1 0 6164 0 -1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_174_58
timestamp 1623621585
transform 1 0 6440 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_70
timestamp 1623621585
transform 1 0 7544 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_82
timestamp 1623621585
transform 1 0 8648 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_94
timestamp 1623621585
transform 1 0 9752 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1650
timestamp 1623621585
transform 1 0 11592 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_106
timestamp 1623621585
transform 1 0 10856 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_115
timestamp 1623621585
transform 1 0 11684 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_127
timestamp 1623621585
transform 1 0 12788 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_139
timestamp 1623621585
transform 1 0 13892 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_151
timestamp 1623621585
transform 1 0 14996 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_163
timestamp 1623621585
transform 1 0 16100 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1651
timestamp 1623621585
transform 1 0 16836 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_174_172
timestamp 1623621585
transform 1 0 16928 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_184
timestamp 1623621585
transform 1 0 18032 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_196
timestamp 1623621585
transform 1 0 19136 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_208
timestamp 1623621585
transform 1 0 20240 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1652
timestamp 1623621585
transform 1 0 22080 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_220
timestamp 1623621585
transform 1 0 21344 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_229
timestamp 1623621585
transform 1 0 22172 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_241
timestamp 1623621585
transform 1 0 23276 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_253
timestamp 1623621585
transform 1 0 24380 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_265
timestamp 1623621585
transform 1 0 25484 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1653
timestamp 1623621585
transform 1 0 27324 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_277
timestamp 1623621585
transform 1 0 26588 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_286
timestamp 1623621585
transform 1 0 27416 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_298
timestamp 1623621585
transform 1 0 28520 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_310
timestamp 1623621585
transform 1 0 29624 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_322
timestamp 1623621585
transform 1 0 30728 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1654
timestamp 1623621585
transform 1 0 32568 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_174_334
timestamp 1623621585
transform 1 0 31832 0 -1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_174_343
timestamp 1623621585
transform 1 0 32660 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_355
timestamp 1623621585
transform 1 0 33764 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_174_367
timestamp 1623621585
transform 1 0 34868 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input310
timestamp 1623621585
transform 1 0 37076 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_174_379
timestamp 1623621585
transform 1 0 35972 0 -1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_174_395
timestamp 1623621585
transform 1 0 37444 0 -1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_349
timestamp 1623621585
transform -1 0 38824 0 -1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1655
timestamp 1623621585
transform 1 0 37812 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_174_400
timestamp 1623621585
transform 1 0 37904 0 -1 97376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_406
timestamp 1623621585
transform 1 0 38456 0 -1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_350
timestamp 1623621585
transform 1 0 1104 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_3
timestamp 1623621585
transform 1 0 1380 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_15
timestamp 1623621585
transform 1 0 2484 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1656
timestamp 1623621585
transform 1 0 3772 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_175_27
timestamp 1623621585
transform 1 0 3588 0 1 97376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_175_30
timestamp 1623621585
transform 1 0 3864 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_42
timestamp 1623621585
transform 1 0 4968 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_54
timestamp 1623621585
transform 1 0 6072 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_66
timestamp 1623621585
transform 1 0 7176 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_78
timestamp 1623621585
transform 1 0 8280 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1657
timestamp 1623621585
transform 1 0 9016 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_87
timestamp 1623621585
transform 1 0 9108 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_99
timestamp 1623621585
transform 1 0 10212 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_111
timestamp 1623621585
transform 1 0 11316 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_123
timestamp 1623621585
transform 1 0 12420 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1658
timestamp 1623621585
transform 1 0 14260 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_175_135
timestamp 1623621585
transform 1 0 13524 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_175_144
timestamp 1623621585
transform 1 0 14352 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0783_
timestamp 1623621585
transform 1 0 16284 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0785_
timestamp 1623621585
transform 1 0 14720 0 1 97376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_175_154
timestamp 1623621585
transform 1 0 15272 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_175_162
timestamp 1623621585
transform 1 0 16008 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_175_169
timestamp 1623621585
transform 1 0 16652 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_181
timestamp 1623621585
transform 1 0 17756 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1659
timestamp 1623621585
transform 1 0 19504 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_175_193
timestamp 1623621585
transform 1 0 18860 0 1 97376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_199
timestamp 1623621585
transform 1 0 19412 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_201
timestamp 1623621585
transform 1 0 19596 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_213
timestamp 1623621585
transform 1 0 20700 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_225
timestamp 1623621585
transform 1 0 21804 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_237
timestamp 1623621585
transform 1 0 22908 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_249
timestamp 1623621585
transform 1 0 24012 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1660
timestamp 1623621585
transform 1 0 24748 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_258
timestamp 1623621585
transform 1 0 24840 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_270
timestamp 1623621585
transform 1 0 25944 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_282
timestamp 1623621585
transform 1 0 27048 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_294
timestamp 1623621585
transform 1 0 28152 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_175_306
timestamp 1623621585
transform 1 0 29256 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1661
timestamp 1623621585
transform 1 0 29992 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_175_315
timestamp 1623621585
transform 1 0 30084 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_327
timestamp 1623621585
transform 1 0 31188 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_339
timestamp 1623621585
transform 1 0 32292 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_351
timestamp 1623621585
transform 1 0 33396 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1662
timestamp 1623621585
transform 1 0 35236 0 1 97376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_175_363
timestamp 1623621585
transform 1 0 34500 0 1 97376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_175_372
timestamp 1623621585
transform 1 0 35328 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_175_384
timestamp 1623621585
transform 1 0 36432 0 1 97376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_351
timestamp 1623621585
transform -1 0 38824 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input321
timestamp 1623621585
transform 1 0 37812 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_175_396
timestamp 1623621585
transform 1 0 37536 0 1 97376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_175_403
timestamp 1623621585
transform 1 0 38180 0 1 97376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_352
timestamp 1623621585
transform 1 0 1104 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input441
timestamp 1623621585
transform 1 0 1748 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_176_3
timestamp 1623621585
transform 1 0 1380 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_176_11
timestamp 1623621585
transform 1 0 2116 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_23
timestamp 1623621585
transform 1 0 3220 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_35
timestamp 1623621585
transform 1 0 4324 0 -1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_41
timestamp 1623621585
transform 1 0 4876 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0935_
timestamp 1623621585
transform 1 0 4968 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1663
timestamp 1623621585
transform 1 0 6348 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_45
timestamp 1623621585
transform 1 0 5244 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_58
timestamp 1623621585
transform 1 0 6440 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_70
timestamp 1623621585
transform 1 0 7544 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_82
timestamp 1623621585
transform 1 0 8648 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_94
timestamp 1623621585
transform 1 0 9752 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1664
timestamp 1623621585
transform 1 0 11592 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_106
timestamp 1623621585
transform 1 0 10856 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_115
timestamp 1623621585
transform 1 0 11684 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_127
timestamp 1623621585
transform 1 0 12788 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_139
timestamp 1623621585
transform 1 0 13892 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_151
timestamp 1623621585
transform 1 0 14996 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_163
timestamp 1623621585
transform 1 0 16100 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1665
timestamp 1623621585
transform 1 0 16836 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_176_172
timestamp 1623621585
transform 1 0 16928 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_184
timestamp 1623621585
transform 1 0 18032 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_196
timestamp 1623621585
transform 1 0 19136 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_208
timestamp 1623621585
transform 1 0 20240 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1666
timestamp 1623621585
transform 1 0 22080 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_220
timestamp 1623621585
transform 1 0 21344 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_229
timestamp 1623621585
transform 1 0 22172 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_241
timestamp 1623621585
transform 1 0 23276 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_253
timestamp 1623621585
transform 1 0 24380 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_265
timestamp 1623621585
transform 1 0 25484 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1667
timestamp 1623621585
transform 1 0 27324 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_277
timestamp 1623621585
transform 1 0 26588 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_286
timestamp 1623621585
transform 1 0 27416 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_298
timestamp 1623621585
transform 1 0 28520 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_310
timestamp 1623621585
transform 1 0 29624 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_322
timestamp 1623621585
transform 1 0 30728 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1668
timestamp 1623621585
transform 1 0 32568 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_176_334
timestamp 1623621585
transform 1 0 31832 0 -1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_176_343
timestamp 1623621585
transform 1 0 32660 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_355
timestamp 1623621585
transform 1 0 33764 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_176_367
timestamp 1623621585
transform 1 0 34868 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input324
timestamp 1623621585
transform 1 0 37076 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_176_379
timestamp 1623621585
transform 1 0 35972 0 -1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_176_395
timestamp 1623621585
transform 1 0 37444 0 -1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_353
timestamp 1623621585
transform -1 0 38824 0 -1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1669
timestamp 1623621585
transform 1 0 37812 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_176_400
timestamp 1623621585
transform 1 0 37904 0 -1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_406
timestamp 1623621585
transform 1 0 38456 0 -1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_354
timestamp 1623621585
transform 1 0 1104 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input442
timestamp 1623621585
transform 1 0 1748 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_177_3
timestamp 1623621585
transform 1 0 1380 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_177_11
timestamp 1623621585
transform 1 0 2116 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1670
timestamp 1623621585
transform 1 0 3772 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_177_23
timestamp 1623621585
transform 1 0 3220 0 1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_177_30
timestamp 1623621585
transform 1 0 3864 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_42
timestamp 1623621585
transform 1 0 4968 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_54
timestamp 1623621585
transform 1 0 6072 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_66
timestamp 1623621585
transform 1 0 7176 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_78
timestamp 1623621585
transform 1 0 8280 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1671
timestamp 1623621585
transform 1 0 9016 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_87
timestamp 1623621585
transform 1 0 9108 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_99
timestamp 1623621585
transform 1 0 10212 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_111
timestamp 1623621585
transform 1 0 11316 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_123
timestamp 1623621585
transform 1 0 12420 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1672
timestamp 1623621585
transform 1 0 14260 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_135
timestamp 1623621585
transform 1 0 13524 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_144
timestamp 1623621585
transform 1 0 14352 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_156
timestamp 1623621585
transform 1 0 15456 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_168
timestamp 1623621585
transform 1 0 16560 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_180
timestamp 1623621585
transform 1 0 17664 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1673
timestamp 1623621585
transform 1 0 19504 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_192
timestamp 1623621585
transform 1 0 18768 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_201
timestamp 1623621585
transform 1 0 19596 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0916_
timestamp 1623621585
transform 1 0 21160 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0928_
timestamp 1623621585
transform 1 0 21896 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_177_213
timestamp 1623621585
transform 1 0 20700 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_217
timestamp 1623621585
transform 1 0 21068 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_177_222
timestamp 1623621585
transform 1 0 21528 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_177_230
timestamp 1623621585
transform 1 0 22264 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_242
timestamp 1623621585
transform 1 0 23368 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1674
timestamp 1623621585
transform 1 0 24748 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_177_254
timestamp 1623621585
transform 1 0 24472 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_177_258
timestamp 1623621585
transform 1 0 24840 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_270
timestamp 1623621585
transform 1 0 25944 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_282
timestamp 1623621585
transform 1 0 27048 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_294
timestamp 1623621585
transform 1 0 28152 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_177_306
timestamp 1623621585
transform 1 0 29256 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1675
timestamp 1623621585
transform 1 0 29992 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_177_315
timestamp 1623621585
transform 1 0 30084 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_327
timestamp 1623621585
transform 1 0 31188 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_339
timestamp 1623621585
transform 1 0 32292 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_177_351
timestamp 1623621585
transform 1 0 33396 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1676
timestamp 1623621585
transform 1 0 35236 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_177_363
timestamp 1623621585
transform 1 0 34500 0 1 98464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_177_372
timestamp 1623621585
transform 1 0 35328 0 1 98464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input326
timestamp 1623621585
transform 1 0 37076 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_177_384
timestamp 1623621585
transform 1 0 36432 0 1 98464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_390
timestamp 1623621585
transform 1 0 36984 0 1 98464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_177_395
timestamp 1623621585
transform 1 0 37444 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_355
timestamp 1623621585
transform -1 0 38824 0 1 98464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input325
timestamp 1623621585
transform 1 0 37812 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_177_403
timestamp 1623621585
transform 1 0 38180 0 1 98464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_356
timestamp 1623621585
transform 1 0 1104 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_358
timestamp 1623621585
transform 1 0 1104 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input443
timestamp 1623621585
transform 1 0 1748 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_178_3
timestamp 1623621585
transform 1 0 1380 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_15
timestamp 1623621585
transform 1 0 2484 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_3
timestamp 1623621585
transform 1 0 1380 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_179_11
timestamp 1623621585
transform 1 0 2116 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1684
timestamp 1623621585
transform 1 0 3772 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_27
timestamp 1623621585
transform 1 0 3588 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_39
timestamp 1623621585
transform 1 0 4692 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_23
timestamp 1623621585
transform 1 0 3220 0 1 99552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_179_30
timestamp 1623621585
transform 1 0 3864 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1677
timestamp 1623621585
transform 1 0 6348 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_178_51
timestamp 1623621585
transform 1 0 5796 0 -1 99552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_178_58
timestamp 1623621585
transform 1 0 6440 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_42
timestamp 1623621585
transform 1 0 4968 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_54
timestamp 1623621585
transform 1 0 6072 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_70
timestamp 1623621585
transform 1 0 7544 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_82
timestamp 1623621585
transform 1 0 8648 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_66
timestamp 1623621585
transform 1 0 7176 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_78
timestamp 1623621585
transform 1 0 8280 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1685
timestamp 1623621585
transform 1 0 9016 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_94
timestamp 1623621585
transform 1 0 9752 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_87
timestamp 1623621585
transform 1 0 9108 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_99
timestamp 1623621585
transform 1 0 10212 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1678
timestamp 1623621585
transform 1 0 11592 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_106
timestamp 1623621585
transform 1 0 10856 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_115
timestamp 1623621585
transform 1 0 11684 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_111
timestamp 1623621585
transform 1 0 11316 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_123
timestamp 1623621585
transform 1 0 12420 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_2  _0800_
timestamp 1623621585
transform 1 0 12880 0 -1 99552
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1686
timestamp 1623621585
transform 1 0 14260 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_178_127
timestamp 1623621585
transform 1 0 12788 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_137
timestamp 1623621585
transform 1 0 13708 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_135
timestamp 1623621585
transform 1 0 13524 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_144
timestamp 1623621585
transform 1 0 14352 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_149
timestamp 1623621585
transform 1 0 14812 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_161
timestamp 1623621585
transform 1 0 15916 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_156
timestamp 1623621585
transform 1 0 15456 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1679
timestamp 1623621585
transform 1 0 16836 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_178_169
timestamp 1623621585
transform 1 0 16652 0 -1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_178_172
timestamp 1623621585
transform 1 0 16928 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_184
timestamp 1623621585
transform 1 0 18032 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_168
timestamp 1623621585
transform 1 0 16560 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_180
timestamp 1623621585
transform 1 0 17664 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1687
timestamp 1623621585
transform 1 0 19504 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_196
timestamp 1623621585
transform 1 0 19136 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_208
timestamp 1623621585
transform 1 0 20240 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_192
timestamp 1623621585
transform 1 0 18768 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_179_201
timestamp 1623621585
transform 1 0 19596 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0917_
timestamp 1623621585
transform 1 0 21804 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1680
timestamp 1623621585
transform 1 0 22080 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_220
timestamp 1623621585
transform 1 0 21344 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_229
timestamp 1623621585
transform 1 0 22172 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_213
timestamp 1623621585
transform 1 0 20700 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_229
timestamp 1623621585
transform 1 0 22172 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_241
timestamp 1623621585
transform 1 0 23276 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_241
timestamp 1623621585
transform 1 0 23276 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1688
timestamp 1623621585
transform 1 0 24748 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_253
timestamp 1623621585
transform 1 0 24380 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_265
timestamp 1623621585
transform 1 0 25484 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_253
timestamp 1623621585
transform 1 0 24380 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_179_258
timestamp 1623621585
transform 1 0 24840 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_270
timestamp 1623621585
transform 1 0 25944 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1681
timestamp 1623621585
transform 1 0 27324 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_277
timestamp 1623621585
transform 1 0 26588 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_286
timestamp 1623621585
transform 1 0 27416 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_282
timestamp 1623621585
transform 1 0 27048 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_298
timestamp 1623621585
transform 1 0 28520 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_310
timestamp 1623621585
transform 1 0 29624 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_294
timestamp 1623621585
transform 1 0 28152 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_179_306
timestamp 1623621585
transform 1 0 29256 0 1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1689
timestamp 1623621585
transform 1 0 29992 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_322
timestamp 1623621585
transform 1 0 30728 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_315
timestamp 1623621585
transform 1 0 30084 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_327
timestamp 1623621585
transform 1 0 31188 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_2  _0814_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 33580 0 1 99552
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1682
timestamp 1623621585
transform 1 0 32568 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_178_334
timestamp 1623621585
transform 1 0 31832 0 -1 99552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_178_343
timestamp 1623621585
transform 1 0 32660 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_179_339
timestamp 1623621585
transform 1 0 32292 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_179_351
timestamp 1623621585
transform 1 0 33396 0 1 99552
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _0815_
timestamp 1623621585
transform 1 0 34408 0 1 99552
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1690
timestamp 1623621585
transform 1 0 35236 0 1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_178_355
timestamp 1623621585
transform 1 0 33764 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_178_367
timestamp 1623621585
transform 1 0 34868 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_358
timestamp 1623621585
transform 1 0 34040 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_179_367
timestamp 1623621585
transform 1 0 34868 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_179_372
timestamp 1623621585
transform 1 0 35328 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input327
timestamp 1623621585
transform 1 0 37076 0 -1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_178_379
timestamp 1623621585
transform 1 0 35972 0 -1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_178_395
timestamp 1623621585
transform 1 0 37444 0 -1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_179_384
timestamp 1623621585
transform 1 0 36432 0 1 99552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_357
timestamp 1623621585
transform -1 0 38824 0 -1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_359
timestamp 1623621585
transform -1 0 38824 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1683
timestamp 1623621585
transform 1 0 37812 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input328
timestamp 1623621585
transform 1 0 37812 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_178_400
timestamp 1623621585
transform 1 0 37904 0 -1 99552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_406
timestamp 1623621585
transform 1 0 38456 0 -1 99552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_179_396
timestamp 1623621585
transform 1 0 37536 0 1 99552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_179_403
timestamp 1623621585
transform 1 0 38180 0 1 99552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_360
timestamp 1623621585
transform 1 0 1104 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input444
timestamp 1623621585
transform 1 0 1748 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_180_3
timestamp 1623621585
transform 1 0 1380 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_180_11
timestamp 1623621585
transform 1 0 2116 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_23
timestamp 1623621585
transform 1 0 3220 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_35
timestamp 1623621585
transform 1 0 4324 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1691
timestamp 1623621585
transform 1 0 6348 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_47
timestamp 1623621585
transform 1 0 5428 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_180_55
timestamp 1623621585
transform 1 0 6164 0 -1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_180_58
timestamp 1623621585
transform 1 0 6440 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_70
timestamp 1623621585
transform 1 0 7544 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_82
timestamp 1623621585
transform 1 0 8648 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_94
timestamp 1623621585
transform 1 0 9752 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1692
timestamp 1623621585
transform 1 0 11592 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_106
timestamp 1623621585
transform 1 0 10856 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_115
timestamp 1623621585
transform 1 0 11684 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_127
timestamp 1623621585
transform 1 0 12788 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_139
timestamp 1623621585
transform 1 0 13892 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_151
timestamp 1623621585
transform 1 0 14996 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_163
timestamp 1623621585
transform 1 0 16100 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1693
timestamp 1623621585
transform 1 0 16836 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_180_172
timestamp 1623621585
transform 1 0 16928 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_184
timestamp 1623621585
transform 1 0 18032 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_196
timestamp 1623621585
transform 1 0 19136 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_208
timestamp 1623621585
transform 1 0 20240 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1694
timestamp 1623621585
transform 1 0 22080 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_220
timestamp 1623621585
transform 1 0 21344 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_180_229
timestamp 1623621585
transform 1 0 22172 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0919_
timestamp 1623621585
transform 1 0 22908 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_180_241
timestamp 1623621585
transform 1 0 23276 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_253
timestamp 1623621585
transform 1 0 24380 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_265
timestamp 1623621585
transform 1 0 25484 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1695
timestamp 1623621585
transform 1 0 27324 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_277
timestamp 1623621585
transform 1 0 26588 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_286
timestamp 1623621585
transform 1 0 27416 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_298
timestamp 1623621585
transform 1 0 28520 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_310
timestamp 1623621585
transform 1 0 29624 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_322
timestamp 1623621585
transform 1 0 30728 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1696
timestamp 1623621585
transform 1 0 32568 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_180_334
timestamp 1623621585
transform 1 0 31832 0 -1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_180_343
timestamp 1623621585
transform 1 0 32660 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_355
timestamp 1623621585
transform 1 0 33764 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_180_367
timestamp 1623621585
transform 1 0 34868 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input329
timestamp 1623621585
transform 1 0 37076 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_180_379
timestamp 1623621585
transform 1 0 35972 0 -1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_180_395
timestamp 1623621585
transform 1 0 37444 0 -1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_361
timestamp 1623621585
transform -1 0 38824 0 -1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1697
timestamp 1623621585
transform 1 0 37812 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_180_400
timestamp 1623621585
transform 1 0 37904 0 -1 100640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_406
timestamp 1623621585
transform 1 0 38456 0 -1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_362
timestamp 1623621585
transform 1 0 1104 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_181_3
timestamp 1623621585
transform 1 0 1380 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_15
timestamp 1623621585
transform 1 0 2484 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1698
timestamp 1623621585
transform 1 0 3772 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_181_27
timestamp 1623621585
transform 1 0 3588 0 1 100640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_181_30
timestamp 1623621585
transform 1 0 3864 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_42
timestamp 1623621585
transform 1 0 4968 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_54
timestamp 1623621585
transform 1 0 6072 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_66
timestamp 1623621585
transform 1 0 7176 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_78
timestamp 1623621585
transform 1 0 8280 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1699
timestamp 1623621585
transform 1 0 9016 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_87
timestamp 1623621585
transform 1 0 9108 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_99
timestamp 1623621585
transform 1 0 10212 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_111
timestamp 1623621585
transform 1 0 11316 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_123
timestamp 1623621585
transform 1 0 12420 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1700
timestamp 1623621585
transform 1 0 14260 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_135
timestamp 1623621585
transform 1 0 13524 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_144
timestamp 1623621585
transform 1 0 14352 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_156
timestamp 1623621585
transform 1 0 15456 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_168
timestamp 1623621585
transform 1 0 16560 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_180
timestamp 1623621585
transform 1 0 17664 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1701
timestamp 1623621585
transform 1 0 19504 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_192
timestamp 1623621585
transform 1 0 18768 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_201
timestamp 1623621585
transform 1 0 19596 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_213
timestamp 1623621585
transform 1 0 20700 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_225
timestamp 1623621585
transform 1 0 21804 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_237
timestamp 1623621585
transform 1 0 22908 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_249
timestamp 1623621585
transform 1 0 24012 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1702
timestamp 1623621585
transform 1 0 24748 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_258
timestamp 1623621585
transform 1 0 24840 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_270
timestamp 1623621585
transform 1 0 25944 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_282
timestamp 1623621585
transform 1 0 27048 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_294
timestamp 1623621585
transform 1 0 28152 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_181_306
timestamp 1623621585
transform 1 0 29256 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1703
timestamp 1623621585
transform 1 0 29992 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_181_315
timestamp 1623621585
transform 1 0 30084 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_327
timestamp 1623621585
transform 1 0 31188 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_339
timestamp 1623621585
transform 1 0 32292 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_181_351
timestamp 1623621585
transform 1 0 33396 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1704
timestamp 1623621585
transform 1 0 35236 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_181_363
timestamp 1623621585
transform 1 0 34500 0 1 100640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_181_372
timestamp 1623621585
transform 1 0 35328 0 1 100640
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input330
timestamp 1623621585
transform 1 0 37076 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_181_384
timestamp 1623621585
transform 1 0 36432 0 1 100640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_390
timestamp 1623621585
transform 1 0 36984 0 1 100640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_181_395
timestamp 1623621585
transform 1 0 37444 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_363
timestamp 1623621585
transform -1 0 38824 0 1 100640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input300
timestamp 1623621585
transform 1 0 37812 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_181_403
timestamp 1623621585
transform 1 0 38180 0 1 100640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_364
timestamp 1623621585
transform 1 0 1104 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input445
timestamp 1623621585
transform 1 0 1748 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_182_3
timestamp 1623621585
transform 1 0 1380 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_11
timestamp 1623621585
transform 1 0 2116 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_23
timestamp 1623621585
transform 1 0 3220 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_35
timestamp 1623621585
transform 1 0 4324 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0925_
timestamp 1623621585
transform 1 0 5704 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1705
timestamp 1623621585
transform 1 0 6348 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_182_47
timestamp 1623621585
transform 1 0 5428 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_182_53
timestamp 1623621585
transform 1 0 5980 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_58
timestamp 1623621585
transform 1 0 6440 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_70
timestamp 1623621585
transform 1 0 7544 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_82
timestamp 1623621585
transform 1 0 8648 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_94
timestamp 1623621585
transform 1 0 9752 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _0798_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623621585
transform 1 0 12052 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1706
timestamp 1623621585
transform 1 0 11592 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_106
timestamp 1623621585
transform 1 0 10856 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_182_115
timestamp 1623621585
transform 1 0 11684 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_127
timestamp 1623621585
transform 1 0 12788 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_139
timestamp 1623621585
transform 1 0 13892 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_151
timestamp 1623621585
transform 1 0 14996 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_163
timestamp 1623621585
transform 1 0 16100 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1707
timestamp 1623621585
transform 1 0 16836 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_182_172
timestamp 1623621585
transform 1 0 16928 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_184
timestamp 1623621585
transform 1 0 18032 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_196
timestamp 1623621585
transform 1 0 19136 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_208
timestamp 1623621585
transform 1 0 20240 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1708
timestamp 1623621585
transform 1 0 22080 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_220
timestamp 1623621585
transform 1 0 21344 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_182_229
timestamp 1623621585
transform 1 0 22172 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0931_
timestamp 1623621585
transform 1 0 23092 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_182_237
timestamp 1623621585
transform 1 0 22908 0 -1 101728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_182_243
timestamp 1623621585
transform 1 0 23460 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_255
timestamp 1623621585
transform 1 0 24564 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_267
timestamp 1623621585
transform 1 0 25668 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1709
timestamp 1623621585
transform 1 0 27324 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_182_279
timestamp 1623621585
transform 1 0 26772 0 -1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_182_286
timestamp 1623621585
transform 1 0 27416 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_298
timestamp 1623621585
transform 1 0 28520 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_310
timestamp 1623621585
transform 1 0 29624 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_322
timestamp 1623621585
transform 1 0 30728 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1710
timestamp 1623621585
transform 1 0 32568 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_334
timestamp 1623621585
transform 1 0 31832 0 -1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_182_343
timestamp 1623621585
transform 1 0 32660 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_355
timestamp 1623621585
transform 1 0 33764 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_182_367
timestamp 1623621585
transform 1 0 34868 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input301
timestamp 1623621585
transform 1 0 37076 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_182_379
timestamp 1623621585
transform 1 0 35972 0 -1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_395
timestamp 1623621585
transform 1 0 37444 0 -1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_365
timestamp 1623621585
transform -1 0 38824 0 -1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1711
timestamp 1623621585
transform 1 0 37812 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_182_400
timestamp 1623621585
transform 1 0 37904 0 -1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_182_406
timestamp 1623621585
transform 1 0 38456 0 -1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_366
timestamp 1623621585
transform 1 0 1104 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input446
timestamp 1623621585
transform 1 0 1748 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_183_3
timestamp 1623621585
transform 1 0 1380 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_183_11
timestamp 1623621585
transform 1 0 2116 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1712
timestamp 1623621585
transform 1 0 3772 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_183_23
timestamp 1623621585
transform 1 0 3220 0 1 101728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_183_30
timestamp 1623621585
transform 1 0 3864 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_42
timestamp 1623621585
transform 1 0 4968 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_54
timestamp 1623621585
transform 1 0 6072 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_66
timestamp 1623621585
transform 1 0 7176 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_78
timestamp 1623621585
transform 1 0 8280 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1713
timestamp 1623621585
transform 1 0 9016 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_87
timestamp 1623621585
transform 1 0 9108 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_99
timestamp 1623621585
transform 1 0 10212 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0786_
timestamp 1623621585
transform 1 0 11224 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_183_107
timestamp 1623621585
transform 1 0 10948 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_183_118
timestamp 1623621585
transform 1 0 11960 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0788_
timestamp 1623621585
transform 1 0 12788 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1714
timestamp 1623621585
transform 1 0 14260 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_183_126
timestamp 1623621585
transform 1 0 12696 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_135
timestamp 1623621585
transform 1 0 13524 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_144
timestamp 1623621585
transform 1 0 14352 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_156
timestamp 1623621585
transform 1 0 15456 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_168
timestamp 1623621585
transform 1 0 16560 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_180
timestamp 1623621585
transform 1 0 17664 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1715
timestamp 1623621585
transform 1 0 19504 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_192
timestamp 1623621585
transform 1 0 18768 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_201
timestamp 1623621585
transform 1 0 19596 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_213
timestamp 1623621585
transform 1 0 20700 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_225
timestamp 1623621585
transform 1 0 21804 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_237
timestamp 1623621585
transform 1 0 22908 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_249
timestamp 1623621585
transform 1 0 24012 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1716
timestamp 1623621585
transform 1 0 24748 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_258
timestamp 1623621585
transform 1 0 24840 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_270
timestamp 1623621585
transform 1 0 25944 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_282
timestamp 1623621585
transform 1 0 27048 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_294
timestamp 1623621585
transform 1 0 28152 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_183_306
timestamp 1623621585
transform 1 0 29256 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1717
timestamp 1623621585
transform 1 0 29992 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_183_315
timestamp 1623621585
transform 1 0 30084 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_327
timestamp 1623621585
transform 1 0 31188 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_339
timestamp 1623621585
transform 1 0 32292 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_351
timestamp 1623621585
transform 1 0 33396 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1718
timestamp 1623621585
transform 1 0 35236 0 1 101728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_183_363
timestamp 1623621585
transform 1 0 34500 0 1 101728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_183_372
timestamp 1623621585
transform 1 0 35328 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_183_384
timestamp 1623621585
transform 1 0 36432 0 1 101728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_367
timestamp 1623621585
transform -1 0 38824 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input302
timestamp 1623621585
transform 1 0 37812 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_183_396
timestamp 1623621585
transform 1 0 37536 0 1 101728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_183_403
timestamp 1623621585
transform 1 0 38180 0 1 101728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_368
timestamp 1623621585
transform 1 0 1104 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_184_3
timestamp 1623621585
transform 1 0 1380 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_15
timestamp 1623621585
transform 1 0 2484 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_27
timestamp 1623621585
transform 1 0 3588 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_39
timestamp 1623621585
transform 1 0 4692 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1719
timestamp 1623621585
transform 1 0 6348 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_184_51
timestamp 1623621585
transform 1 0 5796 0 -1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_184_58
timestamp 1623621585
transform 1 0 6440 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1623621585
transform 1 0 7636 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_184_70
timestamp 1623621585
transform 1 0 7544 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_74
timestamp 1623621585
transform 1 0 7912 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_86
timestamp 1623621585
transform 1 0 9016 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_98
timestamp 1623621585
transform 1 0 10120 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _0790_
timestamp 1623621585
transform 1 0 12052 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1720
timestamp 1623621585
transform 1 0 11592 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_184_110
timestamp 1623621585
transform 1 0 11224 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_184_115
timestamp 1623621585
transform 1 0 11684 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_127
timestamp 1623621585
transform 1 0 12788 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_139
timestamp 1623621585
transform 1 0 13892 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_151
timestamp 1623621585
transform 1 0 14996 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_184_163
timestamp 1623621585
transform 1 0 16100 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1721
timestamp 1623621585
transform 1 0 16836 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_184_172
timestamp 1623621585
transform 1 0 16928 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_184
timestamp 1623621585
transform 1 0 18032 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_196
timestamp 1623621585
transform 1 0 19136 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_208
timestamp 1623621585
transform 1 0 20240 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1722
timestamp 1623621585
transform 1 0 22080 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_220
timestamp 1623621585
transform 1 0 21344 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_184_229
timestamp 1623621585
transform 1 0 22172 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_241
timestamp 1623621585
transform 1 0 23276 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_253
timestamp 1623621585
transform 1 0 24380 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_265
timestamp 1623621585
transform 1 0 25484 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0927_
timestamp 1623621585
transform 1 0 26588 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1723
timestamp 1623621585
transform 1 0 27324 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_184_281
timestamp 1623621585
transform 1 0 26956 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_286
timestamp 1623621585
transform 1 0 27416 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_298
timestamp 1623621585
transform 1 0 28520 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_310
timestamp 1623621585
transform 1 0 29624 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_322
timestamp 1623621585
transform 1 0 30728 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1724
timestamp 1623621585
transform 1 0 32568 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_184_334
timestamp 1623621585
transform 1 0 31832 0 -1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_184_343
timestamp 1623621585
transform 1 0 32660 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_355
timestamp 1623621585
transform 1 0 33764 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_184_367
timestamp 1623621585
transform 1 0 34868 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input303
timestamp 1623621585
transform 1 0 37076 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_184_379
timestamp 1623621585
transform 1 0 35972 0 -1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_184_395
timestamp 1623621585
transform 1 0 37444 0 -1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_369
timestamp 1623621585
transform -1 0 38824 0 -1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1725
timestamp 1623621585
transform 1 0 37812 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_184_400
timestamp 1623621585
transform 1 0 37904 0 -1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_184_406
timestamp 1623621585
transform 1 0 38456 0 -1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_370
timestamp 1623621585
transform 1 0 1104 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_372
timestamp 1623621585
transform 1 0 1104 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input447
timestamp 1623621585
transform 1 0 1748 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input448
timestamp 1623621585
transform 1 0 1748 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_185_3
timestamp 1623621585
transform 1 0 1380 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_185_11
timestamp 1623621585
transform 1 0 2116 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_3
timestamp 1623621585
transform 1 0 1380 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_11
timestamp 1623621585
transform 1 0 2116 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1726
timestamp 1623621585
transform 1 0 3772 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_185_23
timestamp 1623621585
transform 1 0 3220 0 1 102816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_185_30
timestamp 1623621585
transform 1 0 3864 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_23
timestamp 1623621585
transform 1 0 3220 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_35
timestamp 1623621585
transform 1 0 4324 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1623621585
transform 1 0 6164 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0939_
timestamp 1623621585
transform 1 0 6808 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1733
timestamp 1623621585
transform 1 0 6348 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_42
timestamp 1623621585
transform 1 0 4968 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_185_54
timestamp 1623621585
transform 1 0 6072 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_185_58
timestamp 1623621585
transform 1 0 6440 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_186_47
timestamp 1623621585
transform 1 0 5428 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_186_55
timestamp 1623621585
transform 1 0 6164 0 -1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_186_58
timestamp 1623621585
transform 1 0 6440 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_65
timestamp 1623621585
transform 1 0 7084 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_77
timestamp 1623621585
transform 1 0 8188 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_70
timestamp 1623621585
transform 1 0 7544 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_82
timestamp 1623621585
transform 1 0 8648 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1727
timestamp 1623621585
transform 1 0 9016 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_185_85
timestamp 1623621585
transform 1 0 8924 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_87
timestamp 1623621585
transform 1 0 9108 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_99
timestamp 1623621585
transform 1 0 10212 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_94
timestamp 1623621585
transform 1 0 9752 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _0794_
timestamp 1623621585
transform 1 0 12420 0 -1 103904
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1734
timestamp 1623621585
transform 1 0 11592 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_111
timestamp 1623621585
transform 1 0 11316 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_123
timestamp 1623621585
transform 1 0 12420 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_106
timestamp 1623621585
transform 1 0 10856 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_186_115
timestamp 1623621585
transform 1 0 11684 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1728
timestamp 1623621585
transform 1 0 14260 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_185_135
timestamp 1623621585
transform 1 0 13524 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_144
timestamp 1623621585
transform 1 0 14352 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_136
timestamp 1623621585
transform 1 0 13616 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_156
timestamp 1623621585
transform 1 0 15456 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_148
timestamp 1623621585
transform 1 0 14720 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_160
timestamp 1623621585
transform 1 0 15824 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1735
timestamp 1623621585
transform 1 0 16836 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_168
timestamp 1623621585
transform 1 0 16560 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_180
timestamp 1623621585
transform 1 0 17664 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_186_168
timestamp 1623621585
transform 1 0 16560 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_186_172
timestamp 1623621585
transform 1 0 16928 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_184
timestamp 1623621585
transform 1 0 18032 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1729
timestamp 1623621585
transform 1 0 19504 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_185_192
timestamp 1623621585
transform 1 0 18768 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_201
timestamp 1623621585
transform 1 0 19596 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_196
timestamp 1623621585
transform 1 0 19136 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_208
timestamp 1623621585
transform 1 0 20240 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0791_
timestamp 1623621585
transform 1 0 20976 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1736
timestamp 1623621585
transform 1 0 22080 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_213
timestamp 1623621585
transform 1 0 20700 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_225
timestamp 1623621585
transform 1 0 21804 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_224
timestamp 1623621585
transform 1 0 21712 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_186_229
timestamp 1623621585
transform 1 0 22172 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_237
timestamp 1623621585
transform 1 0 22908 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_185_249
timestamp 1623621585
transform 1 0 24012 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_241
timestamp 1623621585
transform 1 0 23276 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1623621585
transform 1 0 24840 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1730
timestamp 1623621585
transform 1 0 24748 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_258
timestamp 1623621585
transform 1 0 24840 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_185_270
timestamp 1623621585
transform 1 0 25944 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_186_253
timestamp 1623621585
transform 1 0 24380 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_186_257
timestamp 1623621585
transform 1 0 24748 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_262
timestamp 1623621585
transform 1 0 25208 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0938_
timestamp 1623621585
transform 1 0 26312 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1737
timestamp 1623621585
transform 1 0 27324 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_278
timestamp 1623621585
transform 1 0 26680 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_290
timestamp 1623621585
transform 1 0 27784 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_274
timestamp 1623621585
transform 1 0 26312 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_186_282
timestamp 1623621585
transform 1 0 27048 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_186_286
timestamp 1623621585
transform 1 0 27416 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_302
timestamp 1623621585
transform 1 0 28888 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_298
timestamp 1623621585
transform 1 0 28520 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_310
timestamp 1623621585
transform 1 0 29624 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1731
timestamp 1623621585
transform 1 0 29992 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_315
timestamp 1623621585
transform 1 0 30084 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_327
timestamp 1623621585
transform 1 0 31188 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_322
timestamp 1623621585
transform 1 0 30728 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1738
timestamp 1623621585
transform 1 0 32568 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_185_339
timestamp 1623621585
transform 1 0 32292 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_185_351
timestamp 1623621585
transform 1 0 33396 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_186_334
timestamp 1623621585
transform 1 0 31832 0 -1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_186_343
timestamp 1623621585
transform 1 0 32660 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1732
timestamp 1623621585
transform 1 0 35236 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_185_363
timestamp 1623621585
transform 1 0 34500 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_185_372
timestamp 1623621585
transform 1 0 35328 0 1 102816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_355
timestamp 1623621585
transform 1 0 33764 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_186_367
timestamp 1623621585
transform 1 0 34868 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input304
timestamp 1623621585
transform 1 0 37260 0 1 102816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input305
timestamp 1623621585
transform 1 0 37076 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_185_384
timestamp 1623621585
transform 1 0 36432 0 1 102816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_185_392
timestamp 1623621585
transform 1 0 37168 0 1 102816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_186_379
timestamp 1623621585
transform 1 0 35972 0 -1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_186_395
timestamp 1623621585
transform 1 0 37444 0 -1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_371
timestamp 1623621585
transform -1 0 38824 0 1 102816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_373
timestamp 1623621585
transform -1 0 38824 0 -1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1739
timestamp 1623621585
transform 1 0 37812 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_185_403
timestamp 1623621585
transform 1 0 38180 0 1 102816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_186_400
timestamp 1623621585
transform 1 0 37904 0 -1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_186_406
timestamp 1623621585
transform 1 0 38456 0 -1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_374
timestamp 1623621585
transform 1 0 1104 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_187_3
timestamp 1623621585
transform 1 0 1380 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_15
timestamp 1623621585
transform 1 0 2484 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1740
timestamp 1623621585
transform 1 0 3772 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_187_27
timestamp 1623621585
transform 1 0 3588 0 1 103904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_187_30
timestamp 1623621585
transform 1 0 3864 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_42
timestamp 1623621585
transform 1 0 4968 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_54
timestamp 1623621585
transform 1 0 6072 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_66
timestamp 1623621585
transform 1 0 7176 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_78
timestamp 1623621585
transform 1 0 8280 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1741
timestamp 1623621585
transform 1 0 9016 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_87
timestamp 1623621585
transform 1 0 9108 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_99
timestamp 1623621585
transform 1 0 10212 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_111
timestamp 1623621585
transform 1 0 11316 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_123
timestamp 1623621585
transform 1 0 12420 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1742
timestamp 1623621585
transform 1 0 14260 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_187_135
timestamp 1623621585
transform 1 0 13524 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_187_144
timestamp 1623621585
transform 1 0 14352 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_156
timestamp 1623621585
transform 1 0 15456 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_168
timestamp 1623621585
transform 1 0 16560 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_180
timestamp 1623621585
transform 1 0 17664 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1743
timestamp 1623621585
transform 1 0 19504 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_187_192
timestamp 1623621585
transform 1 0 18768 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_187_201
timestamp 1623621585
transform 1 0 19596 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_213
timestamp 1623621585
transform 1 0 20700 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_225
timestamp 1623621585
transform 1 0 21804 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_237
timestamp 1623621585
transform 1 0 22908 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_187_249
timestamp 1623621585
transform 1 0 24012 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1744
timestamp 1623621585
transform 1 0 24748 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_258
timestamp 1623621585
transform 1 0 24840 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_270
timestamp 1623621585
transform 1 0 25944 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_282
timestamp 1623621585
transform 1 0 27048 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1623621585
transform 1 0 29348 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_187_294
timestamp 1623621585
transform 1 0 28152 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_187_306
timestamp 1623621585
transform 1 0 29256 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_187_310
timestamp 1623621585
transform 1 0 29624 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1745
timestamp 1623621585
transform 1 0 29992 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_187_315
timestamp 1623621585
transform 1 0 30084 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_327
timestamp 1623621585
transform 1 0 31188 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_339
timestamp 1623621585
transform 1 0 32292 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_187_351
timestamp 1623621585
transform 1 0 33396 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1746
timestamp 1623621585
transform 1 0 35236 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_187_363
timestamp 1623621585
transform 1 0 34500 0 1 103904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_187_372
timestamp 1623621585
transform 1 0 35328 0 1 103904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input307
timestamp 1623621585
transform 1 0 37076 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_187_384
timestamp 1623621585
transform 1 0 36432 0 1 103904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_187_390
timestamp 1623621585
transform 1 0 36984 0 1 103904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_187_395
timestamp 1623621585
transform 1 0 37444 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_375
timestamp 1623621585
transform -1 0 38824 0 1 103904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input306
timestamp 1623621585
transform 1 0 37812 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_187_403
timestamp 1623621585
transform 1 0 38180 0 1 103904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_376
timestamp 1623621585
transform 1 0 1104 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input450
timestamp 1623621585
transform 1 0 1748 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_188_3
timestamp 1623621585
transform 1 0 1380 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_188_11
timestamp 1623621585
transform 1 0 2116 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_23
timestamp 1623621585
transform 1 0 3220 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_35
timestamp 1623621585
transform 1 0 4324 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1747
timestamp 1623621585
transform 1 0 6348 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_47
timestamp 1623621585
transform 1 0 5428 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_188_55
timestamp 1623621585
transform 1 0 6164 0 -1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_188_58
timestamp 1623621585
transform 1 0 6440 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_70
timestamp 1623621585
transform 1 0 7544 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_82
timestamp 1623621585
transform 1 0 8648 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_94
timestamp 1623621585
transform 1 0 9752 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1748
timestamp 1623621585
transform 1 0 11592 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_106
timestamp 1623621585
transform 1 0 10856 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_115
timestamp 1623621585
transform 1 0 11684 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_127
timestamp 1623621585
transform 1 0 12788 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_139
timestamp 1623621585
transform 1 0 13892 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_151
timestamp 1623621585
transform 1 0 14996 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_188_163
timestamp 1623621585
transform 1 0 16100 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1749
timestamp 1623621585
transform 1 0 16836 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_172
timestamp 1623621585
transform 1 0 16928 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_184
timestamp 1623621585
transform 1 0 18032 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_196
timestamp 1623621585
transform 1 0 19136 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_208
timestamp 1623621585
transform 1 0 20240 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1750
timestamp 1623621585
transform 1 0 22080 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_220
timestamp 1623621585
transform 1 0 21344 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_229
timestamp 1623621585
transform 1 0 22172 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_241
timestamp 1623621585
transform 1 0 23276 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _0793_
timestamp 1623621585
transform 1 0 24840 0 -1 104992
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_188_253
timestamp 1623621585
transform 1 0 24380 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_188_257
timestamp 1623621585
transform 1 0 24748 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1751
timestamp 1623621585
transform 1 0 27324 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_188_271
timestamp 1623621585
transform 1 0 26036 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_188_283
timestamp 1623621585
transform 1 0 27140 0 -1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_188_286
timestamp 1623621585
transform 1 0 27416 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_298
timestamp 1623621585
transform 1 0 28520 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_310
timestamp 1623621585
transform 1 0 29624 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_322
timestamp 1623621585
transform 1 0 30728 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1752
timestamp 1623621585
transform 1 0 32568 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_188_334
timestamp 1623621585
transform 1 0 31832 0 -1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_188_343
timestamp 1623621585
transform 1 0 32660 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_355
timestamp 1623621585
transform 1 0 33764 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_188_367
timestamp 1623621585
transform 1 0 34868 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input308
timestamp 1623621585
transform 1 0 37076 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_188_379
timestamp 1623621585
transform 1 0 35972 0 -1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_188_395
timestamp 1623621585
transform 1 0 37444 0 -1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_377
timestamp 1623621585
transform -1 0 38824 0 -1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1753
timestamp 1623621585
transform 1 0 37812 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_188_400
timestamp 1623621585
transform 1 0 37904 0 -1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_188_406
timestamp 1623621585
transform 1 0 38456 0 -1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_378
timestamp 1623621585
transform 1 0 1104 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input451
timestamp 1623621585
transform 1 0 1380 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_189_7
timestamp 1623621585
transform 1 0 1748 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_19
timestamp 1623621585
transform 1 0 2852 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1754
timestamp 1623621585
transform 1 0 3772 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_189_27
timestamp 1623621585
transform 1 0 3588 0 1 104992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_189_30
timestamp 1623621585
transform 1 0 3864 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_42
timestamp 1623621585
transform 1 0 4968 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_54
timestamp 1623621585
transform 1 0 6072 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_66
timestamp 1623621585
transform 1 0 7176 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_78
timestamp 1623621585
transform 1 0 8280 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1755
timestamp 1623621585
transform 1 0 9016 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_87
timestamp 1623621585
transform 1 0 9108 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_99
timestamp 1623621585
transform 1 0 10212 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_111
timestamp 1623621585
transform 1 0 11316 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_123
timestamp 1623621585
transform 1 0 12420 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1756
timestamp 1623621585
transform 1 0 14260 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_135
timestamp 1623621585
transform 1 0 13524 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_144
timestamp 1623621585
transform 1 0 14352 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_156
timestamp 1623621585
transform 1 0 15456 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_168
timestamp 1623621585
transform 1 0 16560 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_180
timestamp 1623621585
transform 1 0 17664 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1757
timestamp 1623621585
transform 1 0 19504 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_192
timestamp 1623621585
transform 1 0 18768 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_201
timestamp 1623621585
transform 1 0 19596 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_213
timestamp 1623621585
transform 1 0 20700 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_225
timestamp 1623621585
transform 1 0 21804 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_237
timestamp 1623621585
transform 1 0 22908 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_249
timestamp 1623621585
transform 1 0 24012 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _0795_
timestamp 1623621585
transform 1 0 25208 0 1 104992
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1758
timestamp 1623621585
transform 1 0 24748 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_189_258
timestamp 1623621585
transform 1 0 24840 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_189_275
timestamp 1623621585
transform 1 0 26404 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_287
timestamp 1623621585
transform 1 0 27508 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_299
timestamp 1623621585
transform 1 0 28612 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_189_311
timestamp 1623621585
transform 1 0 29716 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1759
timestamp 1623621585
transform 1 0 29992 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_315
timestamp 1623621585
transform 1 0 30084 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_189_327
timestamp 1623621585
transform 1 0 31188 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1623621585
transform 1 0 32016 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_189_335
timestamp 1623621585
transform 1 0 31924 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_189_339
timestamp 1623621585
transform 1 0 32292 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_189_351
timestamp 1623621585
transform 1 0 33396 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1760
timestamp 1623621585
transform 1 0 35236 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_189_363
timestamp 1623621585
transform 1 0 34500 0 1 104992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_189_372
timestamp 1623621585
transform 1 0 35328 0 1 104992
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input311
timestamp 1623621585
transform 1 0 37076 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_189_384
timestamp 1623621585
transform 1 0 36432 0 1 104992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_189_390
timestamp 1623621585
transform 1 0 36984 0 1 104992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_189_395
timestamp 1623621585
transform 1 0 37444 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_379
timestamp 1623621585
transform -1 0 38824 0 1 104992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input309
timestamp 1623621585
transform 1 0 37812 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_189_403
timestamp 1623621585
transform 1 0 38180 0 1 104992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_380
timestamp 1623621585
transform 1 0 1104 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_190_3
timestamp 1623621585
transform 1 0 1380 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_15
timestamp 1623621585
transform 1 0 2484 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_27
timestamp 1623621585
transform 1 0 3588 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_39
timestamp 1623621585
transform 1 0 4692 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1761
timestamp 1623621585
transform 1 0 6348 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_190_51
timestamp 1623621585
transform 1 0 5796 0 -1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_190_58
timestamp 1623621585
transform 1 0 6440 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_70
timestamp 1623621585
transform 1 0 7544 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_82
timestamp 1623621585
transform 1 0 8648 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_94
timestamp 1623621585
transform 1 0 9752 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1762
timestamp 1623621585
transform 1 0 11592 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_106
timestamp 1623621585
transform 1 0 10856 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_115
timestamp 1623621585
transform 1 0 11684 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_127
timestamp 1623621585
transform 1 0 12788 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_139
timestamp 1623621585
transform 1 0 13892 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_151
timestamp 1623621585
transform 1 0 14996 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_190_163
timestamp 1623621585
transform 1 0 16100 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1763
timestamp 1623621585
transform 1 0 16836 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_190_172
timestamp 1623621585
transform 1 0 16928 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_184
timestamp 1623621585
transform 1 0 18032 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_196
timestamp 1623621585
transform 1 0 19136 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_208
timestamp 1623621585
transform 1 0 20240 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1764
timestamp 1623621585
transform 1 0 22080 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_220
timestamp 1623621585
transform 1 0 21344 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_229
timestamp 1623621585
transform 1 0 22172 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_241
timestamp 1623621585
transform 1 0 23276 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_253
timestamp 1623621585
transform 1 0 24380 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_265
timestamp 1623621585
transform 1 0 25484 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1765
timestamp 1623621585
transform 1 0 27324 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_277
timestamp 1623621585
transform 1 0 26588 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_286
timestamp 1623621585
transform 1 0 27416 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_298
timestamp 1623621585
transform 1 0 28520 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_310
timestamp 1623621585
transform 1 0 29624 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_322
timestamp 1623621585
transform 1 0 30728 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1766
timestamp 1623621585
transform 1 0 32568 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_190_334
timestamp 1623621585
transform 1 0 31832 0 -1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_190_343
timestamp 1623621585
transform 1 0 32660 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_355
timestamp 1623621585
transform 1 0 33764 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_190_367
timestamp 1623621585
transform 1 0 34868 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input312
timestamp 1623621585
transform 1 0 37076 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_190_379
timestamp 1623621585
transform 1 0 35972 0 -1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_190_395
timestamp 1623621585
transform 1 0 37444 0 -1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_381
timestamp 1623621585
transform -1 0 38824 0 -1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1767
timestamp 1623621585
transform 1 0 37812 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_190_400
timestamp 1623621585
transform 1 0 37904 0 -1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_190_406
timestamp 1623621585
transform 1 0 38456 0 -1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_382
timestamp 1623621585
transform 1 0 1104 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_384
timestamp 1623621585
transform 1 0 1104 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output647
timestamp 1623621585
transform -1 0 2116 0 1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output660
timestamp 1623621585
transform 1 0 1748 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  INSDIODE2_1
timestamp 1623621585
transform -1 0 1748 0 1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_191_3
timestamp 1623621585
transform 1 0 1380 0 1 106080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_191_11
timestamp 1623621585
transform 1 0 2116 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_3
timestamp 1623621585
transform 1 0 1380 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_192_11
timestamp 1623621585
transform 1 0 2116 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1768
timestamp 1623621585
transform 1 0 3772 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_191_23
timestamp 1623621585
transform 1 0 3220 0 1 106080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_191_30
timestamp 1623621585
transform 1 0 3864 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_23
timestamp 1623621585
transform 1 0 3220 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_35
timestamp 1623621585
transform 1 0 4324 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1775
timestamp 1623621585
transform 1 0 6348 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_42
timestamp 1623621585
transform 1 0 4968 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_54
timestamp 1623621585
transform 1 0 6072 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_47
timestamp 1623621585
transform 1 0 5428 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_192_55
timestamp 1623621585
transform 1 0 6164 0 -1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_192_58
timestamp 1623621585
transform 1 0 6440 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_66
timestamp 1623621585
transform 1 0 7176 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_78
timestamp 1623621585
transform 1 0 8280 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_70
timestamp 1623621585
transform 1 0 7544 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_82
timestamp 1623621585
transform 1 0 8648 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1769
timestamp 1623621585
transform 1 0 9016 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_87
timestamp 1623621585
transform 1 0 9108 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_99
timestamp 1623621585
transform 1 0 10212 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_94
timestamp 1623621585
transform 1 0 9752 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1776
timestamp 1623621585
transform 1 0 11592 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_111
timestamp 1623621585
transform 1 0 11316 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_123
timestamp 1623621585
transform 1 0 12420 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_106
timestamp 1623621585
transform 1 0 10856 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_115
timestamp 1623621585
transform 1 0 11684 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1770
timestamp 1623621585
transform 1 0 14260 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_135
timestamp 1623621585
transform 1 0 13524 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_144
timestamp 1623621585
transform 1 0 14352 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_127
timestamp 1623621585
transform 1 0 12788 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_139
timestamp 1623621585
transform 1 0 13892 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_156
timestamp 1623621585
transform 1 0 15456 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_151
timestamp 1623621585
transform 1 0 14996 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_163
timestamp 1623621585
transform 1 0 16100 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1777
timestamp 1623621585
transform 1 0 16836 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_168
timestamp 1623621585
transform 1 0 16560 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_180
timestamp 1623621585
transform 1 0 17664 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_172
timestamp 1623621585
transform 1 0 16928 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_184
timestamp 1623621585
transform 1 0 18032 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1771
timestamp 1623621585
transform 1 0 19504 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_192
timestamp 1623621585
transform 1 0 18768 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_201
timestamp 1623621585
transform 1 0 19596 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_196
timestamp 1623621585
transform 1 0 19136 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_208
timestamp 1623621585
transform 1 0 20240 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1778
timestamp 1623621585
transform 1 0 22080 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_213
timestamp 1623621585
transform 1 0 20700 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_225
timestamp 1623621585
transform 1 0 21804 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_220
timestamp 1623621585
transform 1 0 21344 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_229
timestamp 1623621585
transform 1 0 22172 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_237
timestamp 1623621585
transform 1 0 22908 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_249
timestamp 1623621585
transform 1 0 24012 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_241
timestamp 1623621585
transform 1 0 23276 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1772
timestamp 1623621585
transform 1 0 24748 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_258
timestamp 1623621585
transform 1 0 24840 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_270
timestamp 1623621585
transform 1 0 25944 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_253
timestamp 1623621585
transform 1 0 24380 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_265
timestamp 1623621585
transform 1 0 25484 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1779
timestamp 1623621585
transform 1 0 27324 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_282
timestamp 1623621585
transform 1 0 27048 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_277
timestamp 1623621585
transform 1 0 26588 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_286
timestamp 1623621585
transform 1 0 27416 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_294
timestamp 1623621585
transform 1 0 28152 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_191_306
timestamp 1623621585
transform 1 0 29256 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_298
timestamp 1623621585
transform 1 0 28520 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_310
timestamp 1623621585
transform 1 0 29624 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1773
timestamp 1623621585
transform 1 0 29992 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_315
timestamp 1623621585
transform 1 0 30084 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_327
timestamp 1623621585
transform 1 0 31188 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_322
timestamp 1623621585
transform 1 0 30728 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1780
timestamp 1623621585
transform 1 0 32568 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_191_339
timestamp 1623621585
transform 1 0 32292 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_191_351
timestamp 1623621585
transform 1 0 33396 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_192_334
timestamp 1623621585
transform 1 0 31832 0 -1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_192_343
timestamp 1623621585
transform 1 0 32660 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1774
timestamp 1623621585
transform 1 0 35236 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_191_363
timestamp 1623621585
transform 1 0 34500 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_191_372
timestamp 1623621585
transform 1 0 35328 0 1 106080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_355
timestamp 1623621585
transform 1 0 33764 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_192_367
timestamp 1623621585
transform 1 0 34868 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input313
timestamp 1623621585
transform 1 0 37260 0 1 106080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input314
timestamp 1623621585
transform 1 0 37076 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_191_384
timestamp 1623621585
transform 1 0 36432 0 1 106080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_191_392
timestamp 1623621585
transform 1 0 37168 0 1 106080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_192_379
timestamp 1623621585
transform 1 0 35972 0 -1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_192_395
timestamp 1623621585
transform 1 0 37444 0 -1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_383
timestamp 1623621585
transform -1 0 38824 0 1 106080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_385
timestamp 1623621585
transform -1 0 38824 0 -1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1781
timestamp 1623621585
transform 1 0 37812 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_191_403
timestamp 1623621585
transform 1 0 38180 0 1 106080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_192_400
timestamp 1623621585
transform 1 0 37904 0 -1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_192_406
timestamp 1623621585
transform 1 0 38456 0 -1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_386
timestamp 1623621585
transform 1 0 1104 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_193_3
timestamp 1623621585
transform 1 0 1380 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_15
timestamp 1623621585
transform 1 0 2484 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1782
timestamp 1623621585
transform 1 0 3772 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_193_27
timestamp 1623621585
transform 1 0 3588 0 1 107168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_193_30
timestamp 1623621585
transform 1 0 3864 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_42
timestamp 1623621585
transform 1 0 4968 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_54
timestamp 1623621585
transform 1 0 6072 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_66
timestamp 1623621585
transform 1 0 7176 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_78
timestamp 1623621585
transform 1 0 8280 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1783
timestamp 1623621585
transform 1 0 9016 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_87
timestamp 1623621585
transform 1 0 9108 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_99
timestamp 1623621585
transform 1 0 10212 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_111
timestamp 1623621585
transform 1 0 11316 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_123
timestamp 1623621585
transform 1 0 12420 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1784
timestamp 1623621585
transform 1 0 14260 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_135
timestamp 1623621585
transform 1 0 13524 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_193_144
timestamp 1623621585
transform 1 0 14352 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_156
timestamp 1623621585
transform 1 0 15456 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_168
timestamp 1623621585
transform 1 0 16560 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_180
timestamp 1623621585
transform 1 0 17664 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1785
timestamp 1623621585
transform 1 0 19504 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_192
timestamp 1623621585
transform 1 0 18768 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_193_201
timestamp 1623621585
transform 1 0 19596 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_213
timestamp 1623621585
transform 1 0 20700 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_225
timestamp 1623621585
transform 1 0 21804 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_237
timestamp 1623621585
transform 1 0 22908 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_249
timestamp 1623621585
transform 1 0 24012 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1786
timestamp 1623621585
transform 1 0 24748 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_258
timestamp 1623621585
transform 1 0 24840 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_270
timestamp 1623621585
transform 1 0 25944 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_282
timestamp 1623621585
transform 1 0 27048 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_294
timestamp 1623621585
transform 1 0 28152 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_193_306
timestamp 1623621585
transform 1 0 29256 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1787
timestamp 1623621585
transform 1 0 29992 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_193_315
timestamp 1623621585
transform 1 0 30084 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_327
timestamp 1623621585
transform 1 0 31188 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_339
timestamp 1623621585
transform 1 0 32292 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_193_351
timestamp 1623621585
transform 1 0 33396 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1788
timestamp 1623621585
transform 1 0 35236 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_193_363
timestamp 1623621585
transform 1 0 34500 0 1 107168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_193_372
timestamp 1623621585
transform 1 0 35328 0 1 107168
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input316
timestamp 1623621585
transform 1 0 37076 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_193_384
timestamp 1623621585
transform 1 0 36432 0 1 107168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_193_390
timestamp 1623621585
transform 1 0 36984 0 1 107168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_193_395
timestamp 1623621585
transform 1 0 37444 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_387
timestamp 1623621585
transform -1 0 38824 0 1 107168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input315
timestamp 1623621585
transform 1 0 37812 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_193_403
timestamp 1623621585
transform 1 0 38180 0 1 107168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_388
timestamp 1623621585
transform 1 0 1104 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output663
timestamp 1623621585
transform 1 0 1748 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_194_3
timestamp 1623621585
transform 1 0 1380 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_194_11
timestamp 1623621585
transform 1 0 2116 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_23
timestamp 1623621585
transform 1 0 3220 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_35
timestamp 1623621585
transform 1 0 4324 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1789
timestamp 1623621585
transform 1 0 6348 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_47
timestamp 1623621585
transform 1 0 5428 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_194_55
timestamp 1623621585
transform 1 0 6164 0 -1 108256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_194_58
timestamp 1623621585
transform 1 0 6440 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_70
timestamp 1623621585
transform 1 0 7544 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_82
timestamp 1623621585
transform 1 0 8648 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_94
timestamp 1623621585
transform 1 0 9752 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1790
timestamp 1623621585
transform 1 0 11592 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_106
timestamp 1623621585
transform 1 0 10856 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_115
timestamp 1623621585
transform 1 0 11684 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_127
timestamp 1623621585
transform 1 0 12788 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_139
timestamp 1623621585
transform 1 0 13892 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_151
timestamp 1623621585
transform 1 0 14996 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_194_163
timestamp 1623621585
transform 1 0 16100 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1791
timestamp 1623621585
transform 1 0 16836 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_194_172
timestamp 1623621585
transform 1 0 16928 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_184
timestamp 1623621585
transform 1 0 18032 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_196
timestamp 1623621585
transform 1 0 19136 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_208
timestamp 1623621585
transform 1 0 20240 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1792
timestamp 1623621585
transform 1 0 22080 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_220
timestamp 1623621585
transform 1 0 21344 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_229
timestamp 1623621585
transform 1 0 22172 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_241
timestamp 1623621585
transform 1 0 23276 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_253
timestamp 1623621585
transform 1 0 24380 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_265
timestamp 1623621585
transform 1 0 25484 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1793
timestamp 1623621585
transform 1 0 27324 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_277
timestamp 1623621585
transform 1 0 26588 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_286
timestamp 1623621585
transform 1 0 27416 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_298
timestamp 1623621585
transform 1 0 28520 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_310
timestamp 1623621585
transform 1 0 29624 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_322
timestamp 1623621585
transform 1 0 30728 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1794
timestamp 1623621585
transform 1 0 32568 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_194_334
timestamp 1623621585
transform 1 0 31832 0 -1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_194_343
timestamp 1623621585
transform 1 0 32660 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_355
timestamp 1623621585
transform 1 0 33764 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_194_367
timestamp 1623621585
transform 1 0 34868 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input317
timestamp 1623621585
transform 1 0 37076 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_194_379
timestamp 1623621585
transform 1 0 35972 0 -1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_194_395
timestamp 1623621585
transform 1 0 37444 0 -1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_389
timestamp 1623621585
transform -1 0 38824 0 -1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1795
timestamp 1623621585
transform 1 0 37812 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_194_400
timestamp 1623621585
transform 1 0 37904 0 -1 108256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_194_406
timestamp 1623621585
transform 1 0 38456 0 -1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_390
timestamp 1623621585
transform 1 0 1104 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output664
timestamp 1623621585
transform 1 0 1748 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_195_3
timestamp 1623621585
transform 1 0 1380 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_195_11
timestamp 1623621585
transform 1 0 2116 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1796
timestamp 1623621585
transform 1 0 3772 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_195_23
timestamp 1623621585
transform 1 0 3220 0 1 108256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_195_30
timestamp 1623621585
transform 1 0 3864 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_42
timestamp 1623621585
transform 1 0 4968 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_54
timestamp 1623621585
transform 1 0 6072 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_66
timestamp 1623621585
transform 1 0 7176 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_78
timestamp 1623621585
transform 1 0 8280 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1797
timestamp 1623621585
transform 1 0 9016 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_87
timestamp 1623621585
transform 1 0 9108 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_99
timestamp 1623621585
transform 1 0 10212 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_111
timestamp 1623621585
transform 1 0 11316 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_123
timestamp 1623621585
transform 1 0 12420 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1798
timestamp 1623621585
transform 1 0 14260 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_195_135
timestamp 1623621585
transform 1 0 13524 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_144
timestamp 1623621585
transform 1 0 14352 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_156
timestamp 1623621585
transform 1 0 15456 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_168
timestamp 1623621585
transform 1 0 16560 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_180
timestamp 1623621585
transform 1 0 17664 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1799
timestamp 1623621585
transform 1 0 19504 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_195_192
timestamp 1623621585
transform 1 0 18768 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_201
timestamp 1623621585
transform 1 0 19596 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_213
timestamp 1623621585
transform 1 0 20700 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_225
timestamp 1623621585
transform 1 0 21804 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_237
timestamp 1623621585
transform 1 0 22908 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_249
timestamp 1623621585
transform 1 0 24012 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1800
timestamp 1623621585
transform 1 0 24748 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_258
timestamp 1623621585
transform 1 0 24840 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_270
timestamp 1623621585
transform 1 0 25944 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_282
timestamp 1623621585
transform 1 0 27048 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_294
timestamp 1623621585
transform 1 0 28152 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_195_306
timestamp 1623621585
transform 1 0 29256 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1801
timestamp 1623621585
transform 1 0 29992 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_195_315
timestamp 1623621585
transform 1 0 30084 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_327
timestamp 1623621585
transform 1 0 31188 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_339
timestamp 1623621585
transform 1 0 32292 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_351
timestamp 1623621585
transform 1 0 33396 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1802
timestamp 1623621585
transform 1 0 35236 0 1 108256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_195_363
timestamp 1623621585
transform 1 0 34500 0 1 108256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_195_372
timestamp 1623621585
transform 1 0 35328 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_195_384
timestamp 1623621585
transform 1 0 36432 0 1 108256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_391
timestamp 1623621585
transform -1 0 38824 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input318
timestamp 1623621585
transform 1 0 37812 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_195_396
timestamp 1623621585
transform 1 0 37536 0 1 108256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_195_403
timestamp 1623621585
transform 1 0 38180 0 1 108256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_392
timestamp 1623621585
transform 1 0 1104 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_196_3
timestamp 1623621585
transform 1 0 1380 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_15
timestamp 1623621585
transform 1 0 2484 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_27
timestamp 1623621585
transform 1 0 3588 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_39
timestamp 1623621585
transform 1 0 4692 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1803
timestamp 1623621585
transform 1 0 6348 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_196_51
timestamp 1623621585
transform 1 0 5796 0 -1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_196_58
timestamp 1623621585
transform 1 0 6440 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0943_
timestamp 1623621585
transform 1 0 8464 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_196_70
timestamp 1623621585
transform 1 0 7544 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_196_78
timestamp 1623621585
transform 1 0 8280 0 -1 109344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_196_83
timestamp 1623621585
transform 1 0 8740 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_95
timestamp 1623621585
transform 1 0 9844 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1804
timestamp 1623621585
transform 1 0 11592 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_196_107
timestamp 1623621585
transform 1 0 10948 0 -1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_113
timestamp 1623621585
transform 1 0 11500 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_115
timestamp 1623621585
transform 1 0 11684 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_127
timestamp 1623621585
transform 1 0 12788 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_139
timestamp 1623621585
transform 1 0 13892 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_151
timestamp 1623621585
transform 1 0 14996 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_196_163
timestamp 1623621585
transform 1 0 16100 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1805
timestamp 1623621585
transform 1 0 16836 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_196_172
timestamp 1623621585
transform 1 0 16928 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_184
timestamp 1623621585
transform 1 0 18032 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_196
timestamp 1623621585
transform 1 0 19136 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_208
timestamp 1623621585
transform 1 0 20240 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1806
timestamp 1623621585
transform 1 0 22080 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_220
timestamp 1623621585
transform 1 0 21344 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_229
timestamp 1623621585
transform 1 0 22172 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_241
timestamp 1623621585
transform 1 0 23276 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_253
timestamp 1623621585
transform 1 0 24380 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_265
timestamp 1623621585
transform 1 0 25484 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1807
timestamp 1623621585
transform 1 0 27324 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_277
timestamp 1623621585
transform 1 0 26588 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_286
timestamp 1623621585
transform 1 0 27416 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_298
timestamp 1623621585
transform 1 0 28520 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_310
timestamp 1623621585
transform 1 0 29624 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_322
timestamp 1623621585
transform 1 0 30728 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1808
timestamp 1623621585
transform 1 0 32568 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_196_334
timestamp 1623621585
transform 1 0 31832 0 -1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_196_343
timestamp 1623621585
transform 1 0 32660 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_355
timestamp 1623621585
transform 1 0 33764 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_196_367
timestamp 1623621585
transform 1 0 34868 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input319
timestamp 1623621585
transform 1 0 37076 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_196_379
timestamp 1623621585
transform 1 0 35972 0 -1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_196_395
timestamp 1623621585
transform 1 0 37444 0 -1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_393
timestamp 1623621585
transform -1 0 38824 0 -1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1809
timestamp 1623621585
transform 1 0 37812 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_196_400
timestamp 1623621585
transform 1 0 37904 0 -1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_196_406
timestamp 1623621585
transform 1 0 38456 0 -1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_394
timestamp 1623621585
transform 1 0 1104 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output667
timestamp 1623621585
transform 1 0 1748 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_197_3
timestamp 1623621585
transform 1 0 1380 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_197_11
timestamp 1623621585
transform 1 0 2116 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1810
timestamp 1623621585
transform 1 0 3772 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_197_23
timestamp 1623621585
transform 1 0 3220 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_197_30
timestamp 1623621585
transform 1 0 3864 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_42
timestamp 1623621585
transform 1 0 4968 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_54
timestamp 1623621585
transform 1 0 6072 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_66
timestamp 1623621585
transform 1 0 7176 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_78
timestamp 1623621585
transform 1 0 8280 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1811
timestamp 1623621585
transform 1 0 9016 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_87
timestamp 1623621585
transform 1 0 9108 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_99
timestamp 1623621585
transform 1 0 10212 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_111
timestamp 1623621585
transform 1 0 11316 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_123
timestamp 1623621585
transform 1 0 12420 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1812
timestamp 1623621585
transform 1 0 14260 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_197_135
timestamp 1623621585
transform 1 0 13524 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_144
timestamp 1623621585
transform 1 0 14352 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_156
timestamp 1623621585
transform 1 0 15456 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_168
timestamp 1623621585
transform 1 0 16560 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_180
timestamp 1623621585
transform 1 0 17664 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1813
timestamp 1623621585
transform 1 0 19504 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_197_192
timestamp 1623621585
transform 1 0 18768 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_201
timestamp 1623621585
transform 1 0 19596 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_213
timestamp 1623621585
transform 1 0 20700 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_225
timestamp 1623621585
transform 1 0 21804 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_237
timestamp 1623621585
transform 1 0 22908 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_249
timestamp 1623621585
transform 1 0 24012 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1814
timestamp 1623621585
transform 1 0 24748 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_258
timestamp 1623621585
transform 1 0 24840 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_270
timestamp 1623621585
transform 1 0 25944 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_282
timestamp 1623621585
transform 1 0 27048 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_294
timestamp 1623621585
transform 1 0 28152 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_197_306
timestamp 1623621585
transform 1 0 29256 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1815
timestamp 1623621585
transform 1 0 29992 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_197_315
timestamp 1623621585
transform 1 0 30084 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_327
timestamp 1623621585
transform 1 0 31188 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_339
timestamp 1623621585
transform 1 0 32292 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_197_351
timestamp 1623621585
transform 1 0 33396 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1816
timestamp 1623621585
transform 1 0 35236 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_197_363
timestamp 1623621585
transform 1 0 34500 0 1 109344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_197_372
timestamp 1623621585
transform 1 0 35328 0 1 109344
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input322
timestamp 1623621585
transform 1 0 37076 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_197_384
timestamp 1623621585
transform 1 0 36432 0 1 109344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_197_390
timestamp 1623621585
transform 1 0 36984 0 1 109344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_197_395
timestamp 1623621585
transform 1 0 37444 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_395
timestamp 1623621585
transform -1 0 38824 0 1 109344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input320
timestamp 1623621585
transform 1 0 37812 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_197_403
timestamp 1623621585
transform 1 0 38180 0 1 109344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_396
timestamp 1623621585
transform 1 0 1104 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_398
timestamp 1623621585
transform 1 0 1104 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output701
timestamp 1623621585
transform 1 0 1748 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_198_3
timestamp 1623621585
transform 1 0 1380 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_15
timestamp 1623621585
transform 1 0 2484 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_199_3
timestamp 1623621585
transform 1 0 1380 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_199_11
timestamp 1623621585
transform 1 0 2116 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1824
timestamp 1623621585
transform 1 0 3772 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_27
timestamp 1623621585
transform 1 0 3588 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_39
timestamp 1623621585
transform 1 0 4692 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_199_23
timestamp 1623621585
transform 1 0 3220 0 1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_199_30
timestamp 1623621585
transform 1 0 3864 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1817
timestamp 1623621585
transform 1 0 6348 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_198_51
timestamp 1623621585
transform 1 0 5796 0 -1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_198_58
timestamp 1623621585
transform 1 0 6440 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_42
timestamp 1623621585
transform 1 0 4968 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_54
timestamp 1623621585
transform 1 0 6072 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_70
timestamp 1623621585
transform 1 0 7544 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_82
timestamp 1623621585
transform 1 0 8648 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_66
timestamp 1623621585
transform 1 0 7176 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_78
timestamp 1623621585
transform 1 0 8280 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1825
timestamp 1623621585
transform 1 0 9016 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_94
timestamp 1623621585
transform 1 0 9752 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_87
timestamp 1623621585
transform 1 0 9108 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_99
timestamp 1623621585
transform 1 0 10212 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1818
timestamp 1623621585
transform 1 0 11592 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_106
timestamp 1623621585
transform 1 0 10856 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_115
timestamp 1623621585
transform 1 0 11684 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_111
timestamp 1623621585
transform 1 0 11316 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_123
timestamp 1623621585
transform 1 0 12420 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1826
timestamp 1623621585
transform 1 0 14260 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_127
timestamp 1623621585
transform 1 0 12788 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_139
timestamp 1623621585
transform 1 0 13892 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_135
timestamp 1623621585
transform 1 0 13524 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_144
timestamp 1623621585
transform 1 0 14352 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_151
timestamp 1623621585
transform 1 0 14996 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_198_163
timestamp 1623621585
transform 1 0 16100 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_156
timestamp 1623621585
transform 1 0 15456 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1819
timestamp 1623621585
transform 1 0 16836 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_172
timestamp 1623621585
transform 1 0 16928 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_184
timestamp 1623621585
transform 1 0 18032 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_168
timestamp 1623621585
transform 1 0 16560 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_180
timestamp 1623621585
transform 1 0 17664 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1827
timestamp 1623621585
transform 1 0 19504 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_196
timestamp 1623621585
transform 1 0 19136 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_208
timestamp 1623621585
transform 1 0 20240 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_192
timestamp 1623621585
transform 1 0 18768 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_201
timestamp 1623621585
transform 1 0 19596 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1820
timestamp 1623621585
transform 1 0 22080 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_220
timestamp 1623621585
transform 1 0 21344 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_229
timestamp 1623621585
transform 1 0 22172 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_213
timestamp 1623621585
transform 1 0 20700 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_225
timestamp 1623621585
transform 1 0 21804 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_241
timestamp 1623621585
transform 1 0 23276 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_237
timestamp 1623621585
transform 1 0 22908 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_249
timestamp 1623621585
transform 1 0 24012 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1828
timestamp 1623621585
transform 1 0 24748 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_253
timestamp 1623621585
transform 1 0 24380 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_265
timestamp 1623621585
transform 1 0 25484 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_258
timestamp 1623621585
transform 1 0 24840 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_270
timestamp 1623621585
transform 1 0 25944 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1821
timestamp 1623621585
transform 1 0 27324 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_277
timestamp 1623621585
transform 1 0 26588 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_286
timestamp 1623621585
transform 1 0 27416 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_282
timestamp 1623621585
transform 1 0 27048 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_298
timestamp 1623621585
transform 1 0 28520 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_310
timestamp 1623621585
transform 1 0 29624 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_294
timestamp 1623621585
transform 1 0 28152 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_306
timestamp 1623621585
transform 1 0 29256 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1829
timestamp 1623621585
transform 1 0 29992 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_322
timestamp 1623621585
transform 1 0 30728 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_315
timestamp 1623621585
transform 1 0 30084 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_327
timestamp 1623621585
transform 1 0 31188 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1822
timestamp 1623621585
transform 1 0 32568 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_198_334
timestamp 1623621585
transform 1 0 31832 0 -1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_198_343
timestamp 1623621585
transform 1 0 32660 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_339
timestamp 1623621585
transform 1 0 32292 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_199_351
timestamp 1623621585
transform 1 0 33396 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1830
timestamp 1623621585
transform 1 0 35236 0 1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_198_355
timestamp 1623621585
transform 1 0 33764 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_198_367
timestamp 1623621585
transform 1 0 34868 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_199_363
timestamp 1623621585
transform 1 0 34500 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_199_372
timestamp 1623621585
transform 1 0 35328 0 1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  input63
timestamp 1623621585
transform 1 0 37352 0 1 110432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input323
timestamp 1623621585
transform 1 0 37076 0 -1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_198_379
timestamp 1623621585
transform 1 0 35972 0 -1 110432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_198_395
timestamp 1623621585
transform 1 0 37444 0 -1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_199_384
timestamp 1623621585
transform 1 0 36432 0 1 110432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_199_392
timestamp 1623621585
transform 1 0 37168 0 1 110432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_397
timestamp 1623621585
transform -1 0 38824 0 -1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_399
timestamp 1623621585
transform -1 0 38824 0 1 110432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1823
timestamp 1623621585
transform 1 0 37812 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_198_400
timestamp 1623621585
transform 1 0 37904 0 -1 110432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_198_406
timestamp 1623621585
transform 1 0 38456 0 -1 110432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_199_403
timestamp 1623621585
transform 1 0 38180 0 1 110432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_400
timestamp 1623621585
transform 1 0 1104 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input73
timestamp 1623621585
transform 1 0 1380 0 -1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_200_9
timestamp 1623621585
transform 1 0 1932 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_21
timestamp 1623621585
transform 1 0 3036 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_33
timestamp 1623621585
transform 1 0 4140 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1831
timestamp 1623621585
transform 1 0 6348 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_45
timestamp 1623621585
transform 1 0 5244 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_58
timestamp 1623621585
transform 1 0 6440 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_70
timestamp 1623621585
transform 1 0 7544 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_82
timestamp 1623621585
transform 1 0 8648 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_94
timestamp 1623621585
transform 1 0 9752 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1832
timestamp 1623621585
transform 1 0 11592 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_106
timestamp 1623621585
transform 1 0 10856 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_115
timestamp 1623621585
transform 1 0 11684 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_127
timestamp 1623621585
transform 1 0 12788 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_139
timestamp 1623621585
transform 1 0 13892 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_151
timestamp 1623621585
transform 1 0 14996 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_200_163
timestamp 1623621585
transform 1 0 16100 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1833
timestamp 1623621585
transform 1 0 16836 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_200_172
timestamp 1623621585
transform 1 0 16928 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_184
timestamp 1623621585
transform 1 0 18032 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_196
timestamp 1623621585
transform 1 0 19136 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_208
timestamp 1623621585
transform 1 0 20240 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1834
timestamp 1623621585
transform 1 0 22080 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_220
timestamp 1623621585
transform 1 0 21344 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_229
timestamp 1623621585
transform 1 0 22172 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_241
timestamp 1623621585
transform 1 0 23276 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_253
timestamp 1623621585
transform 1 0 24380 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_265
timestamp 1623621585
transform 1 0 25484 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1835
timestamp 1623621585
transform 1 0 27324 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_277
timestamp 1623621585
transform 1 0 26588 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_286
timestamp 1623621585
transform 1 0 27416 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_298
timestamp 1623621585
transform 1 0 28520 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_310
timestamp 1623621585
transform 1 0 29624 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0950_
timestamp 1623621585
transform 1 0 31556 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_200_322
timestamp 1623621585
transform 1 0 30728 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_200_330
timestamp 1623621585
transform 1 0 31464 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1836
timestamp 1623621585
transform 1 0 32568 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_200_334
timestamp 1623621585
transform 1 0 31832 0 -1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_200_343
timestamp 1623621585
transform 1 0 32660 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_355
timestamp 1623621585
transform 1 0 33764 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_200_367
timestamp 1623621585
transform 1 0 34868 0 -1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output648
timestamp 1623621585
transform 1 0 37076 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output672
timestamp 1623621585
transform 1 0 36340 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_200_379
timestamp 1623621585
transform 1 0 35972 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_200_387
timestamp 1623621585
transform 1 0 36708 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_200_395
timestamp 1623621585
transform 1 0 37444 0 -1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_401
timestamp 1623621585
transform -1 0 38824 0 -1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1837
timestamp 1623621585
transform 1 0 37812 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_200_400
timestamp 1623621585
transform 1 0 37904 0 -1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_200_406
timestamp 1623621585
transform 1 0 38456 0 -1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_402
timestamp 1623621585
transform 1 0 1104 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_201_3
timestamp 1623621585
transform 1 0 1380 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_15
timestamp 1623621585
transform 1 0 2484 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1838
timestamp 1623621585
transform 1 0 3772 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_201_27
timestamp 1623621585
transform 1 0 3588 0 1 111520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_201_30
timestamp 1623621585
transform 1 0 3864 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_42
timestamp 1623621585
transform 1 0 4968 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_54
timestamp 1623621585
transform 1 0 6072 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_66
timestamp 1623621585
transform 1 0 7176 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_78
timestamp 1623621585
transform 1 0 8280 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1839
timestamp 1623621585
transform 1 0 9016 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_87
timestamp 1623621585
transform 1 0 9108 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_99
timestamp 1623621585
transform 1 0 10212 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_111
timestamp 1623621585
transform 1 0 11316 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_123
timestamp 1623621585
transform 1 0 12420 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1840
timestamp 1623621585
transform 1 0 14260 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_135
timestamp 1623621585
transform 1 0 13524 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_144
timestamp 1623621585
transform 1 0 14352 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_156
timestamp 1623621585
transform 1 0 15456 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_168
timestamp 1623621585
transform 1 0 16560 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_180
timestamp 1623621585
transform 1 0 17664 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1841
timestamp 1623621585
transform 1 0 19504 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_192
timestamp 1623621585
transform 1 0 18768 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_201
timestamp 1623621585
transform 1 0 19596 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_213
timestamp 1623621585
transform 1 0 20700 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_225
timestamp 1623621585
transform 1 0 21804 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_237
timestamp 1623621585
transform 1 0 22908 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_249
timestamp 1623621585
transform 1 0 24012 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1842
timestamp 1623621585
transform 1 0 24748 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_258
timestamp 1623621585
transform 1 0 24840 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_270
timestamp 1623621585
transform 1 0 25944 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_282
timestamp 1623621585
transform 1 0 27048 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_294
timestamp 1623621585
transform 1 0 28152 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_201_306
timestamp 1623621585
transform 1 0 29256 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1843
timestamp 1623621585
transform 1 0 29992 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_201_315
timestamp 1623621585
transform 1 0 30084 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_327
timestamp 1623621585
transform 1 0 31188 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_339
timestamp 1623621585
transform 1 0 32292 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_351
timestamp 1623621585
transform 1 0 33396 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1844
timestamp 1623621585
transform 1 0 35236 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_201_363
timestamp 1623621585
transform 1 0 34500 0 1 111520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_201_372
timestamp 1623621585
transform 1 0 35328 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_201_384
timestamp 1623621585
transform 1 0 36432 0 1 111520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_403
timestamp 1623621585
transform -1 0 38824 0 1 111520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1623621585
transform 1 0 37628 0 1 111520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_201_396
timestamp 1623621585
transform 1 0 37536 0 1 111520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_201_403
timestamp 1623621585
transform 1 0 38180 0 1 111520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_404
timestamp 1623621585
transform 1 0 1104 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output670
timestamp 1623621585
transform 1 0 1748 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_3
timestamp 1623621585
transform 1 0 1380 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_202_11
timestamp 1623621585
transform 1 0 2116 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_23
timestamp 1623621585
transform 1 0 3220 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_35
timestamp 1623621585
transform 1 0 4324 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1845
timestamp 1623621585
transform 1 0 6348 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_47
timestamp 1623621585
transform 1 0 5428 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_202_55
timestamp 1623621585
transform 1 0 6164 0 -1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_202_58
timestamp 1623621585
transform 1 0 6440 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_70
timestamp 1623621585
transform 1 0 7544 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_82
timestamp 1623621585
transform 1 0 8648 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_94
timestamp 1623621585
transform 1 0 9752 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1846
timestamp 1623621585
transform 1 0 11592 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_106
timestamp 1623621585
transform 1 0 10856 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_115
timestamp 1623621585
transform 1 0 11684 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_127
timestamp 1623621585
transform 1 0 12788 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_139
timestamp 1623621585
transform 1 0 13892 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_151
timestamp 1623621585
transform 1 0 14996 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_202_163
timestamp 1623621585
transform 1 0 16100 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1847
timestamp 1623621585
transform 1 0 16836 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_202_172
timestamp 1623621585
transform 1 0 16928 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_184
timestamp 1623621585
transform 1 0 18032 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_196
timestamp 1623621585
transform 1 0 19136 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_208
timestamp 1623621585
transform 1 0 20240 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1848
timestamp 1623621585
transform 1 0 22080 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_220
timestamp 1623621585
transform 1 0 21344 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_229
timestamp 1623621585
transform 1 0 22172 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_241
timestamp 1623621585
transform 1 0 23276 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_253
timestamp 1623621585
transform 1 0 24380 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_265
timestamp 1623621585
transform 1 0 25484 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1849
timestamp 1623621585
transform 1 0 27324 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_277
timestamp 1623621585
transform 1 0 26588 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_286
timestamp 1623621585
transform 1 0 27416 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_298
timestamp 1623621585
transform 1 0 28520 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_310
timestamp 1623621585
transform 1 0 29624 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_322
timestamp 1623621585
transform 1 0 30728 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1850
timestamp 1623621585
transform 1 0 32568 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_202_334
timestamp 1623621585
transform 1 0 31832 0 -1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_202_343
timestamp 1623621585
transform 1 0 32660 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_355
timestamp 1623621585
transform 1 0 33764 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_202_367
timestamp 1623621585
transform 1 0 34868 0 -1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output693
timestamp 1623621585
transform 1 0 37076 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output697
timestamp 1623621585
transform 1 0 36340 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_379
timestamp 1623621585
transform 1 0 35972 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_387
timestamp 1623621585
transform 1 0 36708 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_202_395
timestamp 1623621585
transform 1 0 37444 0 -1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_405
timestamp 1623621585
transform -1 0 38824 0 -1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1851
timestamp 1623621585
transform 1 0 37812 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_202_400
timestamp 1623621585
transform 1 0 37904 0 -1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_202_406
timestamp 1623621585
transform 1 0 38456 0 -1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_406
timestamp 1623621585
transform 1 0 1104 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1623621585
transform 1 0 2668 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input74
timestamp 1623621585
transform 1 0 1748 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_203_3
timestamp 1623621585
transform 1 0 1380 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_13
timestamp 1623621585
transform 1 0 2300 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_203_20
timestamp 1623621585
transform 1 0 2944 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1852
timestamp 1623621585
transform 1 0 3772 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1623621585
transform 1 0 4232 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1623621585
transform 1 0 4876 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_203_28
timestamp 1623621585
transform 1 0 3680 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_203_30
timestamp 1623621585
transform 1 0 3864 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_37
timestamp 1623621585
transform 1 0 4508 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1623621585
transform 1 0 5520 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1623621585
transform 1 0 6164 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1623621585
transform 1 0 6808 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_203_44
timestamp 1623621585
transform 1 0 5152 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_51
timestamp 1623621585
transform 1 0 5796 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_58
timestamp 1623621585
transform 1 0 6440 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1623621585
transform 1 0 7452 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_203_65
timestamp 1623621585
transform 1 0 7084 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_203_72
timestamp 1623621585
transform 1 0 7728 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1853
timestamp 1623621585
transform 1 0 9016 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_203_84
timestamp 1623621585
transform 1 0 8832 0 1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_203_87
timestamp 1623621585
transform 1 0 9108 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_99
timestamp 1623621585
transform 1 0 10212 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_111
timestamp 1623621585
transform 1 0 11316 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_123
timestamp 1623621585
transform 1 0 12420 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1854
timestamp 1623621585
transform 1 0 14260 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_203_135
timestamp 1623621585
transform 1 0 13524 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_203_144
timestamp 1623621585
transform 1 0 14352 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_156
timestamp 1623621585
transform 1 0 15456 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_168
timestamp 1623621585
transform 1 0 16560 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_180
timestamp 1623621585
transform 1 0 17664 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1855
timestamp 1623621585
transform 1 0 19504 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_203_192
timestamp 1623621585
transform 1 0 18768 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_203_201
timestamp 1623621585
transform 1 0 19596 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_213
timestamp 1623621585
transform 1 0 20700 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_225
timestamp 1623621585
transform 1 0 21804 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_237
timestamp 1623621585
transform 1 0 22908 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_203_249
timestamp 1623621585
transform 1 0 24012 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1856
timestamp 1623621585
transform 1 0 24748 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_203_258
timestamp 1623621585
transform 1 0 24840 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_270
timestamp 1623621585
transform 1 0 25944 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_203_282
timestamp 1623621585
transform 1 0 27048 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0778_
timestamp 1623621585
transform 1 0 28152 0 1 112608
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_203_303
timestamp 1623621585
transform 1 0 28980 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_203_311
timestamp 1623621585
transform 1 0 29716 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1857
timestamp 1623621585
transform 1 0 29992 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input474
timestamp 1623621585
transform 1 0 31372 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_203_315
timestamp 1623621585
transform 1 0 30084 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_203_327
timestamp 1623621585
transform 1 0 31188 0 1 112608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_203_332
timestamp 1623621585
transform 1 0 31648 0 1 112608
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1623621585
transform 1 0 33304 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_203_344
timestamp 1623621585
transform 1 0 32752 0 1 112608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_203_353
timestamp 1623621585
transform 1 0 33580 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1858
timestamp 1623621585
transform 1 0 35236 0 1 112608
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1623621585
transform 1 0 33948 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_203_360
timestamp 1623621585
transform 1 0 34224 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_203_368
timestamp 1623621585
transform 1 0 34960 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_203_372
timestamp 1623621585
transform 1 0 35328 0 1 112608
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output653
timestamp 1623621585
transform 1 0 37076 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output691
timestamp 1623621585
transform 1 0 36340 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_203_380
timestamp 1623621585
transform 1 0 36064 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_203_387
timestamp 1623621585
transform 1 0 36708 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_395
timestamp 1623621585
transform 1 0 37444 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_407
timestamp 1623621585
transform -1 0 38824 0 1 112608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output651
timestamp 1623621585
transform 1 0 37812 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_203_403
timestamp 1623621585
transform 1 0 38180 0 1 112608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_3
timestamp 1623621585
transform 1 0 1380 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_7
timestamp 1623621585
transform 1 0 1748 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_3
timestamp 1623621585
transform 1 0 1380 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output659
timestamp 1623621585
transform 1 0 1748 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1623621585
transform 1 0 1472 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_410
timestamp 1623621585
transform 1 0 1104 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_408
timestamp 1623621585
transform 1 0 1104 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_205_11
timestamp 1623621585
transform 1 0 2116 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_204_14
timestamp 1623621585
transform 1 0 2392 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0869_
timestamp 1623621585
transform 1 0 2116 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0870_
timestamp 1623621585
transform 1 0 2760 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0849_
timestamp 1623621585
transform 1 0 2852 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_28
timestamp 1623621585
transform 1 0 3680 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_205_22
timestamp 1623621585
transform 1 0 3128 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_204_28
timestamp 1623621585
transform 1 0 3680 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_204_21
timestamp 1623621585
transform 1 0 3036 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1623621585
transform 1 0 3404 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1866
timestamp 1623621585
transform 1 0 3772 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_37
timestamp 1623621585
transform 1 0 4508 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_30
timestamp 1623621585
transform 1 0 3864 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_204_36
timestamp 1623621585
transform 1 0 4416 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1623621585
transform 1 0 4600 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0871_
timestamp 1623621585
transform 1 0 4232 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_204_41
timestamp 1623621585
transform 1 0 4876 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0872_
timestamp 1623621585
transform 1 0 4876 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_48
timestamp 1623621585
transform 1 0 5520 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_44
timestamp 1623621585
transform 1 0 5152 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_204_48
timestamp 1623621585
transform 1 0 5520 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0900_
timestamp 1623621585
transform 1 0 5244 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0874_
timestamp 1623621585
transform 1 0 5612 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_205_52
timestamp 1623621585
transform 1 0 5888 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_204_58
timestamp 1623621585
transform 1 0 6440 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_204_56
timestamp 1623621585
transform 1 0 6256 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1859
timestamp 1623621585
transform 1 0 6348 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_205_60
timestamp 1623621585
transform 1 0 6624 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _0902_
timestamp 1623621585
transform 1 0 6808 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0876_
timestamp 1623621585
transform 1 0 6808 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_65
timestamp 1623621585
transform 1 0 7084 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_65
timestamp 1623621585
transform 1 0 7084 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1623621585
transform 1 0 7452 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1623621585
transform 1 0 7452 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_72
timestamp 1623621585
transform 1 0 7728 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_72
timestamp 1623621585
transform 1 0 7728 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0906_
timestamp 1623621585
transform 1 0 8096 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 1623621585
transform 1 0 8096 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_205_79
timestamp 1623621585
transform 1 0 8372 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_204_79
timestamp 1623621585
transform 1 0 8372 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1623621585
transform 1 0 8740 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1867
timestamp 1623621585
transform 1 0 9016 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1623621585
transform 1 0 9476 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_86
timestamp 1623621585
transform 1 0 9016 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_98
timestamp 1623621585
transform 1 0 10120 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_205_85
timestamp 1623621585
transform 1 0 8924 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_87
timestamp 1623621585
transform 1 0 9108 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_205_94
timestamp 1623621585
transform 1 0 9752 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1860
timestamp 1623621585
transform 1 0 11592 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_204_110
timestamp 1623621585
transform 1 0 11224 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_204_115
timestamp 1623621585
transform 1 0 11684 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_106
timestamp 1623621585
transform 1 0 10856 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_118
timestamp 1623621585
transform 1 0 11960 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1868
timestamp 1623621585
transform 1 0 14260 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_204_127
timestamp 1623621585
transform 1 0 12788 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_139
timestamp 1623621585
transform 1 0 13892 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_130
timestamp 1623621585
transform 1 0 13064 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_205_142
timestamp 1623621585
transform 1 0 14168 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_205_144
timestamp 1623621585
transform 1 0 14352 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1623621585
transform 1 0 15732 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1623621585
transform 1 0 16376 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_151
timestamp 1623621585
transform 1 0 14996 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_204_163
timestamp 1623621585
transform 1 0 16100 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_205_156
timestamp 1623621585
transform 1 0 15456 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_162
timestamp 1623621585
transform 1 0 16008 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1861
timestamp 1623621585
transform 1 0 16836 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1623621585
transform 1 0 17664 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1623621585
transform 1 0 18308 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_172
timestamp 1623621585
transform 1 0 16928 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_184
timestamp 1623621585
transform 1 0 18032 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_169
timestamp 1623621585
transform 1 0 16652 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_205_177
timestamp 1623621585
transform 1 0 17388 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_183
timestamp 1623621585
transform 1 0 17940 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1869
timestamp 1623621585
transform 1 0 19504 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1623621585
transform 1 0 20148 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_196
timestamp 1623621585
transform 1 0 19136 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_208
timestamp 1623621585
transform 1 0 20240 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_205_190
timestamp 1623621585
transform 1 0 18584 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_205_198
timestamp 1623621585
transform 1 0 19320 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_205_201
timestamp 1623621585
transform 1 0 19596 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_205_217
timestamp 1623621585
transform 1 0 21068 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_210
timestamp 1623621585
transform 1 0 20424 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1623621585
transform 1 0 20792 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_205_225
timestamp 1623621585
transform 1 0 21804 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_221
timestamp 1623621585
transform 1 0 21436 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_204_220
timestamp 1623621585
transform 1 0 21344 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1623621585
transform 1 0 22172 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1862
timestamp 1623621585
transform 1 0 22080 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1623621585
transform 1 0 21528 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_229
timestamp 1623621585
transform 1 0 22172 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1623621585
transform 1 0 22816 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1623621585
transform 1 0 23460 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1623621585
transform 1 0 24104 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_241
timestamp 1623621585
transform 1 0 23276 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_205_232
timestamp 1623621585
transform 1 0 22448 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_239
timestamp 1623621585
transform 1 0 23092 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_246
timestamp 1623621585
transform 1 0 23736 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_258
timestamp 1623621585
transform 1 0 24840 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_253
timestamp 1623621585
transform 1 0 24380 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_258
timestamp 1623621585
transform 1 0 24840 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_204_253
timestamp 1623621585
transform 1 0 24380 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1623621585
transform 1 0 24564 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1870
timestamp 1623621585
transform 1 0 24748 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_205_265
timestamp 1623621585
transform 1 0 25484 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1623621585
transform 1 0 25208 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1623621585
transform 1 0 25208 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_265
timestamp 1623621585
transform 1 0 25484 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1623621585
transform 1 0 26220 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1863
timestamp 1623621585
transform 1 0 27324 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_204_277
timestamp 1623621585
transform 1 0 26588 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_204_286
timestamp 1623621585
transform 1 0 27416 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_276
timestamp 1623621585
transform 1 0 26496 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_205_288
timestamp 1623621585
transform 1 0 27600 0 1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input466
timestamp 1623621585
transform 1 0 29256 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_204_298
timestamp 1623621585
transform 1 0 28520 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_204_310
timestamp 1623621585
transform 1 0 29624 0 -1 113696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_205_300
timestamp 1623621585
transform 1 0 28704 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_205_309
timestamp 1623621585
transform 1 0 29532 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_315
timestamp 1623621585
transform 1 0 30084 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_205_313
timestamp 1623621585
transform 1 0 29900 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input468
timestamp 1623621585
transform 1 0 30452 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1871
timestamp 1623621585
transform 1 0 29992 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_329
timestamp 1623621585
transform 1 0 31372 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_322
timestamp 1623621585
transform 1 0 30728 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_325
timestamp 1623621585
transform 1 0 31004 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input473
timestamp 1623621585
transform 1 0 31372 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input471
timestamp 1623621585
transform 1 0 30728 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input470
timestamp 1623621585
transform 1 0 31096 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_204_332
timestamp 1623621585
transform 1 0 31648 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input472
timestamp 1623621585
transform 1 0 31740 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_205_340
timestamp 1623621585
transform 1 0 32384 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_336
timestamp 1623621585
transform 1 0 32016 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_204_340
timestamp 1623621585
transform 1 0 32384 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1623621585
transform 1 0 32476 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1864
timestamp 1623621585
transform 1 0 32568 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_205_344
timestamp 1623621585
transform 1 0 32752 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_204_350
timestamp 1623621585
transform 1 0 33304 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_343
timestamp 1623621585
transform 1 0 32660 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1623621585
transform 1 0 33028 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_205_352
timestamp 1623621585
transform 1 0 33488 0 1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1623621585
transform 1 0 33672 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1623621585
transform 1 0 33672 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_205_357
timestamp 1623621585
transform 1 0 33948 0 1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_204_357
timestamp 1623621585
transform 1 0 33948 0 -1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output702
timestamp 1623621585
transform 1 0 34500 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_367
timestamp 1623621585
transform 1 0 34868 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_371
timestamp 1623621585
transform 1 0 35236 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_204_365
timestamp 1623621585
transform 1 0 34684 0 -1 113696
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output703
timestamp 1623621585
transform 1 0 34868 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1872
timestamp 1623621585
transform 1 0 35236 0 1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_205_372
timestamp 1623621585
transform 1 0 35328 0 1 113696
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output692
timestamp 1623621585
transform 1 0 35604 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_379
timestamp 1623621585
transform 1 0 35972 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_205_380
timestamp 1623621585
transform 1 0 36064 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output687
timestamp 1623621585
transform 1 0 36340 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output680
timestamp 1623621585
transform 1 0 36340 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_387
timestamp 1623621585
transform 1 0 36708 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_387
timestamp 1623621585
transform 1 0 36708 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output666
timestamp 1623621585
transform 1 0 37076 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output665
timestamp 1623621585
transform 1 0 37076 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_205_395
timestamp 1623621585
transform 1 0 37444 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_204_395
timestamp 1623621585
transform 1 0 37444 0 -1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_409
timestamp 1623621585
transform -1 0 38824 0 -1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_411
timestamp 1623621585
transform -1 0 38824 0 1 113696
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1865
timestamp 1623621585
transform 1 0 37812 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output657
timestamp 1623621585
transform 1 0 37812 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_204_400
timestamp 1623621585
transform 1 0 37904 0 -1 113696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_204_406
timestamp 1623621585
transform 1 0 38456 0 -1 113696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_205_403
timestamp 1623621585
transform 1 0 38180 0 1 113696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_412
timestamp 1623621585
transform 1 0 1104 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output649
timestamp 1623621585
transform 1 0 1748 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output684
timestamp 1623621585
transform 1 0 2484 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_3
timestamp 1623621585
transform 1 0 1380 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_11
timestamp 1623621585
transform 1 0 2116 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_19
timestamp 1623621585
transform 1 0 2852 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0851_
timestamp 1623621585
transform 1 0 3956 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0853_
timestamp 1623621585
transform 1 0 4876 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output695
timestamp 1623621585
transform 1 0 3220 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_27
timestamp 1623621585
transform 1 0 3588 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_34
timestamp 1623621585
transform 1 0 4232 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_40
timestamp 1623621585
transform 1 0 4784 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _0857_
timestamp 1623621585
transform 1 0 6808 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0873_
timestamp 1623621585
transform 1 0 5520 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1873
timestamp 1623621585
transform 1 0 6348 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_44
timestamp 1623621585
transform 1 0 5152 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_51
timestamp 1623621585
transform 1 0 5796 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_206_58
timestamp 1623621585
transform 1 0 6440 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0875_
timestamp 1623621585
transform 1 0 7452 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0877_
timestamp 1623621585
transform 1 0 8372 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_65
timestamp 1623621585
transform 1 0 7084 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_72
timestamp 1623621585
transform 1 0 7728 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_78
timestamp 1623621585
transform 1 0 8280 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_82
timestamp 1623621585
transform 1 0 8648 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1623621585
transform 1 0 9016 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1623621585
transform 1 0 9660 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1623621585
transform 1 0 10304 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_89
timestamp 1623621585
transform 1 0 9292 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_96
timestamp 1623621585
transform 1 0 9936 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_103
timestamp 1623621585
transform 1 0 10580 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1874
timestamp 1623621585
transform 1 0 11592 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1623621585
transform 1 0 10948 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1623621585
transform 1 0 12052 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_110
timestamp 1623621585
transform 1 0 11224 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_115
timestamp 1623621585
transform 1 0 11684 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_122
timestamp 1623621585
transform 1 0 12328 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1623621585
transform 1 0 12696 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1623621585
transform 1 0 13340 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1623621585
transform 1 0 13984 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_129
timestamp 1623621585
transform 1 0 12972 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_136
timestamp 1623621585
transform 1 0 13616 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_143
timestamp 1623621585
transform 1 0 14260 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1623621585
transform 1 0 14628 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1623621585
transform 1 0 15272 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1623621585
transform 1 0 15916 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_150
timestamp 1623621585
transform 1 0 14904 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_157
timestamp 1623621585
transform 1 0 15548 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_164
timestamp 1623621585
transform 1 0 16192 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1623621585
transform 1 0 18032 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1875
timestamp 1623621585
transform 1 0 16836 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1623621585
transform 1 0 17296 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_206_170
timestamp 1623621585
transform 1 0 16744 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_172
timestamp 1623621585
transform 1 0 16928 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_179
timestamp 1623621585
transform 1 0 17572 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_206_183
timestamp 1623621585
transform 1 0 17940 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_187
timestamp 1623621585
transform 1 0 18308 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1623621585
transform 1 0 18676 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1623621585
transform 1 0 19320 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1623621585
transform 1 0 19964 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_194
timestamp 1623621585
transform 1 0 18952 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_201
timestamp 1623621585
transform 1 0 19596 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_208
timestamp 1623621585
transform 1 0 20240 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1623621585
transform 1 0 20792 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1623621585
transform 1 0 21436 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1876
timestamp 1623621585
transform 1 0 22080 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_217
timestamp 1623621585
transform 1 0 21068 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_224
timestamp 1623621585
transform 1 0 21712 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_229
timestamp 1623621585
transform 1 0 22172 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1623621585
transform 1 0 24012 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1623621585
transform 1 0 22540 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1623621585
transform 1 0 23184 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_236
timestamp 1623621585
transform 1 0 22816 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_206_243
timestamp 1623621585
transform 1 0 23460 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1623621585
transform 1 0 24932 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1623621585
transform 1 0 25576 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_206_252
timestamp 1623621585
transform 1 0 24288 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_258
timestamp 1623621585
transform 1 0 24840 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_262
timestamp 1623621585
transform 1 0 25208 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_269
timestamp 1623621585
transform 1 0 25852 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1623621585
transform 1 0 26220 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1877
timestamp 1623621585
transform 1 0 27324 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_206_276
timestamp 1623621585
transform 1 0 26496 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_206_284
timestamp 1623621585
transform 1 0 27232 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_206_286
timestamp 1623621585
transform 1 0 27416 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input460
timestamp 1623621585
transform 1 0 27968 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input462
timestamp 1623621585
transform 1 0 28612 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input463
timestamp 1623621585
transform 1 0 29256 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_295
timestamp 1623621585
transform 1 0 28244 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_302
timestamp 1623621585
transform 1 0 28888 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_309
timestamp 1623621585
transform 1 0 29532 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input465
timestamp 1623621585
transform 1 0 29900 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input467
timestamp 1623621585
transform 1 0 30544 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input469
timestamp 1623621585
transform 1 0 31188 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_206_316
timestamp 1623621585
transform 1 0 30176 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_323
timestamp 1623621585
transform 1 0 30820 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_330
timestamp 1623621585
transform 1 0 31464 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1878
timestamp 1623621585
transform 1 0 32568 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1623621585
transform 1 0 31924 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output704
timestamp 1623621585
transform 1 0 33396 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_206_334
timestamp 1623621585
transform 1 0 31832 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_206_338
timestamp 1623621585
transform 1 0 32200 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_206_343
timestamp 1623621585
transform 1 0 32660 0 -1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output681
timestamp 1623621585
transform 1 0 35604 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output689
timestamp 1623621585
transform 1 0 34868 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output698
timestamp 1623621585
transform 1 0 34132 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_355
timestamp 1623621585
transform 1 0 33764 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_363
timestamp 1623621585
transform 1 0 34500 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_371
timestamp 1623621585
transform 1 0 35236 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1623621585
transform 1 0 37076 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output668
timestamp 1623621585
transform 1 0 36340 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_379
timestamp 1623621585
transform 1 0 35972 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_387
timestamp 1623621585
transform 1 0 36708 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_206_395
timestamp 1623621585
transform 1 0 37444 0 -1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_413
timestamp 1623621585
transform -1 0 38824 0 -1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1879
timestamp 1623621585
transform 1 0 37812 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_206_400
timestamp 1623621585
transform 1 0 37904 0 -1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_206_406
timestamp 1623621585
transform 1 0 38456 0 -1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_414
timestamp 1623621585
transform 1 0 1104 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output674
timestamp 1623621585
transform 1 0 1748 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output676
timestamp 1623621585
transform 1 0 2484 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_3
timestamp 1623621585
transform 1 0 1380 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_11
timestamp 1623621585
transform 1 0 2116 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_19
timestamp 1623621585
transform 1 0 2852 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _0850_
timestamp 1623621585
transform 1 0 4232 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0852_
timestamp 1623621585
transform 1 0 4876 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1880
timestamp 1623621585
transform 1 0 3772 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_207_27
timestamp 1623621585
transform 1 0 3588 0 1 114784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_207_30
timestamp 1623621585
transform 1 0 3864 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_37
timestamp 1623621585
transform 1 0 4508 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0854_
timestamp 1623621585
transform 1 0 6256 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output626
timestamp 1623621585
transform 1 0 5520 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_44
timestamp 1623621585
transform 1 0 5152 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_52
timestamp 1623621585
transform 1 0 5888 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_59
timestamp 1623621585
transform 1 0 6532 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0855_
timestamp 1623621585
transform 1 0 6900 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output630
timestamp 1623621585
transform 1 0 7912 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_66
timestamp 1623621585
transform 1 0 7176 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_207_78
timestamp 1623621585
transform 1 0 8280 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _0878_
timestamp 1623621585
transform 1 0 9476 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0879_
timestamp 1623621585
transform 1 0 10120 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1881
timestamp 1623621585
transform 1 0 9016 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_87
timestamp 1623621585
transform 1 0 9108 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_94
timestamp 1623621585
transform 1 0 9752 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_101
timestamp 1623621585
transform 1 0 10396 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0880_
timestamp 1623621585
transform 1 0 10764 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0881_
timestamp 1623621585
transform 1 0 11408 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1623621585
transform 1 0 12052 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_108
timestamp 1623621585
transform 1 0 11040 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_115
timestamp 1623621585
transform 1 0 11684 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_122
timestamp 1623621585
transform 1 0 12328 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0884_
timestamp 1623621585
transform 1 0 12788 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0885_
timestamp 1623621585
transform 1 0 13432 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1882
timestamp 1623621585
transform 1 0 14260 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_207_126
timestamp 1623621585
transform 1 0 12696 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_130
timestamp 1623621585
transform 1 0 13064 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_207_137
timestamp 1623621585
transform 1 0 13708 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_207_144
timestamp 1623621585
transform 1 0 14352 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0886_
timestamp 1623621585
transform 1 0 14720 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0887_
timestamp 1623621585
transform 1 0 15364 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0888_
timestamp 1623621585
transform 1 0 16008 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_151
timestamp 1623621585
transform 1 0 14996 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_158
timestamp 1623621585
transform 1 0 15640 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_165
timestamp 1623621585
transform 1 0 16284 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0889_
timestamp 1623621585
transform 1 0 16652 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0891_
timestamp 1623621585
transform 1 0 17296 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0892_
timestamp 1623621585
transform 1 0 17940 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_172
timestamp 1623621585
transform 1 0 16928 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_179
timestamp 1623621585
transform 1 0 17572 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_186
timestamp 1623621585
transform 1 0 18216 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0893_
timestamp 1623621585
transform 1 0 18584 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0894_
timestamp 1623621585
transform 1 0 19964 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1883
timestamp 1623621585
transform 1 0 19504 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_207_193
timestamp 1623621585
transform 1 0 18860 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_207_199
timestamp 1623621585
transform 1 0 19412 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_201
timestamp 1623621585
transform 1 0 19596 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_208
timestamp 1623621585
transform 1 0 20240 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0862_
timestamp 1623621585
transform 1 0 21436 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1623621585
transform 1 0 20608 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0963_
timestamp 1623621585
transform 1 0 22080 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_207_215
timestamp 1623621585
transform 1 0 20884 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_207_224
timestamp 1623621585
transform 1 0 21712 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 1623621585
transform 1 0 24104 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1623621585
transform 1 0 22724 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1623621585
transform 1 0 23368 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_231
timestamp 1623621585
transform 1 0 22356 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_238
timestamp 1623621585
transform 1 0 23000 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_245
timestamp 1623621585
transform 1 0 23644 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_249
timestamp 1623621585
transform 1 0 24012 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _0895_
timestamp 1623621585
transform 1 0 25208 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0896_
timestamp 1623621585
transform 1 0 25852 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1884
timestamp 1623621585
transform 1 0 24748 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_253
timestamp 1623621585
transform 1 0 24380 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_258
timestamp 1623621585
transform 1 0 24840 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_265
timestamp 1623621585
transform 1 0 25484 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1623621585
transform 1 0 26496 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output713
timestamp 1623621585
transform 1 0 27600 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_272
timestamp 1623621585
transform 1 0 26128 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_279
timestamp 1623621585
transform 1 0 26772 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_207_287
timestamp 1623621585
transform 1 0 27508 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input459
timestamp 1623621585
transform 1 0 28336 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input461
timestamp 1623621585
transform 1 0 28980 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_292
timestamp 1623621585
transform 1 0 27968 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_299
timestamp 1623621585
transform 1 0 28612 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_306
timestamp 1623621585
transform 1 0 29256 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1885
timestamp 1623621585
transform 1 0 29992 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1623621585
transform 1 0 31740 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1623621585
transform 1 0 31096 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input464
timestamp 1623621585
transform 1 0 30452 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_207_315
timestamp 1623621585
transform 1 0 30084 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_322
timestamp 1623621585
transform 1 0 30728 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_329
timestamp 1623621585
transform 1 0 31372 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1623621585
transform 1 0 32384 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output699
timestamp 1623621585
transform 1 0 33028 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_336
timestamp 1623621585
transform 1 0 32016 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_343
timestamp 1623621585
transform 1 0 32660 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_351
timestamp 1623621585
transform 1 0 33396 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1886
timestamp 1623621585
transform 1 0 35236 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output683
timestamp 1623621585
transform 1 0 34500 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output690
timestamp 1623621585
transform 1 0 33764 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_359
timestamp 1623621585
transform 1 0 34132 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_367
timestamp 1623621585
transform 1 0 34868 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_207_372
timestamp 1623621585
transform 1 0 35328 0 1 114784
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output650
timestamp 1623621585
transform 1 0 36892 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output656
timestamp 1623621585
transform 1 0 36156 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_207_380
timestamp 1623621585
transform 1 0 36064 0 1 114784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_207_385
timestamp 1623621585
transform 1 0 36524 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_207_393
timestamp 1623621585
transform 1 0 37260 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_415
timestamp 1623621585
transform -1 0 38824 0 1 114784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input72
timestamp 1623621585
transform 1 0 37628 0 1 114784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_207_403
timestamp 1623621585
transform 1 0 38180 0 1 114784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_416
timestamp 1623621585
transform 1 0 1104 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output661
timestamp 1623621585
transform 1 0 1748 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output678
timestamp 1623621585
transform 1 0 2484 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_3
timestamp 1623621585
transform 1 0 1380 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_11
timestamp 1623621585
transform 1 0 2116 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_208_19
timestamp 1623621585
transform 1 0 2852 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output615
timestamp 1623621585
transform 1 0 4232 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output624
timestamp 1623621585
transform 1 0 3496 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_208_25
timestamp 1623621585
transform 1 0 3404 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_30
timestamp 1623621585
transform 1 0 3864 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_38
timestamp 1623621585
transform 1 0 4600 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0856_
timestamp 1623621585
transform 1 0 6808 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1887
timestamp 1623621585
transform 1 0 6348 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output625
timestamp 1623621585
transform 1 0 4968 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_46
timestamp 1623621585
transform 1 0 5336 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_208_54
timestamp 1623621585
transform 1 0 6072 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_58
timestamp 1623621585
transform 1 0 6440 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output629
timestamp 1623621585
transform 1 0 8096 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_65
timestamp 1623621585
transform 1 0 7084 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_208_73
timestamp 1623621585
transform 1 0 7820 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_80
timestamp 1623621585
transform 1 0 8464 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0831_
timestamp 1623621585
transform 1 0 8832 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0833_
timestamp 1623621585
transform 1 0 9476 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0834_
timestamp 1623621585
transform 1 0 10120 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_87
timestamp 1623621585
transform 1 0 9108 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_94
timestamp 1623621585
transform 1 0 9752 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_101
timestamp 1623621585
transform 1 0 10396 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0835_
timestamp 1623621585
transform 1 0 10764 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0882_
timestamp 1623621585
transform 1 0 12052 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1888
timestamp 1623621585
transform 1 0 11592 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_208_108
timestamp 1623621585
transform 1 0 11040 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_208_115
timestamp 1623621585
transform 1 0 11684 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_122
timestamp 1623621585
transform 1 0 12328 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0839_
timestamp 1623621585
transform 1 0 13340 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0883_
timestamp 1623621585
transform 1 0 12696 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_129
timestamp 1623621585
transform 1 0 12972 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_136
timestamp 1623621585
transform 1 0 13616 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_208_144
timestamp 1623621585
transform 1 0 14352 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _0841_
timestamp 1623621585
transform 1 0 14536 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0842_
timestamp 1623621585
transform 1 0 15180 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0843_
timestamp 1623621585
transform 1 0 15824 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_149
timestamp 1623621585
transform 1 0 14812 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_156
timestamp 1623621585
transform 1 0 15456 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_163
timestamp 1623621585
transform 1 0 16100 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _0890_
timestamp 1623621585
transform 1 0 17296 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1889
timestamp 1623621585
transform 1 0 16836 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_172
timestamp 1623621585
transform 1 0 16928 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_179
timestamp 1623621585
transform 1 0 17572 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_208_187
timestamp 1623621585
transform 1 0 18308 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _0847_
timestamp 1623621585
transform 1 0 18400 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0848_
timestamp 1623621585
transform 1 0 19044 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0859_
timestamp 1623621585
transform 1 0 19688 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_191
timestamp 1623621585
transform 1 0 18676 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_198
timestamp 1623621585
transform 1 0 19320 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_205
timestamp 1623621585
transform 1 0 19964 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0860_
timestamp 1623621585
transform 1 0 20332 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0861_
timestamp 1623621585
transform 1 0 20976 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1890
timestamp 1623621585
transform 1 0 22080 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_212
timestamp 1623621585
transform 1 0 20608 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_219
timestamp 1623621585
transform 1 0 21252 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_208_227
timestamp 1623621585
transform 1 0 21988 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_229
timestamp 1623621585
transform 1 0 22172 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0863_
timestamp 1623621585
transform 1 0 22540 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0864_
timestamp 1623621585
transform 1 0 23184 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0865_
timestamp 1623621585
transform 1 0 23828 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_208_236
timestamp 1623621585
transform 1 0 22816 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_243
timestamp 1623621585
transform 1 0 23460 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_250
timestamp 1623621585
transform 1 0 24104 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0866_
timestamp 1623621585
transform 1 0 24472 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0868_
timestamp 1623621585
transform 1 0 25300 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_208_257
timestamp 1623621585
transform 1 0 24748 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_208_266
timestamp 1623621585
transform 1 0 25576 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1891
timestamp 1623621585
transform 1 0 27324 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output707
timestamp 1623621585
transform 1 0 26312 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output711
timestamp 1623621585
transform 1 0 27784 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_208_278
timestamp 1623621585
transform 1 0 26680 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_284
timestamp 1623621585
transform 1 0 27232 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_286
timestamp 1623621585
transform 1 0 27416 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 1623621585
transform 1 0 28520 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output714
timestamp 1623621585
transform 1 0 29440 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_294
timestamp 1623621585
transform 1 0 28152 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_208_301
timestamp 1623621585
transform 1 0 28796 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_307
timestamp 1623621585
transform 1 0 29348 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_208_312
timestamp 1623621585
transform 1 0 29808 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1623621585
transform 1 0 31556 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1623621585
transform 1 0 30912 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output715
timestamp 1623621585
transform 1 0 30176 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_320
timestamp 1623621585
transform 1 0 30544 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_327
timestamp 1623621585
transform 1 0 31188 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1892
timestamp 1623621585
transform 1 0 32568 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output686
timestamp 1623621585
transform 1 0 33580 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_334
timestamp 1623621585
transform 1 0 31832 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_208_343
timestamp 1623621585
transform 1 0 32660 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_208_351
timestamp 1623621585
transform 1 0 33396 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output673
timestamp 1623621585
transform 1 0 35052 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output682
timestamp 1623621585
transform 1 0 34316 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_357
timestamp 1623621585
transform 1 0 33948 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_365
timestamp 1623621585
transform 1 0 34684 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_373
timestamp 1623621585
transform 1 0 35420 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output644
timestamp 1623621585
transform 1 0 35788 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output645
timestamp 1623621585
transform 1 0 36524 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_208_381
timestamp 1623621585
transform 1 0 36156 0 -1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_208_389
timestamp 1623621585
transform 1 0 36892 0 -1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_417
timestamp 1623621585
transform -1 0 38824 0 -1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1893
timestamp 1623621585
transform 1 0 37812 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_208_397
timestamp 1623621585
transform 1 0 37628 0 -1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_208_400
timestamp 1623621585
transform 1 0 37904 0 -1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_208_406
timestamp 1623621585
transform 1 0 38456 0 -1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_418
timestamp 1623621585
transform 1 0 1104 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output593
timestamp 1623621585
transform 1 0 2208 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output604
timestamp 1623621585
transform 1 0 2944 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_3
timestamp 1623621585
transform 1 0 1380 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_209_11
timestamp 1623621585
transform 1 0 2116 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_16
timestamp 1623621585
transform 1 0 2576 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1894
timestamp 1623621585
transform 1 0 3772 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output588
timestamp 1623621585
transform 1 0 4692 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_24
timestamp 1623621585
transform 1 0 3312 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_28
timestamp 1623621585
transform 1 0 3680 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_209_30
timestamp 1623621585
transform 1 0 3864 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_209_38
timestamp 1623621585
transform 1 0 4600 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output587
timestamp 1623621585
transform 1 0 5428 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output589
timestamp 1623621585
transform 1 0 6164 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_43
timestamp 1623621585
transform 1 0 5060 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_51
timestamp 1623621585
transform 1 0 5796 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_59
timestamp 1623621585
transform 1 0 6532 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output627
timestamp 1623621585
transform 1 0 6900 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output628
timestamp 1623621585
transform 1 0 7636 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_67
timestamp 1623621585
transform 1 0 7268 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_75
timestamp 1623621585
transform 1 0 8004 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_209_83
timestamp 1623621585
transform 1 0 8740 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0832_
timestamp 1623621585
transform 1 0 9476 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1895
timestamp 1623621585
transform 1 0 9016 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output597
timestamp 1623621585
transform 1 0 10396 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_87
timestamp 1623621585
transform 1 0 9108 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_94
timestamp 1623621585
transform 1 0 9752 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_100
timestamp 1623621585
transform 1 0 10304 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _0836_
timestamp 1623621585
transform 1 0 11868 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0837_
timestamp 1623621585
transform 1 0 12512 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output598
timestamp 1623621585
transform 1 0 11132 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_105
timestamp 1623621585
transform 1 0 10764 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_113
timestamp 1623621585
transform 1 0 11500 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_120
timestamp 1623621585
transform 1 0 12144 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0838_
timestamp 1623621585
transform 1 0 13156 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1896
timestamp 1623621585
transform 1 0 14260 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_127
timestamp 1623621585
transform 1 0 12788 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_134
timestamp 1623621585
transform 1 0 13432 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_209_142
timestamp 1623621585
transform 1 0 14168 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_144
timestamp 1623621585
transform 1 0 14352 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0840_
timestamp 1623621585
transform 1 0 14720 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output606
timestamp 1623621585
transform 1 0 15548 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output607
timestamp 1623621585
transform 1 0 16284 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_151
timestamp 1623621585
transform 1 0 14996 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_209_161
timestamp 1623621585
transform 1 0 15916 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0844_
timestamp 1623621585
transform 1 0 17020 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0845_
timestamp 1623621585
transform 1 0 17664 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _0846_
timestamp 1623621585
transform 1 0 18308 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_209_169
timestamp 1623621585
transform 1 0 16652 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_176
timestamp 1623621585
transform 1 0 17296 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_183
timestamp 1623621585
transform 1 0 17940 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1897
timestamp 1623621585
transform 1 0 19504 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output613
timestamp 1623621585
transform 1 0 19964 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_190
timestamp 1623621585
transform 1 0 18584 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_198
timestamp 1623621585
transform 1 0 19320 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_209_201
timestamp 1623621585
transform 1 0 19596 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output616
timestamp 1623621585
transform 1 0 21252 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output617
timestamp 1623621585
transform 1 0 21988 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_209
timestamp 1623621585
transform 1 0 20332 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_209_217
timestamp 1623621585
transform 1 0 21068 0 1 115872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_209_223
timestamp 1623621585
transform 1 0 21620 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output619
timestamp 1623621585
transform 1 0 23092 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output620
timestamp 1623621585
transform 1 0 23828 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_231
timestamp 1623621585
transform 1 0 22356 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_209_243
timestamp 1623621585
transform 1 0 23460 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0867_
timestamp 1623621585
transform 1 0 25208 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1898
timestamp 1623621585
transform 1 0 24748 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output705
timestamp 1623621585
transform 1 0 25852 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_209_251
timestamp 1623621585
transform 1 0 24196 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_209_258
timestamp 1623621585
transform 1 0 24840 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_265
timestamp 1623621585
transform 1 0 25484 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0774_
timestamp 1623621585
transform 1 0 26588 0 1 115872
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output708
timestamp 1623621585
transform 1 0 27416 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_273
timestamp 1623621585
transform 1 0 26220 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_282
timestamp 1623621585
transform 1 0 27048 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_290
timestamp 1623621585
transform 1 0 27784 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output710
timestamp 1623621585
transform 1 0 28152 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output712
timestamp 1623621585
transform 1 0 28888 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_298
timestamp 1623621585
transform 1 0 28520 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_306
timestamp 1623621585
transform 1 0 29256 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0772_
timestamp 1623621585
transform 1 0 30452 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0775_
timestamp 1623621585
transform 1 0 31648 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1899
timestamp 1623621585
transform 1 0 29992 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_315
timestamp 1623621585
transform 1 0 30084 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_328
timestamp 1623621585
transform 1 0 31280 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0777_
timestamp 1623621585
transform 1 0 32844 0 1 115872
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_209_341
timestamp 1623621585
transform 1 0 32476 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_354
timestamp 1623621585
transform 1 0 33672 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1900
timestamp 1623621585
transform 1 0 35236 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output658
timestamp 1623621585
transform 1 0 34500 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_209_362
timestamp 1623621585
transform 1 0 34408 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_367
timestamp 1623621585
transform 1 0 34868 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_372
timestamp 1623621585
transform 1 0 35328 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output641
timestamp 1623621585
transform 1 0 35696 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output643
timestamp 1623621585
transform 1 0 36432 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_209_380
timestamp 1623621585
transform 1 0 36064 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_209_388
timestamp 1623621585
transform 1 0 36800 0 1 115872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_419
timestamp 1623621585
transform -1 0 38824 0 1 115872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1623621585
transform 1 0 37628 0 1 115872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_209_396
timestamp 1623621585
transform 1 0 37536 0 1 115872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_209_403
timestamp 1623621585
transform 1 0 38180 0 1 115872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_420
timestamp 1623621585
transform 1 0 1104 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output553
timestamp 1623621585
transform 1 0 1748 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output555
timestamp 1623621585
transform 1 0 2484 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_3
timestamp 1623621585
transform 1 0 1380 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_11
timestamp 1623621585
transform 1 0 2116 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_19
timestamp 1623621585
transform 1 0 2852 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output549
timestamp 1623621585
transform 1 0 3220 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output566
timestamp 1623621585
transform 1 0 3956 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output577
timestamp 1623621585
transform 1 0 4692 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_27
timestamp 1623621585
transform 1 0 3588 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_35
timestamp 1623621585
transform 1 0 4324 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1901
timestamp 1623621585
transform 1 0 6348 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output586
timestamp 1623621585
transform 1 0 5428 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output590
timestamp 1623621585
transform 1 0 6808 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_43
timestamp 1623621585
transform 1 0 5060 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_210_51
timestamp 1623621585
transform 1 0 5796 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_210_58
timestamp 1623621585
transform 1 0 6440 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output591
timestamp 1623621585
transform 1 0 7544 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output592
timestamp 1623621585
transform 1 0 8280 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_66
timestamp 1623621585
transform 1 0 7176 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_74
timestamp 1623621585
transform 1 0 7912 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_82
timestamp 1623621585
transform 1 0 8648 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output594
timestamp 1623621585
transform 1 0 9016 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output595
timestamp 1623621585
transform 1 0 9752 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output596
timestamp 1623621585
transform 1 0 10488 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_90
timestamp 1623621585
transform 1 0 9384 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_98
timestamp 1623621585
transform 1 0 10120 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1902
timestamp 1623621585
transform 1 0 11592 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output599
timestamp 1623621585
transform 1 0 12052 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_106
timestamp 1623621585
transform 1 0 10856 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_210_115
timestamp 1623621585
transform 1 0 11684 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_123
timestamp 1623621585
transform 1 0 12420 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output600
timestamp 1623621585
transform 1 0 12788 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output601
timestamp 1623621585
transform 1 0 13524 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output602
timestamp 1623621585
transform 1 0 14260 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_131
timestamp 1623621585
transform 1 0 13156 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_139
timestamp 1623621585
transform 1 0 13892 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output603
timestamp 1623621585
transform 1 0 14996 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output605
timestamp 1623621585
transform 1 0 15732 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_147
timestamp 1623621585
transform 1 0 14628 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_155
timestamp 1623621585
transform 1 0 15364 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_163
timestamp 1623621585
transform 1 0 16100 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1903
timestamp 1623621585
transform 1 0 16836 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output608
timestamp 1623621585
transform 1 0 17296 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output609
timestamp 1623621585
transform 1 0 18032 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_172
timestamp 1623621585
transform 1 0 16928 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_180
timestamp 1623621585
transform 1 0 17664 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output610
timestamp 1623621585
transform 1 0 18768 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output611
timestamp 1623621585
transform 1 0 19504 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output612
timestamp 1623621585
transform 1 0 20240 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_188
timestamp 1623621585
transform 1 0 18400 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_196
timestamp 1623621585
transform 1 0 19136 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_204
timestamp 1623621585
transform 1 0 19872 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1904
timestamp 1623621585
transform 1 0 22080 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output614
timestamp 1623621585
transform 1 0 20976 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_212
timestamp 1623621585
transform 1 0 20608 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_210_220
timestamp 1623621585
transform 1 0 21344 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_210_229
timestamp 1623621585
transform 1 0 22172 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output580
timestamp 1623621585
transform 1 0 22540 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output618
timestamp 1623621585
transform 1 0 23276 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_237
timestamp 1623621585
transform 1 0 22908 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_210_245
timestamp 1623621585
transform 1 0 23644 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output583
timestamp 1623621585
transform 1 0 24196 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output621
timestamp 1623621585
transform 1 0 24932 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output622
timestamp 1623621585
transform 1 0 25668 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_255
timestamp 1623621585
transform 1 0 24564 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_263
timestamp 1623621585
transform 1 0 25300 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1905
timestamp 1623621585
transform 1 0 27324 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output623
timestamp 1623621585
transform 1 0 26404 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output706
timestamp 1623621585
transform 1 0 27784 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_271
timestamp 1623621585
transform 1 0 26036 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_210_279
timestamp 1623621585
transform 1 0 26772 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_210_286
timestamp 1623621585
transform 1 0 27416 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0773_
timestamp 1623621585
transform 1 0 29256 0 -1 116960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output709
timestamp 1623621585
transform 1 0 28520 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_294
timestamp 1623621585
transform 1 0 28152 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_302
timestamp 1623621585
transform 1 0 28888 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0776_
timestamp 1623621585
transform 1 0 30912 0 -1 116960
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_210_315
timestamp 1623621585
transform 1 0 30084 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_210_323
timestamp 1623621585
transform 1 0 30820 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_210_333
timestamp 1623621585
transform 1 0 31740 0 -1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1906
timestamp 1623621585
transform 1 0 32568 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output679
timestamp 1623621585
transform 1 0 33120 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_210_341
timestamp 1623621585
transform 1 0 32476 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_343
timestamp 1623621585
transform 1 0 32660 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_210_347
timestamp 1623621585
transform 1 0 33028 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_210_352
timestamp 1623621585
transform 1 0 33488 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output638
timestamp 1623621585
transform 1 0 34592 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output639
timestamp 1623621585
transform 1 0 35328 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output677
timestamp 1623621585
transform 1 0 33856 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_360
timestamp 1623621585
transform 1 0 34224 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_368
timestamp 1623621585
transform 1 0 34960 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output640
timestamp 1623621585
transform 1 0 36064 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output642
timestamp 1623621585
transform 1 0 36800 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_376
timestamp 1623621585
transform 1 0 35696 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_210_384
timestamp 1623621585
transform 1 0 36432 0 -1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_210_392
timestamp 1623621585
transform 1 0 37168 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_421
timestamp 1623621585
transform -1 0 38824 0 -1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1907
timestamp 1623621585
transform 1 0 37812 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_210_398
timestamp 1623621585
transform 1 0 37720 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_210_400
timestamp 1623621585
transform 1 0 37904 0 -1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_210_406
timestamp 1623621585
transform 1 0 38456 0 -1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_422
timestamp 1623621585
transform 1 0 1104 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output547
timestamp 1623621585
transform 1 0 1748 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output548
timestamp 1623621585
transform 1 0 2484 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_3
timestamp 1623621585
transform 1 0 1380 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_11
timestamp 1623621585
transform 1 0 2116 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_211_19
timestamp 1623621585
transform 1 0 2852 0 1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1908
timestamp 1623621585
transform 1 0 3772 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output550
timestamp 1623621585
transform 1 0 4232 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_211_27
timestamp 1623621585
transform 1 0 3588 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_211_30
timestamp 1623621585
transform 1 0 3864 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_38
timestamp 1623621585
transform 1 0 4600 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1909
timestamp 1623621585
transform 1 0 6440 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output551
timestamp 1623621585
transform 1 0 4968 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output552
timestamp 1623621585
transform 1 0 5704 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_46
timestamp 1623621585
transform 1 0 5336 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_54
timestamp 1623621585
transform 1 0 6072 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_59
timestamp 1623621585
transform 1 0 6532 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _0858_
timestamp 1623621585
transform 1 0 7636 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output554
timestamp 1623621585
transform 1 0 6900 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output556
timestamp 1623621585
transform 1 0 8280 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_67
timestamp 1623621585
transform 1 0 7268 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_74
timestamp 1623621585
transform 1 0 7912 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_82
timestamp 1623621585
transform 1 0 8648 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1910
timestamp 1623621585
transform 1 0 9108 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output557
timestamp 1623621585
transform 1 0 9568 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output558
timestamp 1623621585
transform 1 0 10304 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_86
timestamp 1623621585
transform 1 0 9016 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_211_88
timestamp 1623621585
transform 1 0 9200 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_96
timestamp 1623621585
transform 1 0 9936 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_104
timestamp 1623621585
transform 1 0 10672 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1911
timestamp 1623621585
transform 1 0 11776 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output559
timestamp 1623621585
transform 1 0 11040 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output560
timestamp 1623621585
transform 1 0 12236 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_112
timestamp 1623621585
transform 1 0 11408 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_117
timestamp 1623621585
transform 1 0 11868 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_125
timestamp 1623621585
transform 1 0 12604 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1912
timestamp 1623621585
transform 1 0 14444 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output561
timestamp 1623621585
transform 1 0 12972 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output562
timestamp 1623621585
transform 1 0 13708 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_133
timestamp 1623621585
transform 1 0 13340 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_141
timestamp 1623621585
transform 1 0 14076 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output563
timestamp 1623621585
transform 1 0 14904 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output564
timestamp 1623621585
transform 1 0 15640 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output565
timestamp 1623621585
transform 1 0 16376 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_146
timestamp 1623621585
transform 1 0 14536 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_154
timestamp 1623621585
transform 1 0 15272 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_162
timestamp 1623621585
transform 1 0 16008 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1913
timestamp 1623621585
transform 1 0 17112 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output567
timestamp 1623621585
transform 1 0 17572 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output568
timestamp 1623621585
transform 1 0 18308 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_170
timestamp 1623621585
transform 1 0 16744 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_175
timestamp 1623621585
transform 1 0 17204 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_183
timestamp 1623621585
transform 1 0 17940 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1914
timestamp 1623621585
transform 1 0 19780 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output569
timestamp 1623621585
transform 1 0 19044 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output570
timestamp 1623621585
transform 1 0 20240 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_191
timestamp 1623621585
transform 1 0 18676 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_199
timestamp 1623621585
transform 1 0 19412 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_204
timestamp 1623621585
transform 1 0 19872 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output571
timestamp 1623621585
transform 1 0 20976 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output572
timestamp 1623621585
transform 1 0 21712 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_212
timestamp 1623621585
transform 1 0 20608 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_220
timestamp 1623621585
transform 1 0 21344 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_228
timestamp 1623621585
transform 1 0 22080 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1915
timestamp 1623621585
transform 1 0 22448 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output573
timestamp 1623621585
transform 1 0 22908 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output574
timestamp 1623621585
transform 1 0 23644 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_233
timestamp 1623621585
transform 1 0 22540 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_241
timestamp 1623621585
transform 1 0 23276 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_249
timestamp 1623621585
transform 1 0 24012 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1916
timestamp 1623621585
transform 1 0 25116 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output575
timestamp 1623621585
transform 1 0 24380 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output576
timestamp 1623621585
transform 1 0 25576 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_257
timestamp 1623621585
transform 1 0 24748 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_262
timestamp 1623621585
transform 1 0 25208 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_270
timestamp 1623621585
transform 1 0 25944 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1917
timestamp 1623621585
transform 1 0 27784 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output578
timestamp 1623621585
transform 1 0 26312 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output579
timestamp 1623621585
transform 1 0 27048 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_278
timestamp 1623621585
transform 1 0 26680 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_286
timestamp 1623621585
transform 1 0 27416 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_291
timestamp 1623621585
transform 1 0 27876 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output581
timestamp 1623621585
transform 1 0 28244 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output582
timestamp 1623621585
transform 1 0 28980 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output584
timestamp 1623621585
transform 1 0 29716 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_299
timestamp 1623621585
transform 1 0 28612 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_307
timestamp 1623621585
transform 1 0 29348 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1918
timestamp 1623621585
transform 1 0 30452 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output585
timestamp 1623621585
transform 1 0 30912 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output637
timestamp 1623621585
transform 1 0 31648 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_315
timestamp 1623621585
transform 1 0 30084 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_320
timestamp 1623621585
transform 1 0 30544 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_328
timestamp 1623621585
transform 1 0 31280 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1919
timestamp 1623621585
transform 1 0 33120 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output636
timestamp 1623621585
transform 1 0 32384 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_336
timestamp 1623621585
transform 1 0 32016 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_211_344
timestamp 1623621585
transform 1 0 32752 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_211_349
timestamp 1623621585
transform 1 0 33212 0 1 116960
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output634
timestamp 1623621585
transform 1 0 34132 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output635
timestamp 1623621585
transform 1 0 35052 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_211_357
timestamp 1623621585
transform 1 0 33948 0 1 116960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_211_363
timestamp 1623621585
transform 1 0 34500 0 1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_211_373
timestamp 1623621585
transform 1 0 35420 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1920
timestamp 1623621585
transform 1 0 35788 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  input68
timestamp 1623621585
transform 1 0 36340 0 1 116960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input71
timestamp 1623621585
transform 1 0 37260 0 1 116960
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_211_378
timestamp 1623621585
transform 1 0 35880 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_211_382
timestamp 1623621585
transform 1 0 36248 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_211_389
timestamp 1623621585
transform 1 0 36892 0 1 116960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_423
timestamp 1623621585
transform -1 0 38824 0 1 116960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1921
timestamp 1623621585
transform 1 0 38456 0 1 116960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_211_402
timestamp 1623621585
transform 1 0 38088 0 1 116960
box -38 -48 406 592
<< labels >>
rlabel metal2 s 110 119200 166 120800 6 dsi[0]
port 0 nsew signal tristate
rlabel metal2 s 294 119200 350 120800 6 dsi[1]
port 1 nsew signal tristate
rlabel metal2 s 478 119200 534 120800 6 dsi[2]
port 2 nsew signal tristate
rlabel metal2 s 662 119200 718 120800 6 dsi[3]
port 3 nsew signal tristate
rlabel metal2 s 938 119200 994 120800 6 dsi[4]
port 4 nsew signal tristate
rlabel metal2 s 1122 119200 1178 120800 6 dsi[5]
port 5 nsew signal tristate
rlabel metal2 s 1306 119200 1362 120800 6 dsi[6]
port 6 nsew signal tristate
rlabel metal2 s 1582 119200 1638 120800 6 dsi[7]
port 7 nsew signal tristate
rlabel metal2 s 1766 119200 1822 120800 6 io_in[0]
port 8 nsew signal input
rlabel metal2 s 8114 119200 8170 120800 6 io_in[10]
port 9 nsew signal input
rlabel metal2 s 8758 119200 8814 120800 6 io_in[11]
port 10 nsew signal input
rlabel metal2 s 9402 119200 9458 120800 6 io_in[12]
port 11 nsew signal input
rlabel metal2 s 10046 119200 10102 120800 6 io_in[13]
port 12 nsew signal input
rlabel metal2 s 10690 119200 10746 120800 6 io_in[14]
port 13 nsew signal input
rlabel metal2 s 11242 119200 11298 120800 6 io_in[15]
port 14 nsew signal input
rlabel metal2 s 11886 119200 11942 120800 6 io_in[16]
port 15 nsew signal input
rlabel metal2 s 12530 119200 12586 120800 6 io_in[17]
port 16 nsew signal input
rlabel metal2 s 13174 119200 13230 120800 6 io_in[18]
port 17 nsew signal input
rlabel metal2 s 13818 119200 13874 120800 6 io_in[19]
port 18 nsew signal input
rlabel metal2 s 2410 119200 2466 120800 6 io_in[1]
port 19 nsew signal input
rlabel metal2 s 14462 119200 14518 120800 6 io_in[20]
port 20 nsew signal input
rlabel metal2 s 15106 119200 15162 120800 6 io_in[21]
port 21 nsew signal input
rlabel metal2 s 15750 119200 15806 120800 6 io_in[22]
port 22 nsew signal input
rlabel metal2 s 16394 119200 16450 120800 6 io_in[23]
port 23 nsew signal input
rlabel metal2 s 17038 119200 17094 120800 6 io_in[24]
port 24 nsew signal input
rlabel metal2 s 17682 119200 17738 120800 6 io_in[25]
port 25 nsew signal input
rlabel metal2 s 18234 119200 18290 120800 6 io_in[26]
port 26 nsew signal input
rlabel metal2 s 18878 119200 18934 120800 6 io_in[27]
port 27 nsew signal input
rlabel metal2 s 19522 119200 19578 120800 6 io_in[28]
port 28 nsew signal input
rlabel metal2 s 20166 119200 20222 120800 6 io_in[29]
port 29 nsew signal input
rlabel metal2 s 3054 119200 3110 120800 6 io_in[2]
port 30 nsew signal input
rlabel metal2 s 20810 119200 20866 120800 6 io_in[30]
port 31 nsew signal input
rlabel metal2 s 21454 119200 21510 120800 6 io_in[31]
port 32 nsew signal input
rlabel metal2 s 22098 119200 22154 120800 6 io_in[32]
port 33 nsew signal input
rlabel metal2 s 22742 119200 22798 120800 6 io_in[33]
port 34 nsew signal input
rlabel metal2 s 23386 119200 23442 120800 6 io_in[34]
port 35 nsew signal input
rlabel metal2 s 24030 119200 24086 120800 6 io_in[35]
port 36 nsew signal input
rlabel metal2 s 24582 119200 24638 120800 6 io_in[36]
port 37 nsew signal input
rlabel metal2 s 25226 119200 25282 120800 6 io_in[37]
port 38 nsew signal input
rlabel metal2 s 3698 119200 3754 120800 6 io_in[3]
port 39 nsew signal input
rlabel metal2 s 4342 119200 4398 120800 6 io_in[4]
port 40 nsew signal input
rlabel metal2 s 4894 119200 4950 120800 6 io_in[5]
port 41 nsew signal input
rlabel metal2 s 5538 119200 5594 120800 6 io_in[6]
port 42 nsew signal input
rlabel metal2 s 6182 119200 6238 120800 6 io_in[7]
port 43 nsew signal input
rlabel metal2 s 6826 119200 6882 120800 6 io_in[8]
port 44 nsew signal input
rlabel metal2 s 7470 119200 7526 120800 6 io_in[9]
port 45 nsew signal input
rlabel metal2 s 1950 119200 2006 120800 6 io_oeb[0]
port 46 nsew signal tristate
rlabel metal2 s 8298 119200 8354 120800 6 io_oeb[10]
port 47 nsew signal tristate
rlabel metal2 s 8942 119200 8998 120800 6 io_oeb[11]
port 48 nsew signal tristate
rlabel metal2 s 9586 119200 9642 120800 6 io_oeb[12]
port 49 nsew signal tristate
rlabel metal2 s 10230 119200 10286 120800 6 io_oeb[13]
port 50 nsew signal tristate
rlabel metal2 s 10874 119200 10930 120800 6 io_oeb[14]
port 51 nsew signal tristate
rlabel metal2 s 11518 119200 11574 120800 6 io_oeb[15]
port 52 nsew signal tristate
rlabel metal2 s 12162 119200 12218 120800 6 io_oeb[16]
port 53 nsew signal tristate
rlabel metal2 s 12806 119200 12862 120800 6 io_oeb[17]
port 54 nsew signal tristate
rlabel metal2 s 13450 119200 13506 120800 6 io_oeb[18]
port 55 nsew signal tristate
rlabel metal2 s 14002 119200 14058 120800 6 io_oeb[19]
port 56 nsew signal tristate
rlabel metal2 s 2594 119200 2650 120800 6 io_oeb[1]
port 57 nsew signal tristate
rlabel metal2 s 14646 119200 14702 120800 6 io_oeb[20]
port 58 nsew signal tristate
rlabel metal2 s 15290 119200 15346 120800 6 io_oeb[21]
port 59 nsew signal tristate
rlabel metal2 s 15934 119200 15990 120800 6 io_oeb[22]
port 60 nsew signal tristate
rlabel metal2 s 16578 119200 16634 120800 6 io_oeb[23]
port 61 nsew signal tristate
rlabel metal2 s 17222 119200 17278 120800 6 io_oeb[24]
port 62 nsew signal tristate
rlabel metal2 s 17866 119200 17922 120800 6 io_oeb[25]
port 63 nsew signal tristate
rlabel metal2 s 18510 119200 18566 120800 6 io_oeb[26]
port 64 nsew signal tristate
rlabel metal2 s 19154 119200 19210 120800 6 io_oeb[27]
port 65 nsew signal tristate
rlabel metal2 s 19798 119200 19854 120800 6 io_oeb[28]
port 66 nsew signal tristate
rlabel metal2 s 20350 119200 20406 120800 6 io_oeb[29]
port 67 nsew signal tristate
rlabel metal2 s 3238 119200 3294 120800 6 io_oeb[2]
port 68 nsew signal tristate
rlabel metal2 s 20994 119200 21050 120800 6 io_oeb[30]
port 69 nsew signal tristate
rlabel metal2 s 21638 119200 21694 120800 6 io_oeb[31]
port 70 nsew signal tristate
rlabel metal2 s 22282 119200 22338 120800 6 io_oeb[32]
port 71 nsew signal tristate
rlabel metal2 s 22926 119200 22982 120800 6 io_oeb[33]
port 72 nsew signal tristate
rlabel metal2 s 23570 119200 23626 120800 6 io_oeb[34]
port 73 nsew signal tristate
rlabel metal2 s 24214 119200 24270 120800 6 io_oeb[35]
port 74 nsew signal tristate
rlabel metal2 s 24858 119200 24914 120800 6 io_oeb[36]
port 75 nsew signal tristate
rlabel metal2 s 25502 119200 25558 120800 6 io_oeb[37]
port 76 nsew signal tristate
rlabel metal2 s 3882 119200 3938 120800 6 io_oeb[3]
port 77 nsew signal tristate
rlabel metal2 s 4526 119200 4582 120800 6 io_oeb[4]
port 78 nsew signal tristate
rlabel metal2 s 5170 119200 5226 120800 6 io_oeb[5]
port 79 nsew signal tristate
rlabel metal2 s 5814 119200 5870 120800 6 io_oeb[6]
port 80 nsew signal tristate
rlabel metal2 s 6458 119200 6514 120800 6 io_oeb[7]
port 81 nsew signal tristate
rlabel metal2 s 7010 119200 7066 120800 6 io_oeb[8]
port 82 nsew signal tristate
rlabel metal2 s 7654 119200 7710 120800 6 io_oeb[9]
port 83 nsew signal tristate
rlabel metal2 s 2226 119200 2282 120800 6 io_out[0]
port 84 nsew signal tristate
rlabel metal2 s 8574 119200 8630 120800 6 io_out[10]
port 85 nsew signal tristate
rlabel metal2 s 9126 119200 9182 120800 6 io_out[11]
port 86 nsew signal tristate
rlabel metal2 s 9770 119200 9826 120800 6 io_out[12]
port 87 nsew signal tristate
rlabel metal2 s 10414 119200 10470 120800 6 io_out[13]
port 88 nsew signal tristate
rlabel metal2 s 11058 119200 11114 120800 6 io_out[14]
port 89 nsew signal tristate
rlabel metal2 s 11702 119200 11758 120800 6 io_out[15]
port 90 nsew signal tristate
rlabel metal2 s 12346 119200 12402 120800 6 io_out[16]
port 91 nsew signal tristate
rlabel metal2 s 12990 119200 13046 120800 6 io_out[17]
port 92 nsew signal tristate
rlabel metal2 s 13634 119200 13690 120800 6 io_out[18]
port 93 nsew signal tristate
rlabel metal2 s 14278 119200 14334 120800 6 io_out[19]
port 94 nsew signal tristate
rlabel metal2 s 2778 119200 2834 120800 6 io_out[1]
port 95 nsew signal tristate
rlabel metal2 s 14922 119200 14978 120800 6 io_out[20]
port 96 nsew signal tristate
rlabel metal2 s 15566 119200 15622 120800 6 io_out[21]
port 97 nsew signal tristate
rlabel metal2 s 16118 119200 16174 120800 6 io_out[22]
port 98 nsew signal tristate
rlabel metal2 s 16762 119200 16818 120800 6 io_out[23]
port 99 nsew signal tristate
rlabel metal2 s 17406 119200 17462 120800 6 io_out[24]
port 100 nsew signal tristate
rlabel metal2 s 18050 119200 18106 120800 6 io_out[25]
port 101 nsew signal tristate
rlabel metal2 s 18694 119200 18750 120800 6 io_out[26]
port 102 nsew signal tristate
rlabel metal2 s 19338 119200 19394 120800 6 io_out[27]
port 103 nsew signal tristate
rlabel metal2 s 19982 119200 20038 120800 6 io_out[28]
port 104 nsew signal tristate
rlabel metal2 s 20626 119200 20682 120800 6 io_out[29]
port 105 nsew signal tristate
rlabel metal2 s 3422 119200 3478 120800 6 io_out[2]
port 106 nsew signal tristate
rlabel metal2 s 21270 119200 21326 120800 6 io_out[30]
port 107 nsew signal tristate
rlabel metal2 s 21914 119200 21970 120800 6 io_out[31]
port 108 nsew signal tristate
rlabel metal2 s 22466 119200 22522 120800 6 io_out[32]
port 109 nsew signal tristate
rlabel metal2 s 23110 119200 23166 120800 6 io_out[33]
port 110 nsew signal tristate
rlabel metal2 s 23754 119200 23810 120800 6 io_out[34]
port 111 nsew signal tristate
rlabel metal2 s 24398 119200 24454 120800 6 io_out[35]
port 112 nsew signal tristate
rlabel metal2 s 25042 119200 25098 120800 6 io_out[36]
port 113 nsew signal tristate
rlabel metal2 s 25686 119200 25742 120800 6 io_out[37]
port 114 nsew signal tristate
rlabel metal2 s 4066 119200 4122 120800 6 io_out[3]
port 115 nsew signal tristate
rlabel metal2 s 4710 119200 4766 120800 6 io_out[4]
port 116 nsew signal tristate
rlabel metal2 s 5354 119200 5410 120800 6 io_out[5]
port 117 nsew signal tristate
rlabel metal2 s 5998 119200 6054 120800 6 io_out[6]
port 118 nsew signal tristate
rlabel metal2 s 6642 119200 6698 120800 6 io_out[7]
port 119 nsew signal tristate
rlabel metal2 s 7286 119200 7342 120800 6 io_out[8]
port 120 nsew signal tristate
rlabel metal2 s 7930 119200 7986 120800 6 io_out[9]
port 121 nsew signal tristate
rlabel metal2 s 662 -800 718 800 8 irq[0]
port 122 nsew signal tristate
rlabel metal2 s 938 -800 994 800 8 irq[1]
port 123 nsew signal tristate
rlabel metal2 s 1214 -800 1270 800 8 irq[2]
port 124 nsew signal tristate
rlabel metal2 s 31942 -800 31998 800 8 la_reset[0]
port 125 nsew signal input
rlabel metal2 s 34794 -800 34850 800 8 la_reset[10]
port 126 nsew signal input
rlabel metal2 s 35162 -800 35218 800 8 la_reset[11]
port 127 nsew signal input
rlabel metal2 s 32218 -800 32274 800 8 la_reset[1]
port 128 nsew signal input
rlabel metal2 s 32494 -800 32550 800 8 la_reset[2]
port 129 nsew signal input
rlabel metal2 s 32770 -800 32826 800 8 la_reset[3]
port 130 nsew signal input
rlabel metal2 s 33046 -800 33102 800 8 la_reset[4]
port 131 nsew signal input
rlabel metal2 s 33322 -800 33378 800 8 la_reset[5]
port 132 nsew signal input
rlabel metal2 s 33690 -800 33746 800 8 la_reset[6]
port 133 nsew signal input
rlabel metal2 s 33966 -800 34022 800 8 la_reset[7]
port 134 nsew signal input
rlabel metal2 s 34242 -800 34298 800 8 la_reset[8]
port 135 nsew signal input
rlabel metal2 s 34518 -800 34574 800 8 la_reset[9]
port 136 nsew signal input
rlabel metal2 s 31574 119200 31630 120800 6 m_irqs[0]
port 137 nsew signal input
rlabel metal2 s 33690 119200 33746 120800 6 m_irqs[10]
port 138 nsew signal input
rlabel metal2 s 33966 119200 34022 120800 6 m_irqs[11]
port 139 nsew signal input
rlabel metal2 s 31850 119200 31906 120800 6 m_irqs[1]
port 140 nsew signal input
rlabel metal2 s 32034 119200 32090 120800 6 m_irqs[2]
port 141 nsew signal input
rlabel metal2 s 32218 119200 32274 120800 6 m_irqs[3]
port 142 nsew signal input
rlabel metal2 s 32494 119200 32550 120800 6 m_irqs[4]
port 143 nsew signal input
rlabel metal2 s 32678 119200 32734 120800 6 m_irqs[5]
port 144 nsew signal input
rlabel metal2 s 32862 119200 32918 120800 6 m_irqs[6]
port 145 nsew signal input
rlabel metal2 s 33138 119200 33194 120800 6 m_irqs[7]
port 146 nsew signal input
rlabel metal2 s 33322 119200 33378 120800 6 m_irqs[8]
port 147 nsew signal input
rlabel metal2 s 33506 119200 33562 120800 6 m_irqs[9]
port 148 nsew signal input
rlabel metal2 s 34150 119200 34206 120800 6 m_la_reset[0]
port 149 nsew signal tristate
rlabel metal2 s 36266 119200 36322 120800 6 m_la_reset[10]
port 150 nsew signal tristate
rlabel metal2 s 36450 119200 36506 120800 6 m_la_reset[11]
port 151 nsew signal tristate
rlabel metal2 s 34334 119200 34390 120800 6 m_la_reset[1]
port 152 nsew signal tristate
rlabel metal2 s 34610 119200 34666 120800 6 m_la_reset[2]
port 153 nsew signal tristate
rlabel metal2 s 34794 119200 34850 120800 6 m_la_reset[3]
port 154 nsew signal tristate
rlabel metal2 s 34978 119200 35034 120800 6 m_la_reset[4]
port 155 nsew signal tristate
rlabel metal2 s 35254 119200 35310 120800 6 m_la_reset[5]
port 156 nsew signal tristate
rlabel metal2 s 35438 119200 35494 120800 6 m_la_reset[6]
port 157 nsew signal tristate
rlabel metal2 s 35622 119200 35678 120800 6 m_la_reset[7]
port 158 nsew signal tristate
rlabel metal2 s 35806 119200 35862 120800 6 m_la_reset[8]
port 159 nsew signal tristate
rlabel metal2 s 36082 119200 36138 120800 6 m_la_reset[9]
port 160 nsew signal tristate
rlabel metal2 s 35438 -800 35494 800 8 m_wb_clk_i
port 161 nsew signal tristate
rlabel metal3 s -800 106224 800 106344 4 m_wb_rst_i
port 162 nsew signal tristate
rlabel metal3 s 39200 110576 40800 110696 6 m_wbs_ack_o[0]
port 163 nsew signal input
rlabel metal2 s 38290 -800 38346 800 8 m_wbs_ack_o[10]
port 164 nsew signal input
rlabel metal3 s 39200 116560 40800 116680 6 m_wbs_ack_o[11]
port 165 nsew signal input
rlabel metal3 s 39200 111800 40800 111920 6 m_wbs_ack_o[1]
port 166 nsew signal input
rlabel metal2 s 35714 -800 35770 800 8 m_wbs_ack_o[2]
port 167 nsew signal input
rlabel metal2 s 37094 119200 37150 120800 6 m_wbs_ack_o[3]
port 168 nsew signal input
rlabel metal2 s 36542 -800 36598 800 8 m_wbs_ack_o[4]
port 169 nsew signal input
rlabel metal3 s 39200 114384 40800 114504 6 m_wbs_ack_o[5]
port 170 nsew signal input
rlabel metal2 s 37738 119200 37794 120800 6 m_wbs_ack_o[6]
port 171 nsew signal input
rlabel metal3 s 39200 115336 40800 115456 6 m_wbs_ack_o[7]
port 172 nsew signal input
rlabel metal3 s -800 111256 800 111376 4 m_wbs_ack_o[8]
port 173 nsew signal input
rlabel metal3 s -800 112888 800 113008 4 m_wbs_ack_o[9]
port 174 nsew signal input
rlabel metal3 s 39200 110984 40800 111104 6 m_wbs_adr_i[0]
port 175 nsew signal tristate
rlabel metal3 s -800 114520 800 114640 4 m_wbs_adr_i[10]
port 176 nsew signal tristate
rlabel metal3 s 39200 116968 40800 117088 6 m_wbs_adr_i[11]
port 177 nsew signal tristate
rlabel metal3 s 39200 112208 40800 112328 6 m_wbs_adr_i[1]
port 178 nsew signal tristate
rlabel metal2 s 35990 -800 36046 800 8 m_wbs_adr_i[2]
port 179 nsew signal tristate
rlabel metal3 s 39200 112752 40800 112872 6 m_wbs_adr_i[3]
port 180 nsew signal tristate
rlabel metal2 s 36910 -800 36966 800 8 m_wbs_adr_i[4]
port 181 nsew signal tristate
rlabel metal2 s 37186 -800 37242 800 8 m_wbs_adr_i[5]
port 182 nsew signal tristate
rlabel metal2 s 37922 119200 37978 120800 6 m_wbs_adr_i[6]
port 183 nsew signal tristate
rlabel metal3 s 39200 115744 40800 115864 6 m_wbs_adr_i[7]
port 184 nsew signal tristate
rlabel metal2 s 38198 119200 38254 120800 6 m_wbs_adr_i[8]
port 185 nsew signal tristate
rlabel metal3 s -800 113704 800 113824 4 m_wbs_adr_i[9]
port 186 nsew signal tristate
rlabel metal3 s -800 107040 800 107160 4 m_wbs_cs_i[0]
port 187 nsew signal tristate
rlabel metal3 s -800 115336 800 115456 4 m_wbs_cs_i[10]
port 188 nsew signal tristate
rlabel metal2 s 38658 -800 38714 800 8 m_wbs_cs_i[11]
port 189 nsew signal tristate
rlabel metal3 s -800 107856 800 107976 4 m_wbs_cs_i[1]
port 190 nsew signal tristate
rlabel metal3 s -800 108672 800 108792 4 m_wbs_cs_i[2]
port 191 nsew signal tristate
rlabel metal3 s 39200 113160 40800 113280 6 m_wbs_cs_i[3]
port 192 nsew signal tristate
rlabel metal3 s 39200 113976 40800 114096 6 m_wbs_cs_i[4]
port 193 nsew signal tristate
rlabel metal3 s -800 109488 800 109608 4 m_wbs_cs_i[5]
port 194 nsew signal tristate
rlabel metal3 s 39200 114792 40800 114912 6 m_wbs_cs_i[6]
port 195 nsew signal tristate
rlabel metal2 s 37738 -800 37794 800 8 m_wbs_cs_i[7]
port 196 nsew signal tristate
rlabel metal3 s -800 112072 800 112192 4 m_wbs_cs_i[8]
port 197 nsew signal tristate
rlabel metal2 s 38014 -800 38070 800 8 m_wbs_cs_i[9]
port 198 nsew signal tristate
rlabel metal3 s 39200 111392 40800 111512 6 m_wbs_dat_i[0]
port 199 nsew signal tristate
rlabel metal3 s 39200 116152 40800 116272 6 m_wbs_dat_i[10]
port 200 nsew signal tristate
rlabel metal3 s -800 116152 800 116272 4 m_wbs_dat_i[11]
port 201 nsew signal tristate
rlabel metal2 s 38934 -800 38990 800 8 m_wbs_dat_i[12]
port 202 nsew signal tristate
rlabel metal3 s -800 116968 800 117088 4 m_wbs_dat_i[13]
port 203 nsew signal tristate
rlabel metal2 s 38842 119200 38898 120800 6 m_wbs_dat_i[14]
port 204 nsew signal tristate
rlabel metal3 s -800 117784 800 117904 4 m_wbs_dat_i[15]
port 205 nsew signal tristate
rlabel metal2 s 39026 119200 39082 120800 6 m_wbs_dat_i[16]
port 206 nsew signal tristate
rlabel metal3 s 39200 117376 40800 117496 6 m_wbs_dat_i[17]
port 207 nsew signal tristate
rlabel metal2 s 39210 119200 39266 120800 6 m_wbs_dat_i[18]
port 208 nsew signal tristate
rlabel metal2 s 39486 119200 39542 120800 6 m_wbs_dat_i[19]
port 209 nsew signal tristate
rlabel metal2 s 36910 119200 36966 120800 6 m_wbs_dat_i[1]
port 210 nsew signal tristate
rlabel metal3 s -800 118600 800 118720 4 m_wbs_dat_i[20]
port 211 nsew signal tristate
rlabel metal2 s 39210 -800 39266 800 8 m_wbs_dat_i[21]
port 212 nsew signal tristate
rlabel metal3 s 39200 117920 40800 118040 6 m_wbs_dat_i[22]
port 213 nsew signal tristate
rlabel metal3 s 39200 118328 40800 118448 6 m_wbs_dat_i[23]
port 214 nsew signal tristate
rlabel metal2 s 39486 -800 39542 800 8 m_wbs_dat_i[24]
port 215 nsew signal tristate
rlabel metal2 s 39670 119200 39726 120800 6 m_wbs_dat_i[25]
port 216 nsew signal tristate
rlabel metal3 s 39200 118736 40800 118856 6 m_wbs_dat_i[26]
port 217 nsew signal tristate
rlabel metal3 s 39200 119144 40800 119264 6 m_wbs_dat_i[27]
port 218 nsew signal tristate
rlabel metal3 s 39200 119552 40800 119672 6 m_wbs_dat_i[28]
port 219 nsew signal tristate
rlabel metal2 s 39854 119200 39910 120800 6 m_wbs_dat_i[29]
port 220 nsew signal tristate
rlabel metal2 s 36266 -800 36322 800 8 m_wbs_dat_i[2]
port 221 nsew signal tristate
rlabel metal3 s -800 119416 800 119536 4 m_wbs_dat_i[30]
port 222 nsew signal tristate
rlabel metal2 s 39762 -800 39818 800 8 m_wbs_dat_i[31]
port 223 nsew signal tristate
rlabel metal3 s 39200 113568 40800 113688 6 m_wbs_dat_i[3]
port 224 nsew signal tristate
rlabel metal2 s 37370 119200 37426 120800 6 m_wbs_dat_i[4]
port 225 nsew signal tristate
rlabel metal2 s 37554 119200 37610 120800 6 m_wbs_dat_i[5]
port 226 nsew signal tristate
rlabel metal2 s 37462 -800 37518 800 8 m_wbs_dat_i[6]
port 227 nsew signal tristate
rlabel metal3 s -800 110440 800 110560 4 m_wbs_dat_i[7]
port 228 nsew signal tristate
rlabel metal2 s 38382 119200 38438 120800 6 m_wbs_dat_i[8]
port 229 nsew signal tristate
rlabel metal2 s 38566 119200 38622 120800 6 m_wbs_dat_i[9]
port 230 nsew signal tristate
rlabel metal3 s 39200 144 40800 264 6 m_wbs_dat_o_0[0]
port 231 nsew signal input
rlabel metal3 s 39200 4360 40800 4480 6 m_wbs_dat_o_0[10]
port 232 nsew signal input
rlabel metal3 s 39200 4768 40800 4888 6 m_wbs_dat_o_0[11]
port 233 nsew signal input
rlabel metal3 s 39200 5312 40800 5432 6 m_wbs_dat_o_0[12]
port 234 nsew signal input
rlabel metal3 s 39200 5720 40800 5840 6 m_wbs_dat_o_0[13]
port 235 nsew signal input
rlabel metal3 s 39200 6128 40800 6248 6 m_wbs_dat_o_0[14]
port 236 nsew signal input
rlabel metal3 s 39200 6536 40800 6656 6 m_wbs_dat_o_0[15]
port 237 nsew signal input
rlabel metal3 s 39200 6944 40800 7064 6 m_wbs_dat_o_0[16]
port 238 nsew signal input
rlabel metal3 s 39200 7352 40800 7472 6 m_wbs_dat_o_0[17]
port 239 nsew signal input
rlabel metal3 s 39200 7896 40800 8016 6 m_wbs_dat_o_0[18]
port 240 nsew signal input
rlabel metal3 s 39200 8304 40800 8424 6 m_wbs_dat_o_0[19]
port 241 nsew signal input
rlabel metal3 s 39200 552 40800 672 6 m_wbs_dat_o_0[1]
port 242 nsew signal input
rlabel metal3 s 39200 8712 40800 8832 6 m_wbs_dat_o_0[20]
port 243 nsew signal input
rlabel metal3 s 39200 9120 40800 9240 6 m_wbs_dat_o_0[21]
port 244 nsew signal input
rlabel metal3 s 39200 9528 40800 9648 6 m_wbs_dat_o_0[22]
port 245 nsew signal input
rlabel metal3 s 39200 9936 40800 10056 6 m_wbs_dat_o_0[23]
port 246 nsew signal input
rlabel metal3 s 39200 10480 40800 10600 6 m_wbs_dat_o_0[24]
port 247 nsew signal input
rlabel metal3 s 39200 10888 40800 11008 6 m_wbs_dat_o_0[25]
port 248 nsew signal input
rlabel metal3 s 39200 11296 40800 11416 6 m_wbs_dat_o_0[26]
port 249 nsew signal input
rlabel metal3 s 39200 11704 40800 11824 6 m_wbs_dat_o_0[27]
port 250 nsew signal input
rlabel metal3 s 39200 12112 40800 12232 6 m_wbs_dat_o_0[28]
port 251 nsew signal input
rlabel metal3 s 39200 12656 40800 12776 6 m_wbs_dat_o_0[29]
port 252 nsew signal input
rlabel metal3 s 39200 960 40800 1080 6 m_wbs_dat_o_0[2]
port 253 nsew signal input
rlabel metal3 s 39200 13064 40800 13184 6 m_wbs_dat_o_0[30]
port 254 nsew signal input
rlabel metal3 s 39200 13472 40800 13592 6 m_wbs_dat_o_0[31]
port 255 nsew signal input
rlabel metal3 s 39200 1368 40800 1488 6 m_wbs_dat_o_0[3]
port 256 nsew signal input
rlabel metal3 s 39200 1776 40800 1896 6 m_wbs_dat_o_0[4]
port 257 nsew signal input
rlabel metal3 s 39200 2184 40800 2304 6 m_wbs_dat_o_0[5]
port 258 nsew signal input
rlabel metal3 s 39200 2728 40800 2848 6 m_wbs_dat_o_0[6]
port 259 nsew signal input
rlabel metal3 s 39200 3136 40800 3256 6 m_wbs_dat_o_0[7]
port 260 nsew signal input
rlabel metal3 s 39200 3544 40800 3664 6 m_wbs_dat_o_0[8]
port 261 nsew signal input
rlabel metal3 s 39200 3952 40800 4072 6 m_wbs_dat_o_0[9]
port 262 nsew signal input
rlabel metal3 s 39200 14288 40800 14408 6 m_wbs_dat_o_10[0]
port 263 nsew signal input
rlabel metal3 s 39200 27208 40800 27328 6 m_wbs_dat_o_10[10]
port 264 nsew signal input
rlabel metal3 s 39200 28568 40800 28688 6 m_wbs_dat_o_10[11]
port 265 nsew signal input
rlabel metal3 s 39200 29792 40800 29912 6 m_wbs_dat_o_10[12]
port 266 nsew signal input
rlabel metal3 s 39200 31152 40800 31272 6 m_wbs_dat_o_10[13]
port 267 nsew signal input
rlabel metal3 s 39200 32376 40800 32496 6 m_wbs_dat_o_10[14]
port 268 nsew signal input
rlabel metal3 s 39200 33736 40800 33856 6 m_wbs_dat_o_10[15]
port 269 nsew signal input
rlabel metal3 s 39200 34960 40800 35080 6 m_wbs_dat_o_10[16]
port 270 nsew signal input
rlabel metal3 s 39200 36320 40800 36440 6 m_wbs_dat_o_10[17]
port 271 nsew signal input
rlabel metal3 s 39200 37680 40800 37800 6 m_wbs_dat_o_10[18]
port 272 nsew signal input
rlabel metal3 s 39200 38904 40800 39024 6 m_wbs_dat_o_10[19]
port 273 nsew signal input
rlabel metal3 s 39200 15648 40800 15768 6 m_wbs_dat_o_10[1]
port 274 nsew signal input
rlabel metal3 s 39200 40264 40800 40384 6 m_wbs_dat_o_10[20]
port 275 nsew signal input
rlabel metal3 s 39200 41488 40800 41608 6 m_wbs_dat_o_10[21]
port 276 nsew signal input
rlabel metal3 s 39200 42848 40800 42968 6 m_wbs_dat_o_10[22]
port 277 nsew signal input
rlabel metal3 s 39200 44072 40800 44192 6 m_wbs_dat_o_10[23]
port 278 nsew signal input
rlabel metal3 s 39200 45432 40800 45552 6 m_wbs_dat_o_10[24]
port 279 nsew signal input
rlabel metal3 s 39200 46656 40800 46776 6 m_wbs_dat_o_10[25]
port 280 nsew signal input
rlabel metal3 s 39200 48016 40800 48136 6 m_wbs_dat_o_10[26]
port 281 nsew signal input
rlabel metal3 s 39200 49240 40800 49360 6 m_wbs_dat_o_10[27]
port 282 nsew signal input
rlabel metal3 s 39200 50600 40800 50720 6 m_wbs_dat_o_10[28]
port 283 nsew signal input
rlabel metal3 s 39200 51824 40800 51944 6 m_wbs_dat_o_10[29]
port 284 nsew signal input
rlabel metal3 s 39200 16872 40800 16992 6 m_wbs_dat_o_10[2]
port 285 nsew signal input
rlabel metal3 s 39200 53184 40800 53304 6 m_wbs_dat_o_10[30]
port 286 nsew signal input
rlabel metal3 s 39200 54408 40800 54528 6 m_wbs_dat_o_10[31]
port 287 nsew signal input
rlabel metal3 s 39200 18232 40800 18352 6 m_wbs_dat_o_10[3]
port 288 nsew signal input
rlabel metal3 s 39200 19456 40800 19576 6 m_wbs_dat_o_10[4]
port 289 nsew signal input
rlabel metal3 s 39200 20816 40800 20936 6 m_wbs_dat_o_10[5]
port 290 nsew signal input
rlabel metal3 s 39200 22040 40800 22160 6 m_wbs_dat_o_10[6]
port 291 nsew signal input
rlabel metal3 s 39200 23400 40800 23520 6 m_wbs_dat_o_10[7]
port 292 nsew signal input
rlabel metal3 s 39200 24624 40800 24744 6 m_wbs_dat_o_10[8]
port 293 nsew signal input
rlabel metal3 s 39200 25984 40800 26104 6 m_wbs_dat_o_10[9]
port 294 nsew signal input
rlabel metal3 s 39200 14696 40800 14816 6 m_wbs_dat_o_11[0]
port 295 nsew signal input
rlabel metal3 s 39200 27752 40800 27872 6 m_wbs_dat_o_11[10]
port 296 nsew signal input
rlabel metal3 s 39200 28976 40800 29096 6 m_wbs_dat_o_11[11]
port 297 nsew signal input
rlabel metal3 s 39200 30336 40800 30456 6 m_wbs_dat_o_11[12]
port 298 nsew signal input
rlabel metal3 s 39200 31560 40800 31680 6 m_wbs_dat_o_11[13]
port 299 nsew signal input
rlabel metal3 s 39200 32920 40800 33040 6 m_wbs_dat_o_11[14]
port 300 nsew signal input
rlabel metal3 s 39200 34144 40800 34264 6 m_wbs_dat_o_11[15]
port 301 nsew signal input
rlabel metal3 s 39200 35504 40800 35624 6 m_wbs_dat_o_11[16]
port 302 nsew signal input
rlabel metal3 s 39200 36728 40800 36848 6 m_wbs_dat_o_11[17]
port 303 nsew signal input
rlabel metal3 s 39200 38088 40800 38208 6 m_wbs_dat_o_11[18]
port 304 nsew signal input
rlabel metal3 s 39200 39312 40800 39432 6 m_wbs_dat_o_11[19]
port 305 nsew signal input
rlabel metal3 s 39200 16056 40800 16176 6 m_wbs_dat_o_11[1]
port 306 nsew signal input
rlabel metal3 s 39200 40672 40800 40792 6 m_wbs_dat_o_11[20]
port 307 nsew signal input
rlabel metal3 s 39200 41896 40800 42016 6 m_wbs_dat_o_11[21]
port 308 nsew signal input
rlabel metal3 s 39200 43256 40800 43376 6 m_wbs_dat_o_11[22]
port 309 nsew signal input
rlabel metal3 s 39200 44480 40800 44600 6 m_wbs_dat_o_11[23]
port 310 nsew signal input
rlabel metal3 s 39200 45840 40800 45960 6 m_wbs_dat_o_11[24]
port 311 nsew signal input
rlabel metal3 s 39200 47064 40800 47184 6 m_wbs_dat_o_11[25]
port 312 nsew signal input
rlabel metal3 s 39200 48424 40800 48544 6 m_wbs_dat_o_11[26]
port 313 nsew signal input
rlabel metal3 s 39200 49648 40800 49768 6 m_wbs_dat_o_11[27]
port 314 nsew signal input
rlabel metal3 s 39200 51008 40800 51128 6 m_wbs_dat_o_11[28]
port 315 nsew signal input
rlabel metal3 s 39200 52232 40800 52352 6 m_wbs_dat_o_11[29]
port 316 nsew signal input
rlabel metal3 s 39200 17280 40800 17400 6 m_wbs_dat_o_11[2]
port 317 nsew signal input
rlabel metal3 s 39200 53592 40800 53712 6 m_wbs_dat_o_11[30]
port 318 nsew signal input
rlabel metal3 s 39200 54816 40800 54936 6 m_wbs_dat_o_11[31]
port 319 nsew signal input
rlabel metal3 s 39200 18640 40800 18760 6 m_wbs_dat_o_11[3]
port 320 nsew signal input
rlabel metal3 s 39200 19864 40800 19984 6 m_wbs_dat_o_11[4]
port 321 nsew signal input
rlabel metal3 s 39200 21224 40800 21344 6 m_wbs_dat_o_11[5]
port 322 nsew signal input
rlabel metal3 s 39200 22448 40800 22568 6 m_wbs_dat_o_11[6]
port 323 nsew signal input
rlabel metal3 s 39200 23808 40800 23928 6 m_wbs_dat_o_11[7]
port 324 nsew signal input
rlabel metal3 s 39200 25168 40800 25288 6 m_wbs_dat_o_11[8]
port 325 nsew signal input
rlabel metal3 s 39200 26392 40800 26512 6 m_wbs_dat_o_11[9]
port 326 nsew signal input
rlabel metal3 s 39200 13880 40800 14000 6 m_wbs_dat_o_1[0]
port 327 nsew signal input
rlabel metal3 s 39200 26800 40800 26920 6 m_wbs_dat_o_1[10]
port 328 nsew signal input
rlabel metal3 s 39200 28160 40800 28280 6 m_wbs_dat_o_1[11]
port 329 nsew signal input
rlabel metal3 s 39200 29384 40800 29504 6 m_wbs_dat_o_1[12]
port 330 nsew signal input
rlabel metal3 s 39200 30744 40800 30864 6 m_wbs_dat_o_1[13]
port 331 nsew signal input
rlabel metal3 s 39200 31968 40800 32088 6 m_wbs_dat_o_1[14]
port 332 nsew signal input
rlabel metal3 s 39200 33328 40800 33448 6 m_wbs_dat_o_1[15]
port 333 nsew signal input
rlabel metal3 s 39200 34552 40800 34672 6 m_wbs_dat_o_1[16]
port 334 nsew signal input
rlabel metal3 s 39200 35912 40800 36032 6 m_wbs_dat_o_1[17]
port 335 nsew signal input
rlabel metal3 s 39200 37136 40800 37256 6 m_wbs_dat_o_1[18]
port 336 nsew signal input
rlabel metal3 s 39200 38496 40800 38616 6 m_wbs_dat_o_1[19]
port 337 nsew signal input
rlabel metal3 s 39200 15240 40800 15360 6 m_wbs_dat_o_1[1]
port 338 nsew signal input
rlabel metal3 s 39200 39720 40800 39840 6 m_wbs_dat_o_1[20]
port 339 nsew signal input
rlabel metal3 s 39200 41080 40800 41200 6 m_wbs_dat_o_1[21]
port 340 nsew signal input
rlabel metal3 s 39200 42304 40800 42424 6 m_wbs_dat_o_1[22]
port 341 nsew signal input
rlabel metal3 s 39200 43664 40800 43784 6 m_wbs_dat_o_1[23]
port 342 nsew signal input
rlabel metal3 s 39200 44888 40800 45008 6 m_wbs_dat_o_1[24]
port 343 nsew signal input
rlabel metal3 s 39200 46248 40800 46368 6 m_wbs_dat_o_1[25]
port 344 nsew signal input
rlabel metal3 s 39200 47472 40800 47592 6 m_wbs_dat_o_1[26]
port 345 nsew signal input
rlabel metal3 s 39200 48832 40800 48952 6 m_wbs_dat_o_1[27]
port 346 nsew signal input
rlabel metal3 s 39200 50192 40800 50312 6 m_wbs_dat_o_1[28]
port 347 nsew signal input
rlabel metal3 s 39200 51416 40800 51536 6 m_wbs_dat_o_1[29]
port 348 nsew signal input
rlabel metal3 s 39200 16464 40800 16584 6 m_wbs_dat_o_1[2]
port 349 nsew signal input
rlabel metal3 s 39200 52776 40800 52896 6 m_wbs_dat_o_1[30]
port 350 nsew signal input
rlabel metal3 s 39200 54000 40800 54120 6 m_wbs_dat_o_1[31]
port 351 nsew signal input
rlabel metal3 s 39200 17824 40800 17944 6 m_wbs_dat_o_1[3]
port 352 nsew signal input
rlabel metal3 s 39200 19048 40800 19168 6 m_wbs_dat_o_1[4]
port 353 nsew signal input
rlabel metal3 s 39200 20408 40800 20528 6 m_wbs_dat_o_1[5]
port 354 nsew signal input
rlabel metal3 s 39200 21632 40800 21752 6 m_wbs_dat_o_1[6]
port 355 nsew signal input
rlabel metal3 s 39200 22992 40800 23112 6 m_wbs_dat_o_1[7]
port 356 nsew signal input
rlabel metal3 s 39200 24216 40800 24336 6 m_wbs_dat_o_1[8]
port 357 nsew signal input
rlabel metal3 s 39200 25576 40800 25696 6 m_wbs_dat_o_1[9]
port 358 nsew signal input
rlabel metal3 s 39200 55360 40800 55480 6 m_wbs_dat_o_2[0]
port 359 nsew signal input
rlabel metal3 s 39200 59576 40800 59696 6 m_wbs_dat_o_2[10]
port 360 nsew signal input
rlabel metal3 s 39200 60120 40800 60240 6 m_wbs_dat_o_2[11]
port 361 nsew signal input
rlabel metal3 s 39200 60528 40800 60648 6 m_wbs_dat_o_2[12]
port 362 nsew signal input
rlabel metal3 s 39200 60936 40800 61056 6 m_wbs_dat_o_2[13]
port 363 nsew signal input
rlabel metal3 s 39200 61344 40800 61464 6 m_wbs_dat_o_2[14]
port 364 nsew signal input
rlabel metal3 s 39200 61752 40800 61872 6 m_wbs_dat_o_2[15]
port 365 nsew signal input
rlabel metal3 s 39200 62160 40800 62280 6 m_wbs_dat_o_2[16]
port 366 nsew signal input
rlabel metal3 s 39200 62704 40800 62824 6 m_wbs_dat_o_2[17]
port 367 nsew signal input
rlabel metal3 s 39200 63112 40800 63232 6 m_wbs_dat_o_2[18]
port 368 nsew signal input
rlabel metal3 s 39200 63520 40800 63640 6 m_wbs_dat_o_2[19]
port 369 nsew signal input
rlabel metal3 s 39200 55768 40800 55888 6 m_wbs_dat_o_2[1]
port 370 nsew signal input
rlabel metal3 s 39200 63928 40800 64048 6 m_wbs_dat_o_2[20]
port 371 nsew signal input
rlabel metal3 s 39200 64336 40800 64456 6 m_wbs_dat_o_2[21]
port 372 nsew signal input
rlabel metal3 s 39200 64744 40800 64864 6 m_wbs_dat_o_2[22]
port 373 nsew signal input
rlabel metal3 s 39200 65288 40800 65408 6 m_wbs_dat_o_2[23]
port 374 nsew signal input
rlabel metal3 s 39200 65696 40800 65816 6 m_wbs_dat_o_2[24]
port 375 nsew signal input
rlabel metal3 s 39200 66104 40800 66224 6 m_wbs_dat_o_2[25]
port 376 nsew signal input
rlabel metal3 s 39200 66512 40800 66632 6 m_wbs_dat_o_2[26]
port 377 nsew signal input
rlabel metal3 s 39200 66920 40800 67040 6 m_wbs_dat_o_2[27]
port 378 nsew signal input
rlabel metal3 s 39200 67328 40800 67448 6 m_wbs_dat_o_2[28]
port 379 nsew signal input
rlabel metal3 s 39200 67872 40800 67992 6 m_wbs_dat_o_2[29]
port 380 nsew signal input
rlabel metal3 s 39200 56176 40800 56296 6 m_wbs_dat_o_2[2]
port 381 nsew signal input
rlabel metal3 s 39200 68280 40800 68400 6 m_wbs_dat_o_2[30]
port 382 nsew signal input
rlabel metal3 s 39200 68688 40800 68808 6 m_wbs_dat_o_2[31]
port 383 nsew signal input
rlabel metal3 s 39200 56584 40800 56704 6 m_wbs_dat_o_2[3]
port 384 nsew signal input
rlabel metal3 s 39200 56992 40800 57112 6 m_wbs_dat_o_2[4]
port 385 nsew signal input
rlabel metal3 s 39200 57400 40800 57520 6 m_wbs_dat_o_2[5]
port 386 nsew signal input
rlabel metal3 s 39200 57944 40800 58064 6 m_wbs_dat_o_2[6]
port 387 nsew signal input
rlabel metal3 s 39200 58352 40800 58472 6 m_wbs_dat_o_2[7]
port 388 nsew signal input
rlabel metal3 s 39200 58760 40800 58880 6 m_wbs_dat_o_2[8]
port 389 nsew signal input
rlabel metal3 s 39200 59168 40800 59288 6 m_wbs_dat_o_2[9]
port 390 nsew signal input
rlabel metal3 s 39200 69096 40800 69216 6 m_wbs_dat_o_3[0]
port 391 nsew signal input
rlabel metal3 s 39200 73448 40800 73568 6 m_wbs_dat_o_3[10]
port 392 nsew signal input
rlabel metal3 s 39200 73856 40800 73976 6 m_wbs_dat_o_3[11]
port 393 nsew signal input
rlabel metal3 s 39200 74264 40800 74384 6 m_wbs_dat_o_3[12]
port 394 nsew signal input
rlabel metal3 s 39200 74672 40800 74792 6 m_wbs_dat_o_3[13]
port 395 nsew signal input
rlabel metal3 s 39200 75216 40800 75336 6 m_wbs_dat_o_3[14]
port 396 nsew signal input
rlabel metal3 s 39200 75624 40800 75744 6 m_wbs_dat_o_3[15]
port 397 nsew signal input
rlabel metal3 s 39200 76032 40800 76152 6 m_wbs_dat_o_3[16]
port 398 nsew signal input
rlabel metal3 s 39200 76440 40800 76560 6 m_wbs_dat_o_3[17]
port 399 nsew signal input
rlabel metal3 s 39200 76848 40800 76968 6 m_wbs_dat_o_3[18]
port 400 nsew signal input
rlabel metal3 s 39200 77256 40800 77376 6 m_wbs_dat_o_3[19]
port 401 nsew signal input
rlabel metal3 s 39200 69504 40800 69624 6 m_wbs_dat_o_3[1]
port 402 nsew signal input
rlabel metal3 s 39200 77800 40800 77920 6 m_wbs_dat_o_3[20]
port 403 nsew signal input
rlabel metal3 s 39200 78208 40800 78328 6 m_wbs_dat_o_3[21]
port 404 nsew signal input
rlabel metal3 s 39200 78616 40800 78736 6 m_wbs_dat_o_3[22]
port 405 nsew signal input
rlabel metal3 s 39200 79024 40800 79144 6 m_wbs_dat_o_3[23]
port 406 nsew signal input
rlabel metal3 s 39200 79432 40800 79552 6 m_wbs_dat_o_3[24]
port 407 nsew signal input
rlabel metal3 s 39200 79840 40800 79960 6 m_wbs_dat_o_3[25]
port 408 nsew signal input
rlabel metal3 s 39200 80384 40800 80504 6 m_wbs_dat_o_3[26]
port 409 nsew signal input
rlabel metal3 s 39200 80792 40800 80912 6 m_wbs_dat_o_3[27]
port 410 nsew signal input
rlabel metal3 s 39200 81200 40800 81320 6 m_wbs_dat_o_3[28]
port 411 nsew signal input
rlabel metal3 s 39200 81608 40800 81728 6 m_wbs_dat_o_3[29]
port 412 nsew signal input
rlabel metal3 s 39200 69912 40800 70032 6 m_wbs_dat_o_3[2]
port 413 nsew signal input
rlabel metal3 s 39200 82016 40800 82136 6 m_wbs_dat_o_3[30]
port 414 nsew signal input
rlabel metal3 s 39200 82424 40800 82544 6 m_wbs_dat_o_3[31]
port 415 nsew signal input
rlabel metal3 s 39200 70456 40800 70576 6 m_wbs_dat_o_3[3]
port 416 nsew signal input
rlabel metal3 s 39200 70864 40800 70984 6 m_wbs_dat_o_3[4]
port 417 nsew signal input
rlabel metal3 s 39200 71272 40800 71392 6 m_wbs_dat_o_3[5]
port 418 nsew signal input
rlabel metal3 s 39200 71680 40800 71800 6 m_wbs_dat_o_3[6]
port 419 nsew signal input
rlabel metal3 s 39200 72088 40800 72208 6 m_wbs_dat_o_3[7]
port 420 nsew signal input
rlabel metal3 s 39200 72632 40800 72752 6 m_wbs_dat_o_3[8]
port 421 nsew signal input
rlabel metal3 s 39200 73040 40800 73160 6 m_wbs_dat_o_3[9]
port 422 nsew signal input
rlabel metal3 s 39200 82968 40800 83088 6 m_wbs_dat_o_4[0]
port 423 nsew signal input
rlabel metal3 s 39200 87184 40800 87304 6 m_wbs_dat_o_4[10]
port 424 nsew signal input
rlabel metal3 s 39200 87728 40800 87848 6 m_wbs_dat_o_4[11]
port 425 nsew signal input
rlabel metal3 s 39200 88136 40800 88256 6 m_wbs_dat_o_4[12]
port 426 nsew signal input
rlabel metal3 s 39200 88544 40800 88664 6 m_wbs_dat_o_4[13]
port 427 nsew signal input
rlabel metal3 s 39200 88952 40800 89072 6 m_wbs_dat_o_4[14]
port 428 nsew signal input
rlabel metal3 s 39200 89360 40800 89480 6 m_wbs_dat_o_4[15]
port 429 nsew signal input
rlabel metal3 s 39200 89768 40800 89888 6 m_wbs_dat_o_4[16]
port 430 nsew signal input
rlabel metal3 s 39200 90312 40800 90432 6 m_wbs_dat_o_4[17]
port 431 nsew signal input
rlabel metal3 s 39200 90720 40800 90840 6 m_wbs_dat_o_4[18]
port 432 nsew signal input
rlabel metal3 s 39200 91128 40800 91248 6 m_wbs_dat_o_4[19]
port 433 nsew signal input
rlabel metal3 s 39200 83376 40800 83496 6 m_wbs_dat_o_4[1]
port 434 nsew signal input
rlabel metal3 s 39200 91536 40800 91656 6 m_wbs_dat_o_4[20]
port 435 nsew signal input
rlabel metal3 s 39200 91944 40800 92064 6 m_wbs_dat_o_4[21]
port 436 nsew signal input
rlabel metal3 s 39200 92352 40800 92472 6 m_wbs_dat_o_4[22]
port 437 nsew signal input
rlabel metal3 s 39200 92896 40800 93016 6 m_wbs_dat_o_4[23]
port 438 nsew signal input
rlabel metal3 s 39200 93304 40800 93424 6 m_wbs_dat_o_4[24]
port 439 nsew signal input
rlabel metal3 s 39200 93712 40800 93832 6 m_wbs_dat_o_4[25]
port 440 nsew signal input
rlabel metal3 s 39200 94120 40800 94240 6 m_wbs_dat_o_4[26]
port 441 nsew signal input
rlabel metal3 s 39200 94528 40800 94648 6 m_wbs_dat_o_4[27]
port 442 nsew signal input
rlabel metal3 s 39200 94936 40800 95056 6 m_wbs_dat_o_4[28]
port 443 nsew signal input
rlabel metal3 s 39200 95480 40800 95600 6 m_wbs_dat_o_4[29]
port 444 nsew signal input
rlabel metal3 s 39200 83784 40800 83904 6 m_wbs_dat_o_4[2]
port 445 nsew signal input
rlabel metal3 s 39200 95888 40800 96008 6 m_wbs_dat_o_4[30]
port 446 nsew signal input
rlabel metal3 s 39200 96296 40800 96416 6 m_wbs_dat_o_4[31]
port 447 nsew signal input
rlabel metal3 s 39200 84192 40800 84312 6 m_wbs_dat_o_4[3]
port 448 nsew signal input
rlabel metal3 s 39200 84600 40800 84720 6 m_wbs_dat_o_4[4]
port 449 nsew signal input
rlabel metal3 s 39200 85144 40800 85264 6 m_wbs_dat_o_4[5]
port 450 nsew signal input
rlabel metal3 s 39200 85552 40800 85672 6 m_wbs_dat_o_4[6]
port 451 nsew signal input
rlabel metal3 s 39200 85960 40800 86080 6 m_wbs_dat_o_4[7]
port 452 nsew signal input
rlabel metal3 s 39200 86368 40800 86488 6 m_wbs_dat_o_4[8]
port 453 nsew signal input
rlabel metal3 s 39200 86776 40800 86896 6 m_wbs_dat_o_4[9]
port 454 nsew signal input
rlabel metal3 s 39200 96704 40800 96824 6 m_wbs_dat_o_5[0]
port 455 nsew signal input
rlabel metal3 s 39200 101056 40800 101176 6 m_wbs_dat_o_5[10]
port 456 nsew signal input
rlabel metal3 s 39200 101464 40800 101584 6 m_wbs_dat_o_5[11]
port 457 nsew signal input
rlabel metal3 s 39200 101872 40800 101992 6 m_wbs_dat_o_5[12]
port 458 nsew signal input
rlabel metal3 s 39200 102280 40800 102400 6 m_wbs_dat_o_5[13]
port 459 nsew signal input
rlabel metal3 s 39200 102824 40800 102944 6 m_wbs_dat_o_5[14]
port 460 nsew signal input
rlabel metal3 s 39200 103232 40800 103352 6 m_wbs_dat_o_5[15]
port 461 nsew signal input
rlabel metal3 s 39200 103640 40800 103760 6 m_wbs_dat_o_5[16]
port 462 nsew signal input
rlabel metal3 s 39200 104048 40800 104168 6 m_wbs_dat_o_5[17]
port 463 nsew signal input
rlabel metal3 s 39200 104456 40800 104576 6 m_wbs_dat_o_5[18]
port 464 nsew signal input
rlabel metal3 s 39200 104864 40800 104984 6 m_wbs_dat_o_5[19]
port 465 nsew signal input
rlabel metal3 s 39200 97112 40800 97232 6 m_wbs_dat_o_5[1]
port 466 nsew signal input
rlabel metal3 s 39200 105408 40800 105528 6 m_wbs_dat_o_5[20]
port 467 nsew signal input
rlabel metal3 s 39200 105816 40800 105936 6 m_wbs_dat_o_5[21]
port 468 nsew signal input
rlabel metal3 s 39200 106224 40800 106344 6 m_wbs_dat_o_5[22]
port 469 nsew signal input
rlabel metal3 s 39200 106632 40800 106752 6 m_wbs_dat_o_5[23]
port 470 nsew signal input
rlabel metal3 s 39200 107040 40800 107160 6 m_wbs_dat_o_5[24]
port 471 nsew signal input
rlabel metal3 s 39200 107448 40800 107568 6 m_wbs_dat_o_5[25]
port 472 nsew signal input
rlabel metal3 s 39200 107992 40800 108112 6 m_wbs_dat_o_5[26]
port 473 nsew signal input
rlabel metal3 s 39200 108400 40800 108520 6 m_wbs_dat_o_5[27]
port 474 nsew signal input
rlabel metal3 s 39200 108808 40800 108928 6 m_wbs_dat_o_5[28]
port 475 nsew signal input
rlabel metal3 s 39200 109216 40800 109336 6 m_wbs_dat_o_5[29]
port 476 nsew signal input
rlabel metal3 s 39200 97656 40800 97776 6 m_wbs_dat_o_5[2]
port 477 nsew signal input
rlabel metal3 s 39200 109624 40800 109744 6 m_wbs_dat_o_5[30]
port 478 nsew signal input
rlabel metal3 s 39200 110168 40800 110288 6 m_wbs_dat_o_5[31]
port 479 nsew signal input
rlabel metal3 s 39200 98064 40800 98184 6 m_wbs_dat_o_5[3]
port 480 nsew signal input
rlabel metal3 s 39200 98472 40800 98592 6 m_wbs_dat_o_5[4]
port 481 nsew signal input
rlabel metal3 s 39200 98880 40800 99000 6 m_wbs_dat_o_5[5]
port 482 nsew signal input
rlabel metal3 s 39200 99288 40800 99408 6 m_wbs_dat_o_5[6]
port 483 nsew signal input
rlabel metal3 s 39200 99696 40800 99816 6 m_wbs_dat_o_5[7]
port 484 nsew signal input
rlabel metal3 s 39200 100240 40800 100360 6 m_wbs_dat_o_5[8]
port 485 nsew signal input
rlabel metal3 s 39200 100648 40800 100768 6 m_wbs_dat_o_5[9]
port 486 nsew signal input
rlabel metal3 s -800 416 800 536 4 m_wbs_dat_o_6[0]
port 487 nsew signal input
rlabel metal3 s -800 8576 800 8696 4 m_wbs_dat_o_6[10]
port 488 nsew signal input
rlabel metal3 s -800 9392 800 9512 4 m_wbs_dat_o_6[11]
port 489 nsew signal input
rlabel metal3 s -800 10208 800 10328 4 m_wbs_dat_o_6[12]
port 490 nsew signal input
rlabel metal3 s -800 11160 800 11280 4 m_wbs_dat_o_6[13]
port 491 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 m_wbs_dat_o_6[14]
port 492 nsew signal input
rlabel metal3 s -800 12792 800 12912 4 m_wbs_dat_o_6[15]
port 493 nsew signal input
rlabel metal3 s -800 13608 800 13728 4 m_wbs_dat_o_6[16]
port 494 nsew signal input
rlabel metal3 s -800 14424 800 14544 4 m_wbs_dat_o_6[17]
port 495 nsew signal input
rlabel metal3 s -800 15240 800 15360 4 m_wbs_dat_o_6[18]
port 496 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 m_wbs_dat_o_6[19]
port 497 nsew signal input
rlabel metal3 s -800 1232 800 1352 4 m_wbs_dat_o_6[1]
port 498 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 m_wbs_dat_o_6[20]
port 499 nsew signal input
rlabel metal3 s -800 17688 800 17808 4 m_wbs_dat_o_6[21]
port 500 nsew signal input
rlabel metal3 s -800 18504 800 18624 4 m_wbs_dat_o_6[22]
port 501 nsew signal input
rlabel metal3 s -800 19320 800 19440 4 m_wbs_dat_o_6[23]
port 502 nsew signal input
rlabel metal3 s -800 20136 800 20256 4 m_wbs_dat_o_6[24]
port 503 nsew signal input
rlabel metal3 s -800 21088 800 21208 4 m_wbs_dat_o_6[25]
port 504 nsew signal input
rlabel metal3 s -800 21904 800 22024 4 m_wbs_dat_o_6[26]
port 505 nsew signal input
rlabel metal3 s -800 22720 800 22840 4 m_wbs_dat_o_6[27]
port 506 nsew signal input
rlabel metal3 s -800 23536 800 23656 4 m_wbs_dat_o_6[28]
port 507 nsew signal input
rlabel metal3 s -800 24352 800 24472 4 m_wbs_dat_o_6[29]
port 508 nsew signal input
rlabel metal3 s -800 2048 800 2168 4 m_wbs_dat_o_6[2]
port 509 nsew signal input
rlabel metal3 s -800 25168 800 25288 4 m_wbs_dat_o_6[30]
port 510 nsew signal input
rlabel metal3 s -800 25984 800 26104 4 m_wbs_dat_o_6[31]
port 511 nsew signal input
rlabel metal3 s -800 2864 800 2984 4 m_wbs_dat_o_6[3]
port 512 nsew signal input
rlabel metal3 s -800 3680 800 3800 4 m_wbs_dat_o_6[4]
port 513 nsew signal input
rlabel metal3 s -800 4496 800 4616 4 m_wbs_dat_o_6[5]
port 514 nsew signal input
rlabel metal3 s -800 5312 800 5432 4 m_wbs_dat_o_6[6]
port 515 nsew signal input
rlabel metal3 s -800 6128 800 6248 4 m_wbs_dat_o_6[7]
port 516 nsew signal input
rlabel metal3 s -800 6944 800 7064 4 m_wbs_dat_o_6[8]
port 517 nsew signal input
rlabel metal3 s -800 7760 800 7880 4 m_wbs_dat_o_6[9]
port 518 nsew signal input
rlabel metal3 s -800 26800 800 26920 4 m_wbs_dat_o_7[0]
port 519 nsew signal input
rlabel metal3 s -800 35096 800 35216 4 m_wbs_dat_o_7[10]
port 520 nsew signal input
rlabel metal3 s -800 35912 800 36032 4 m_wbs_dat_o_7[11]
port 521 nsew signal input
rlabel metal3 s -800 36728 800 36848 4 m_wbs_dat_o_7[12]
port 522 nsew signal input
rlabel metal3 s -800 37544 800 37664 4 m_wbs_dat_o_7[13]
port 523 nsew signal input
rlabel metal3 s -800 38360 800 38480 4 m_wbs_dat_o_7[14]
port 524 nsew signal input
rlabel metal3 s -800 39176 800 39296 4 m_wbs_dat_o_7[15]
port 525 nsew signal input
rlabel metal3 s -800 39992 800 40112 4 m_wbs_dat_o_7[16]
port 526 nsew signal input
rlabel metal3 s -800 40944 800 41064 4 m_wbs_dat_o_7[17]
port 527 nsew signal input
rlabel metal3 s -800 41760 800 41880 4 m_wbs_dat_o_7[18]
port 528 nsew signal input
rlabel metal3 s -800 42576 800 42696 4 m_wbs_dat_o_7[19]
port 529 nsew signal input
rlabel metal3 s -800 27616 800 27736 4 m_wbs_dat_o_7[1]
port 530 nsew signal input
rlabel metal3 s -800 43392 800 43512 4 m_wbs_dat_o_7[20]
port 531 nsew signal input
rlabel metal3 s -800 44208 800 44328 4 m_wbs_dat_o_7[21]
port 532 nsew signal input
rlabel metal3 s -800 45024 800 45144 4 m_wbs_dat_o_7[22]
port 533 nsew signal input
rlabel metal3 s -800 45840 800 45960 4 m_wbs_dat_o_7[23]
port 534 nsew signal input
rlabel metal3 s -800 46656 800 46776 4 m_wbs_dat_o_7[24]
port 535 nsew signal input
rlabel metal3 s -800 47472 800 47592 4 m_wbs_dat_o_7[25]
port 536 nsew signal input
rlabel metal3 s -800 48288 800 48408 4 m_wbs_dat_o_7[26]
port 537 nsew signal input
rlabel metal3 s -800 49104 800 49224 4 m_wbs_dat_o_7[27]
port 538 nsew signal input
rlabel metal3 s -800 49920 800 50040 4 m_wbs_dat_o_7[28]
port 539 nsew signal input
rlabel metal3 s -800 50872 800 50992 4 m_wbs_dat_o_7[29]
port 540 nsew signal input
rlabel metal3 s -800 28432 800 28552 4 m_wbs_dat_o_7[2]
port 541 nsew signal input
rlabel metal3 s -800 51688 800 51808 4 m_wbs_dat_o_7[30]
port 542 nsew signal input
rlabel metal3 s -800 52504 800 52624 4 m_wbs_dat_o_7[31]
port 543 nsew signal input
rlabel metal3 s -800 29248 800 29368 4 m_wbs_dat_o_7[3]
port 544 nsew signal input
rlabel metal3 s -800 30064 800 30184 4 m_wbs_dat_o_7[4]
port 545 nsew signal input
rlabel metal3 s -800 31016 800 31136 4 m_wbs_dat_o_7[5]
port 546 nsew signal input
rlabel metal3 s -800 31832 800 31952 4 m_wbs_dat_o_7[6]
port 547 nsew signal input
rlabel metal3 s -800 32648 800 32768 4 m_wbs_dat_o_7[7]
port 548 nsew signal input
rlabel metal3 s -800 33464 800 33584 4 m_wbs_dat_o_7[8]
port 549 nsew signal input
rlabel metal3 s -800 34280 800 34400 4 m_wbs_dat_o_7[9]
port 550 nsew signal input
rlabel metal3 s -800 53320 800 53440 4 m_wbs_dat_o_8[0]
port 551 nsew signal input
rlabel metal3 s -800 61616 800 61736 4 m_wbs_dat_o_8[10]
port 552 nsew signal input
rlabel metal3 s -800 62432 800 62552 4 m_wbs_dat_o_8[11]
port 553 nsew signal input
rlabel metal3 s -800 63248 800 63368 4 m_wbs_dat_o_8[12]
port 554 nsew signal input
rlabel metal3 s -800 64064 800 64184 4 m_wbs_dat_o_8[13]
port 555 nsew signal input
rlabel metal3 s -800 64880 800 65000 4 m_wbs_dat_o_8[14]
port 556 nsew signal input
rlabel metal3 s -800 65696 800 65816 4 m_wbs_dat_o_8[15]
port 557 nsew signal input
rlabel metal3 s -800 66512 800 66632 4 m_wbs_dat_o_8[16]
port 558 nsew signal input
rlabel metal3 s -800 67328 800 67448 4 m_wbs_dat_o_8[17]
port 559 nsew signal input
rlabel metal3 s -800 68144 800 68264 4 m_wbs_dat_o_8[18]
port 560 nsew signal input
rlabel metal3 s -800 68960 800 69080 4 m_wbs_dat_o_8[19]
port 561 nsew signal input
rlabel metal3 s -800 54136 800 54256 4 m_wbs_dat_o_8[1]
port 562 nsew signal input
rlabel metal3 s -800 69776 800 69896 4 m_wbs_dat_o_8[20]
port 563 nsew signal input
rlabel metal3 s -800 70728 800 70848 4 m_wbs_dat_o_8[21]
port 564 nsew signal input
rlabel metal3 s -800 71544 800 71664 4 m_wbs_dat_o_8[22]
port 565 nsew signal input
rlabel metal3 s -800 72360 800 72480 4 m_wbs_dat_o_8[23]
port 566 nsew signal input
rlabel metal3 s -800 73176 800 73296 4 m_wbs_dat_o_8[24]
port 567 nsew signal input
rlabel metal3 s -800 73992 800 74112 4 m_wbs_dat_o_8[25]
port 568 nsew signal input
rlabel metal3 s -800 74808 800 74928 4 m_wbs_dat_o_8[26]
port 569 nsew signal input
rlabel metal3 s -800 75624 800 75744 4 m_wbs_dat_o_8[27]
port 570 nsew signal input
rlabel metal3 s -800 76440 800 76560 4 m_wbs_dat_o_8[28]
port 571 nsew signal input
rlabel metal3 s -800 77256 800 77376 4 m_wbs_dat_o_8[29]
port 572 nsew signal input
rlabel metal3 s -800 54952 800 55072 4 m_wbs_dat_o_8[2]
port 573 nsew signal input
rlabel metal3 s -800 78072 800 78192 4 m_wbs_dat_o_8[30]
port 574 nsew signal input
rlabel metal3 s -800 78888 800 79008 4 m_wbs_dat_o_8[31]
port 575 nsew signal input
rlabel metal3 s -800 55768 800 55888 4 m_wbs_dat_o_8[3]
port 576 nsew signal input
rlabel metal3 s -800 56584 800 56704 4 m_wbs_dat_o_8[4]
port 577 nsew signal input
rlabel metal3 s -800 57400 800 57520 4 m_wbs_dat_o_8[5]
port 578 nsew signal input
rlabel metal3 s -800 58216 800 58336 4 m_wbs_dat_o_8[6]
port 579 nsew signal input
rlabel metal3 s -800 59032 800 59152 4 m_wbs_dat_o_8[7]
port 580 nsew signal input
rlabel metal3 s -800 59848 800 59968 4 m_wbs_dat_o_8[8]
port 581 nsew signal input
rlabel metal3 s -800 60800 800 60920 4 m_wbs_dat_o_8[9]
port 582 nsew signal input
rlabel metal3 s -800 79704 800 79824 4 m_wbs_dat_o_9[0]
port 583 nsew signal input
rlabel metal3 s -800 88000 800 88120 4 m_wbs_dat_o_9[10]
port 584 nsew signal input
rlabel metal3 s -800 88816 800 88936 4 m_wbs_dat_o_9[11]
port 585 nsew signal input
rlabel metal3 s -800 89632 800 89752 4 m_wbs_dat_o_9[12]
port 586 nsew signal input
rlabel metal3 s -800 90584 800 90704 4 m_wbs_dat_o_9[13]
port 587 nsew signal input
rlabel metal3 s -800 91400 800 91520 4 m_wbs_dat_o_9[14]
port 588 nsew signal input
rlabel metal3 s -800 92216 800 92336 4 m_wbs_dat_o_9[15]
port 589 nsew signal input
rlabel metal3 s -800 93032 800 93152 4 m_wbs_dat_o_9[16]
port 590 nsew signal input
rlabel metal3 s -800 93848 800 93968 4 m_wbs_dat_o_9[17]
port 591 nsew signal input
rlabel metal3 s -800 94664 800 94784 4 m_wbs_dat_o_9[18]
port 592 nsew signal input
rlabel metal3 s -800 95480 800 95600 4 m_wbs_dat_o_9[19]
port 593 nsew signal input
rlabel metal3 s -800 80656 800 80776 4 m_wbs_dat_o_9[1]
port 594 nsew signal input
rlabel metal3 s -800 96296 800 96416 4 m_wbs_dat_o_9[20]
port 595 nsew signal input
rlabel metal3 s -800 97112 800 97232 4 m_wbs_dat_o_9[21]
port 596 nsew signal input
rlabel metal3 s -800 97928 800 98048 4 m_wbs_dat_o_9[22]
port 597 nsew signal input
rlabel metal3 s -800 98744 800 98864 4 m_wbs_dat_o_9[23]
port 598 nsew signal input
rlabel metal3 s -800 99560 800 99680 4 m_wbs_dat_o_9[24]
port 599 nsew signal input
rlabel metal3 s -800 100512 800 100632 4 m_wbs_dat_o_9[25]
port 600 nsew signal input
rlabel metal3 s -800 101328 800 101448 4 m_wbs_dat_o_9[26]
port 601 nsew signal input
rlabel metal3 s -800 102144 800 102264 4 m_wbs_dat_o_9[27]
port 602 nsew signal input
rlabel metal3 s -800 102960 800 103080 4 m_wbs_dat_o_9[28]
port 603 nsew signal input
rlabel metal3 s -800 103776 800 103896 4 m_wbs_dat_o_9[29]
port 604 nsew signal input
rlabel metal3 s -800 81472 800 81592 4 m_wbs_dat_o_9[2]
port 605 nsew signal input
rlabel metal3 s -800 104592 800 104712 4 m_wbs_dat_o_9[30]
port 606 nsew signal input
rlabel metal3 s -800 105408 800 105528 4 m_wbs_dat_o_9[31]
port 607 nsew signal input
rlabel metal3 s -800 82288 800 82408 4 m_wbs_dat_o_9[3]
port 608 nsew signal input
rlabel metal3 s -800 83104 800 83224 4 m_wbs_dat_o_9[4]
port 609 nsew signal input
rlabel metal3 s -800 83920 800 84040 4 m_wbs_dat_o_9[5]
port 610 nsew signal input
rlabel metal3 s -800 84736 800 84856 4 m_wbs_dat_o_9[6]
port 611 nsew signal input
rlabel metal3 s -800 85552 800 85672 4 m_wbs_dat_o_9[7]
port 612 nsew signal input
rlabel metal3 s -800 86368 800 86488 4 m_wbs_dat_o_9[8]
port 613 nsew signal input
rlabel metal3 s -800 87184 800 87304 4 m_wbs_dat_o_9[9]
port 614 nsew signal input
rlabel metal2 s 36726 119200 36782 120800 6 m_wbs_we_i
port 615 nsew signal tristate
rlabel metal2 s 25870 119200 25926 120800 6 mt_QEI_ChA_0
port 616 nsew signal tristate
rlabel metal2 s 26146 119200 26202 120800 6 mt_QEI_ChA_1
port 617 nsew signal tristate
rlabel metal2 s 26330 119200 26386 120800 6 mt_QEI_ChA_2
port 618 nsew signal tristate
rlabel metal2 s 26514 119200 26570 120800 6 mt_QEI_ChA_3
port 619 nsew signal tristate
rlabel metal2 s 26790 119200 26846 120800 6 mt_QEI_ChB_0
port 620 nsew signal tristate
rlabel metal2 s 26974 119200 27030 120800 6 mt_QEI_ChB_1
port 621 nsew signal tristate
rlabel metal2 s 27158 119200 27214 120800 6 mt_QEI_ChB_2
port 622 nsew signal tristate
rlabel metal2 s 27342 119200 27398 120800 6 mt_QEI_ChB_3
port 623 nsew signal tristate
rlabel metal2 s 27618 119200 27674 120800 6 mt_clo_test
port 624 nsew signal tristate
rlabel metal2 s 27802 119200 27858 120800 6 mt_pwm_h_0
port 625 nsew signal input
rlabel metal2 s 27986 119200 28042 120800 6 mt_pwm_h_1
port 626 nsew signal input
rlabel metal2 s 28262 119200 28318 120800 6 mt_pwm_h_2
port 627 nsew signal input
rlabel metal2 s 28446 119200 28502 120800 6 mt_pwm_h_3
port 628 nsew signal input
rlabel metal2 s 28630 119200 28686 120800 6 mt_pwm_l_0
port 629 nsew signal input
rlabel metal2 s 28906 119200 28962 120800 6 mt_pwm_l_1
port 630 nsew signal input
rlabel metal2 s 29090 119200 29146 120800 6 mt_pwm_l_2
port 631 nsew signal input
rlabel metal2 s 29274 119200 29330 120800 6 mt_pwm_l_3
port 632 nsew signal input
rlabel metal2 s 29458 119200 29514 120800 6 mt_pwm_test
port 633 nsew signal tristate
rlabel metal2 s 29918 119200 29974 120800 6 mt_sync_in[0]
port 634 nsew signal input
rlabel metal2 s 30102 119200 30158 120800 6 mt_sync_in[1]
port 635 nsew signal input
rlabel metal2 s 30378 119200 30434 120800 6 mt_sync_in[2]
port 636 nsew signal input
rlabel metal2 s 30562 119200 30618 120800 6 mt_sync_in[3]
port 637 nsew signal input
rlabel metal2 s 30746 119200 30802 120800 6 mt_sync_in[4]
port 638 nsew signal input
rlabel metal2 s 31022 119200 31078 120800 6 mt_sync_in[5]
port 639 nsew signal input
rlabel metal2 s 31206 119200 31262 120800 6 mt_sync_in[6]
port 640 nsew signal input
rlabel metal2 s 31390 119200 31446 120800 6 mt_sync_in[7]
port 641 nsew signal input
rlabel metal2 s 29734 119200 29790 120800 6 mt_sync_out
port 642 nsew signal tristate
rlabel metal2 s 110 -800 166 800 8 wb_clk_i
port 643 nsew signal input
rlabel metal2 s 386 -800 442 800 8 wb_rst_i
port 644 nsew signal input
rlabel metal2 s 1490 -800 1546 800 8 wbs_ack_o
port 645 nsew signal tristate
rlabel metal2 s 2686 -800 2742 800 8 wbs_adr_i[0]
port 646 nsew signal input
rlabel metal2 s 12622 -800 12678 800 8 wbs_adr_i[10]
port 647 nsew signal input
rlabel metal2 s 13542 -800 13598 800 8 wbs_adr_i[11]
port 648 nsew signal input
rlabel metal2 s 14370 -800 14426 800 8 wbs_adr_i[12]
port 649 nsew signal input
rlabel metal2 s 15290 -800 15346 800 8 wbs_adr_i[13]
port 650 nsew signal input
rlabel metal2 s 16118 -800 16174 800 8 wbs_adr_i[14]
port 651 nsew signal input
rlabel metal2 s 17038 -800 17094 800 8 wbs_adr_i[15]
port 652 nsew signal input
rlabel metal2 s 17866 -800 17922 800 8 wbs_adr_i[16]
port 653 nsew signal input
rlabel metal2 s 18786 -800 18842 800 8 wbs_adr_i[17]
port 654 nsew signal input
rlabel metal2 s 19614 -800 19670 800 8 wbs_adr_i[18]
port 655 nsew signal input
rlabel metal2 s 20534 -800 20590 800 8 wbs_adr_i[19]
port 656 nsew signal input
rlabel metal2 s 3882 -800 3938 800 8 wbs_adr_i[1]
port 657 nsew signal input
rlabel metal2 s 21362 -800 21418 800 8 wbs_adr_i[20]
port 658 nsew signal input
rlabel metal2 s 22282 -800 22338 800 8 wbs_adr_i[21]
port 659 nsew signal input
rlabel metal2 s 23110 -800 23166 800 8 wbs_adr_i[22]
port 660 nsew signal input
rlabel metal2 s 24030 -800 24086 800 8 wbs_adr_i[23]
port 661 nsew signal input
rlabel metal2 s 24858 -800 24914 800 8 wbs_adr_i[24]
port 662 nsew signal input
rlabel metal2 s 25778 -800 25834 800 8 wbs_adr_i[25]
port 663 nsew signal input
rlabel metal2 s 26606 -800 26662 800 8 wbs_adr_i[26]
port 664 nsew signal input
rlabel metal2 s 27526 -800 27582 800 8 wbs_adr_i[27]
port 665 nsew signal input
rlabel metal2 s 28354 -800 28410 800 8 wbs_adr_i[28]
port 666 nsew signal input
rlabel metal2 s 29274 -800 29330 800 8 wbs_adr_i[29]
port 667 nsew signal input
rlabel metal2 s 4986 -800 5042 800 8 wbs_adr_i[2]
port 668 nsew signal input
rlabel metal2 s 30194 -800 30250 800 8 wbs_adr_i[30]
port 669 nsew signal input
rlabel metal2 s 31022 -800 31078 800 8 wbs_adr_i[31]
port 670 nsew signal input
rlabel metal2 s 6182 -800 6238 800 8 wbs_adr_i[3]
port 671 nsew signal input
rlabel metal2 s 7378 -800 7434 800 8 wbs_adr_i[4]
port 672 nsew signal input
rlabel metal2 s 8206 -800 8262 800 8 wbs_adr_i[5]
port 673 nsew signal input
rlabel metal2 s 9126 -800 9182 800 8 wbs_adr_i[6]
port 674 nsew signal input
rlabel metal2 s 9954 -800 10010 800 8 wbs_adr_i[7]
port 675 nsew signal input
rlabel metal2 s 10874 -800 10930 800 8 wbs_adr_i[8]
port 676 nsew signal input
rlabel metal2 s 11794 -800 11850 800 8 wbs_adr_i[9]
port 677 nsew signal input
rlabel metal2 s 1858 -800 1914 800 8 wbs_cyc_i
port 678 nsew signal input
rlabel metal2 s 2962 -800 3018 800 8 wbs_dat_i[0]
port 679 nsew signal input
rlabel metal2 s 12898 -800 12954 800 8 wbs_dat_i[10]
port 680 nsew signal input
rlabel metal2 s 13818 -800 13874 800 8 wbs_dat_i[11]
port 681 nsew signal input
rlabel metal2 s 14646 -800 14702 800 8 wbs_dat_i[12]
port 682 nsew signal input
rlabel metal2 s 15566 -800 15622 800 8 wbs_dat_i[13]
port 683 nsew signal input
rlabel metal2 s 16394 -800 16450 800 8 wbs_dat_i[14]
port 684 nsew signal input
rlabel metal2 s 17314 -800 17370 800 8 wbs_dat_i[15]
port 685 nsew signal input
rlabel metal2 s 18142 -800 18198 800 8 wbs_dat_i[16]
port 686 nsew signal input
rlabel metal2 s 19062 -800 19118 800 8 wbs_dat_i[17]
port 687 nsew signal input
rlabel metal2 s 19890 -800 19946 800 8 wbs_dat_i[18]
port 688 nsew signal input
rlabel metal2 s 20810 -800 20866 800 8 wbs_dat_i[19]
port 689 nsew signal input
rlabel metal2 s 4158 -800 4214 800 8 wbs_dat_i[1]
port 690 nsew signal input
rlabel metal2 s 21638 -800 21694 800 8 wbs_dat_i[20]
port 691 nsew signal input
rlabel metal2 s 22558 -800 22614 800 8 wbs_dat_i[21]
port 692 nsew signal input
rlabel metal2 s 23478 -800 23534 800 8 wbs_dat_i[22]
port 693 nsew signal input
rlabel metal2 s 24306 -800 24362 800 8 wbs_dat_i[23]
port 694 nsew signal input
rlabel metal2 s 25226 -800 25282 800 8 wbs_dat_i[24]
port 695 nsew signal input
rlabel metal2 s 26054 -800 26110 800 8 wbs_dat_i[25]
port 696 nsew signal input
rlabel metal2 s 26974 -800 27030 800 8 wbs_dat_i[26]
port 697 nsew signal input
rlabel metal2 s 27802 -800 27858 800 8 wbs_dat_i[27]
port 698 nsew signal input
rlabel metal2 s 28722 -800 28778 800 8 wbs_dat_i[28]
port 699 nsew signal input
rlabel metal2 s 29550 -800 29606 800 8 wbs_dat_i[29]
port 700 nsew signal input
rlabel metal2 s 5354 -800 5410 800 8 wbs_dat_i[2]
port 701 nsew signal input
rlabel metal2 s 30470 -800 30526 800 8 wbs_dat_i[30]
port 702 nsew signal input
rlabel metal2 s 31298 -800 31354 800 8 wbs_dat_i[31]
port 703 nsew signal input
rlabel metal2 s 6458 -800 6514 800 8 wbs_dat_i[3]
port 704 nsew signal input
rlabel metal2 s 7654 -800 7710 800 8 wbs_dat_i[4]
port 705 nsew signal input
rlabel metal2 s 8574 -800 8630 800 8 wbs_dat_i[5]
port 706 nsew signal input
rlabel metal2 s 9402 -800 9458 800 8 wbs_dat_i[6]
port 707 nsew signal input
rlabel metal2 s 10322 -800 10378 800 8 wbs_dat_i[7]
port 708 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 wbs_dat_i[8]
port 709 nsew signal input
rlabel metal2 s 12070 -800 12126 800 8 wbs_dat_i[9]
port 710 nsew signal input
rlabel metal2 s 3238 -800 3294 800 8 wbs_dat_o[0]
port 711 nsew signal tristate
rlabel metal2 s 13174 -800 13230 800 8 wbs_dat_o[10]
port 712 nsew signal tristate
rlabel metal2 s 14094 -800 14150 800 8 wbs_dat_o[11]
port 713 nsew signal tristate
rlabel metal2 s 14922 -800 14978 800 8 wbs_dat_o[12]
port 714 nsew signal tristate
rlabel metal2 s 15842 -800 15898 800 8 wbs_dat_o[13]
port 715 nsew signal tristate
rlabel metal2 s 16670 -800 16726 800 8 wbs_dat_o[14]
port 716 nsew signal tristate
rlabel metal2 s 17590 -800 17646 800 8 wbs_dat_o[15]
port 717 nsew signal tristate
rlabel metal2 s 18510 -800 18566 800 8 wbs_dat_o[16]
port 718 nsew signal tristate
rlabel metal2 s 19338 -800 19394 800 8 wbs_dat_o[17]
port 719 nsew signal tristate
rlabel metal2 s 20258 -800 20314 800 8 wbs_dat_o[18]
port 720 nsew signal tristate
rlabel metal2 s 21086 -800 21142 800 8 wbs_dat_o[19]
port 721 nsew signal tristate
rlabel metal2 s 4434 -800 4490 800 8 wbs_dat_o[1]
port 722 nsew signal tristate
rlabel metal2 s 22006 -800 22062 800 8 wbs_dat_o[20]
port 723 nsew signal tristate
rlabel metal2 s 22834 -800 22890 800 8 wbs_dat_o[21]
port 724 nsew signal tristate
rlabel metal2 s 23754 -800 23810 800 8 wbs_dat_o[22]
port 725 nsew signal tristate
rlabel metal2 s 24582 -800 24638 800 8 wbs_dat_o[23]
port 726 nsew signal tristate
rlabel metal2 s 25502 -800 25558 800 8 wbs_dat_o[24]
port 727 nsew signal tristate
rlabel metal2 s 26330 -800 26386 800 8 wbs_dat_o[25]
port 728 nsew signal tristate
rlabel metal2 s 27250 -800 27306 800 8 wbs_dat_o[26]
port 729 nsew signal tristate
rlabel metal2 s 28078 -800 28134 800 8 wbs_dat_o[27]
port 730 nsew signal tristate
rlabel metal2 s 28998 -800 29054 800 8 wbs_dat_o[28]
port 731 nsew signal tristate
rlabel metal2 s 29826 -800 29882 800 8 wbs_dat_o[29]
port 732 nsew signal tristate
rlabel metal2 s 5630 -800 5686 800 8 wbs_dat_o[2]
port 733 nsew signal tristate
rlabel metal2 s 30746 -800 30802 800 8 wbs_dat_o[30]
port 734 nsew signal tristate
rlabel metal2 s 31574 -800 31630 800 8 wbs_dat_o[31]
port 735 nsew signal tristate
rlabel metal2 s 6826 -800 6882 800 8 wbs_dat_o[3]
port 736 nsew signal tristate
rlabel metal2 s 7930 -800 7986 800 8 wbs_dat_o[4]
port 737 nsew signal tristate
rlabel metal2 s 8850 -800 8906 800 8 wbs_dat_o[5]
port 738 nsew signal tristate
rlabel metal2 s 9678 -800 9734 800 8 wbs_dat_o[6]
port 739 nsew signal tristate
rlabel metal2 s 10598 -800 10654 800 8 wbs_dat_o[7]
port 740 nsew signal tristate
rlabel metal2 s 11426 -800 11482 800 8 wbs_dat_o[8]
port 741 nsew signal tristate
rlabel metal2 s 12346 -800 12402 800 8 wbs_dat_o[9]
port 742 nsew signal tristate
rlabel metal2 s 3606 -800 3662 800 8 wbs_sel_i[0]
port 743 nsew signal input
rlabel metal2 s 4710 -800 4766 800 8 wbs_sel_i[1]
port 744 nsew signal input
rlabel metal2 s 5906 -800 5962 800 8 wbs_sel_i[2]
port 745 nsew signal input
rlabel metal2 s 7102 -800 7158 800 8 wbs_sel_i[3]
port 746 nsew signal input
rlabel metal2 s 2134 -800 2190 800 8 wbs_stb_i
port 747 nsew signal input
rlabel metal2 s 2410 -800 2466 800 8 wbs_we_i
port 748 nsew signal input
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 749 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 750 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 751 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 120000
<< end >>
