* NGSPICE file created from cic_con.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt cic_con io_ack_o io_adr_i[0] io_adr_i[10] io_adr_i[11] io_adr_i[1] io_adr_i[2]
+ io_adr_i[3] io_adr_i[4] io_adr_i[5] io_adr_i[6] io_adr_i[7] io_adr_i[8] io_adr_i[9]
+ io_b_adr_i[0] io_b_adr_i[1] io_b_cs_i_0 io_b_cs_i_1 io_b_cs_i_10 io_b_cs_i_2 io_b_cs_i_3
+ io_b_cs_i_4 io_b_cs_i_5 io_b_cs_i_6 io_b_cs_i_7 io_b_cs_i_8 io_b_cs_i_9 io_b_dat_i[0]
+ io_b_dat_i[10] io_b_dat_i[11] io_b_dat_i[12] io_b_dat_i[13] io_b_dat_i[14] io_b_dat_i[15]
+ io_b_dat_i[1] io_b_dat_i[2] io_b_dat_i[3] io_b_dat_i[4] io_b_dat_i[5] io_b_dat_i[6]
+ io_b_dat_i[7] io_b_dat_i[8] io_b_dat_i[9] io_b_dat_o_0[0] io_b_dat_o_0[10] io_b_dat_o_0[11]
+ io_b_dat_o_0[12] io_b_dat_o_0[13] io_b_dat_o_0[14] io_b_dat_o_0[15] io_b_dat_o_0[1]
+ io_b_dat_o_0[2] io_b_dat_o_0[3] io_b_dat_o_0[4] io_b_dat_o_0[5] io_b_dat_o_0[6]
+ io_b_dat_o_0[7] io_b_dat_o_0[8] io_b_dat_o_0[9] io_b_dat_o_10[0] io_b_dat_o_10[10]
+ io_b_dat_o_10[11] io_b_dat_o_10[12] io_b_dat_o_10[13] io_b_dat_o_10[14] io_b_dat_o_10[15]
+ io_b_dat_o_10[1] io_b_dat_o_10[2] io_b_dat_o_10[3] io_b_dat_o_10[4] io_b_dat_o_10[5]
+ io_b_dat_o_10[6] io_b_dat_o_10[7] io_b_dat_o_10[8] io_b_dat_o_10[9] io_b_dat_o_1[0]
+ io_b_dat_o_1[10] io_b_dat_o_1[11] io_b_dat_o_1[12] io_b_dat_o_1[13] io_b_dat_o_1[14]
+ io_b_dat_o_1[15] io_b_dat_o_1[1] io_b_dat_o_1[2] io_b_dat_o_1[3] io_b_dat_o_1[4]
+ io_b_dat_o_1[5] io_b_dat_o_1[6] io_b_dat_o_1[7] io_b_dat_o_1[8] io_b_dat_o_1[9]
+ io_b_dat_o_2[0] io_b_dat_o_2[10] io_b_dat_o_2[11] io_b_dat_o_2[12] io_b_dat_o_2[13]
+ io_b_dat_o_2[14] io_b_dat_o_2[15] io_b_dat_o_2[1] io_b_dat_o_2[2] io_b_dat_o_2[3]
+ io_b_dat_o_2[4] io_b_dat_o_2[5] io_b_dat_o_2[6] io_b_dat_o_2[7] io_b_dat_o_2[8]
+ io_b_dat_o_2[9] io_b_dat_o_3[0] io_b_dat_o_3[10] io_b_dat_o_3[11] io_b_dat_o_3[12]
+ io_b_dat_o_3[13] io_b_dat_o_3[14] io_b_dat_o_3[15] io_b_dat_o_3[1] io_b_dat_o_3[2]
+ io_b_dat_o_3[3] io_b_dat_o_3[4] io_b_dat_o_3[5] io_b_dat_o_3[6] io_b_dat_o_3[7]
+ io_b_dat_o_3[8] io_b_dat_o_3[9] io_b_dat_o_4[0] io_b_dat_o_4[10] io_b_dat_o_4[11]
+ io_b_dat_o_4[12] io_b_dat_o_4[13] io_b_dat_o_4[14] io_b_dat_o_4[15] io_b_dat_o_4[1]
+ io_b_dat_o_4[2] io_b_dat_o_4[3] io_b_dat_o_4[4] io_b_dat_o_4[5] io_b_dat_o_4[6]
+ io_b_dat_o_4[7] io_b_dat_o_4[8] io_b_dat_o_4[9] io_b_dat_o_5[0] io_b_dat_o_5[10]
+ io_b_dat_o_5[11] io_b_dat_o_5[12] io_b_dat_o_5[13] io_b_dat_o_5[14] io_b_dat_o_5[15]
+ io_b_dat_o_5[1] io_b_dat_o_5[2] io_b_dat_o_5[3] io_b_dat_o_5[4] io_b_dat_o_5[5]
+ io_b_dat_o_5[6] io_b_dat_o_5[7] io_b_dat_o_5[8] io_b_dat_o_5[9] io_b_dat_o_6[0]
+ io_b_dat_o_6[10] io_b_dat_o_6[11] io_b_dat_o_6[12] io_b_dat_o_6[13] io_b_dat_o_6[14]
+ io_b_dat_o_6[15] io_b_dat_o_6[1] io_b_dat_o_6[2] io_b_dat_o_6[3] io_b_dat_o_6[4]
+ io_b_dat_o_6[5] io_b_dat_o_6[6] io_b_dat_o_6[7] io_b_dat_o_6[8] io_b_dat_o_6[9]
+ io_b_dat_o_7[0] io_b_dat_o_7[10] io_b_dat_o_7[11] io_b_dat_o_7[12] io_b_dat_o_7[13]
+ io_b_dat_o_7[14] io_b_dat_o_7[15] io_b_dat_o_7[1] io_b_dat_o_7[2] io_b_dat_o_7[3]
+ io_b_dat_o_7[4] io_b_dat_o_7[5] io_b_dat_o_7[6] io_b_dat_o_7[7] io_b_dat_o_7[8]
+ io_b_dat_o_7[9] io_b_dat_o_8[0] io_b_dat_o_8[10] io_b_dat_o_8[11] io_b_dat_o_8[12]
+ io_b_dat_o_8[13] io_b_dat_o_8[14] io_b_dat_o_8[15] io_b_dat_o_8[1] io_b_dat_o_8[2]
+ io_b_dat_o_8[3] io_b_dat_o_8[4] io_b_dat_o_8[5] io_b_dat_o_8[6] io_b_dat_o_8[7]
+ io_b_dat_o_8[8] io_b_dat_o_8[9] io_b_dat_o_9[0] io_b_dat_o_9[10] io_b_dat_o_9[11]
+ io_b_dat_o_9[12] io_b_dat_o_9[13] io_b_dat_o_9[14] io_b_dat_o_9[15] io_b_dat_o_9[1]
+ io_b_dat_o_9[2] io_b_dat_o_9[3] io_b_dat_o_9[4] io_b_dat_o_9[5] io_b_dat_o_9[6]
+ io_b_dat_o_9[7] io_b_dat_o_9[8] io_b_dat_o_9[9] io_b_we_i io_cs_i io_dat_i[0] io_dat_i[10]
+ io_dat_i[11] io_dat_i[12] io_dat_i[13] io_dat_i[14] io_dat_i[15] io_dat_i[16] io_dat_i[17]
+ io_dat_i[18] io_dat_i[19] io_dat_i[1] io_dat_i[20] io_dat_i[21] io_dat_i[22] io_dat_i[23]
+ io_dat_i[24] io_dat_i[25] io_dat_i[26] io_dat_i[27] io_dat_i[28] io_dat_i[29] io_dat_i[2]
+ io_dat_i[30] io_dat_i[31] io_dat_i[3] io_dat_i[4] io_dat_i[5] io_dat_i[6] io_dat_i[7]
+ io_dat_i[8] io_dat_i[9] io_dat_o[0] io_dat_o[10] io_dat_o[11] io_dat_o[12] io_dat_o[13]
+ io_dat_o[14] io_dat_o[15] io_dat_o[16] io_dat_o[17] io_dat_o[18] io_dat_o[19] io_dat_o[1]
+ io_dat_o[20] io_dat_o[21] io_dat_o[22] io_dat_o[23] io_dat_o[24] io_dat_o[25] io_dat_o[26]
+ io_dat_o[27] io_dat_o[28] io_dat_o[29] io_dat_o[2] io_dat_o[30] io_dat_o[31] io_dat_o[3]
+ io_dat_o[4] io_dat_o[5] io_dat_o[6] io_dat_o[7] io_dat_o[8] io_dat_o[9] io_dataLastBlock[0]
+ io_dataLastBlock[10] io_dataLastBlock[11] io_dataLastBlock[12] io_dataLastBlock[13]
+ io_dataLastBlock[14] io_dataLastBlock[15] io_dataLastBlock[16] io_dataLastBlock[17]
+ io_dataLastBlock[18] io_dataLastBlock[19] io_dataLastBlock[1] io_dataLastBlock[20]
+ io_dataLastBlock[21] io_dataLastBlock[22] io_dataLastBlock[23] io_dataLastBlock[24]
+ io_dataLastBlock[25] io_dataLastBlock[26] io_dataLastBlock[27] io_dataLastBlock[28]
+ io_dataLastBlock[29] io_dataLastBlock[2] io_dataLastBlock[30] io_dataLastBlock[31]
+ io_dataLastBlock[32] io_dataLastBlock[33] io_dataLastBlock[34] io_dataLastBlock[35]
+ io_dataLastBlock[36] io_dataLastBlock[37] io_dataLastBlock[38] io_dataLastBlock[39]
+ io_dataLastBlock[3] io_dataLastBlock[40] io_dataLastBlock[41] io_dataLastBlock[42]
+ io_dataLastBlock[43] io_dataLastBlock[44] io_dataLastBlock[45] io_dataLastBlock[46]
+ io_dataLastBlock[47] io_dataLastBlock[48] io_dataLastBlock[49] io_dataLastBlock[4]
+ io_dataLastBlock[50] io_dataLastBlock[51] io_dataLastBlock[52] io_dataLastBlock[53]
+ io_dataLastBlock[54] io_dataLastBlock[55] io_dataLastBlock[56] io_dataLastBlock[57]
+ io_dataLastBlock[58] io_dataLastBlock[59] io_dataLastBlock[5] io_dataLastBlock[60]
+ io_dataLastBlock[61] io_dataLastBlock[62] io_dataLastBlock[63] io_dataLastBlock[6]
+ io_dataLastBlock[7] io_dataLastBlock[8] io_dataLastBlock[9] io_dsi_in[0] io_dsi_in[1]
+ io_dsi_in[2] io_dsi_in[3] io_dsi_in[4] io_dsi_in[5] io_dsi_in[6] io_dsi_in[7] io_dsi_o
+ io_irq io_sync_out io_vout[0] io_vout[10] io_vout[1] io_vout[2] io_vout[3] io_vout[4]
+ io_vout[5] io_vout[6] io_vout[7] io_vout[8] io_vout[9] io_we_i wb_clk_i wb_rst_i
+ vccd1 vssd1
XFILLER_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3155_ _3180_/CLK _3155_/D vssd1 vssd1 vccd1 vccd1 _3155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2106_ _2190_/A _2544_/A vssd1 vssd1 vccd1 vccd1 _2122_/A sky130_fd_sc_hd__or2_4
X_3086_ _3087_/CLK _3086_/D vssd1 vssd1 vccd1 vccd1 _3086_/Q sky130_fd_sc_hd__dfxtp_1
X_2037_ _3245_/Q _2031_/X _1967_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2939_ _3093_/Q _3069_/Q _3045_/Q _3349_/Q _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2939_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_60_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3301_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2724_ _3144_/Q _3120_/Q _3192_/Q _3440_/Q _2750_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2724_/X sky130_fd_sc_hd__mux4_1
X_2655_ _2906_/X _2654_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__mux2_2
X_1606_ _1609_/A _2961_/X vssd1 vssd1 vccd1 vccd1 _3460_/D sky130_fd_sc_hd__and2_1
X_2586_ _2585_/X _2493_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__mux2_1
X_1537_ _1626_/D _1678_/D vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__or2_4
XFILLER_47_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3207_ _3279_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3138_ _3346_/CLK _3138_/D vssd1 vssd1 vccd1 vccd1 _3138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3069_ _3437_/CLK _3069_/D vssd1 vssd1 vccd1 vccd1 _3069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2440_ _3414_/Q vssd1 vssd1 vccd1 vccd1 _2440_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2371_ _3037_/Q _2367_/X _2332_/X _2368_/X vssd1 vssd1 vccd1 vccd1 _3037_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2707_ _2703_/X _2704_/X _2705_/X _2706_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2707_/X sky130_fd_sc_hd__mux4_2
X_2638_ _2856_/X _2857_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__mux2_1
X_2569_ _2569_/A vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__buf_1
XINSDIODE2_4 _2759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput297 _2556_/X vssd1 vssd1 vccd1 vccd1 io_b_adr_i[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_75_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1940_ _3304_/Q _1931_/X _1939_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _3304_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1871_ _3345_/Q _1864_/A _1826_/X _1865_/A vssd1 vssd1 vccd1 vccd1 _3345_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3472_ _3500_/CLK _3472_/D vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfxtp_1
X_2423_ _2430_/A _2611_/X vssd1 vssd1 vccd1 vccd1 _2423_/X sky130_fd_sc_hd__and2_1
X_2354_ _3050_/Q _2351_/X _2330_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3050_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2285_ _3093_/Q _2282_/X _2250_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _3093_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2070_ _3226_/Q _2063_/A _2053_/X _2064_/A vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ input21/X input53/X input69/X input85/X _2610_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2972_/X sky130_fd_sc_hd__mux4_1
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1923_ _1943_/A vssd1 vssd1 vccd1 vccd1 _1945_/A sky130_fd_sc_hd__inv_2
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1854_ _3358_/Q _1849_/X _1636_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__a22o_1
X_1785_ _3392_/Q _1782_/X _1770_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__a22o_1
X_3455_ _3455_/CLK _3455_/D vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfxtp_1
X_2406_ _3008_/Q _1736_/X _2038_/A _1738_/X vssd1 vssd1 vccd1 vccd1 _3008_/D sky130_fd_sc_hd__a22o_1
X_3386_ _3420_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
X_2337_ _3059_/Q _2326_/X _2336_/X _2328_/X vssd1 vssd1 vccd1 vccd1 _3059_/D sky130_fd_sc_hd__a22o_1
X_2268_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__inv_2
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2199_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3485_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ _1582_/A vssd1 vssd1 vccd1 vccd1 _1575_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3240_ _3307_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
X_3171_ _3335_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2122_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2053_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2053_/X sky130_fd_sc_hd__buf_2
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _3380_/Q _3416_/Q _3432_/Q _3428_/Q _2610_/S _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2955_/X sky130_fd_sc_hd__mux4_2
X_2886_ input28/X input60/X input76/X input92/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2886_/X sky130_fd_sc_hd__mux4_1
X_1906_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1906_/X sky130_fd_sc_hd__clkbuf_2
X_1837_ _1837_/A vssd1 vssd1 vccd1 vccd1 _1837_/X sky130_fd_sc_hd__buf_2
X_3507_ _3509_/CLK _3507_/D vssd1 vssd1 vccd1 vccd1 _3507_/Q sky130_fd_sc_hd__dfxtp_1
X_1768_ _2224_/A _1798_/B _2224_/C _1828_/B vssd1 vssd1 vccd1 vccd1 _2377_/A sky130_fd_sc_hd__or4_4
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1699_ _3425_/Q _1693_/X _1670_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3438_ _3438_/CLK _3438_/D vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfxtp_1
X_3369_ _3371_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater383 _2992_/S1 vssd1 vssd1 vccd1 vccd1 _2997_/S1 sky130_fd_sc_hd__buf_8
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater394 _1700_/B vssd1 vssd1 vccd1 vccd1 _2611_/S sky130_fd_sc_hd__buf_8
XFILLER_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput120 io_b_dat_o_5[5] vssd1 vssd1 vccd1 vccd1 _2934_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput142 io_b_dat_o_7[10] vssd1 vssd1 vccd1 vccd1 _2879_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput131 io_b_dat_o_6[15] vssd1 vssd1 vccd1 vccd1 _2854_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput153 io_b_dat_o_7[6] vssd1 vssd1 vccd1 vccd1 _2921_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput175 io_b_dat_o_9[11] vssd1 vssd1 vccd1 vccd1 _2588_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput186 io_b_dat_o_9[7] vssd1 vssd1 vccd1 vccd1 _2596_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput164 io_b_dat_o_8[1] vssd1 vssd1 vccd1 vccd1 _2608_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput197 io_dat_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_1
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ _3243_/Q _3219_/Q _3291_/Q _3267_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2740_/X sky130_fd_sc_hd__mux4_2
X_2671_ _2958_/X _2670_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2671_/X sky130_fd_sc_hd__mux2_1
X_1622_ _1676_/A vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__inv_2
X_1553_ _3497_/Q _1539_/A _1939_/A _1541_/A _1544_/X vssd1 vssd1 vccd1 vccd1 _3497_/D
+ sky130_fd_sc_hd__o221a_1
X_1484_ _1484_/A vssd1 vssd1 vccd1 vccd1 _1484_/Y sky130_fd_sc_hd__inv_2
X_3223_ _3296_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3154_ _3501_/CLK _3154_/D vssd1 vssd1 vccd1 vccd1 _3154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2105_ _3201_/Q _2097_/A _2056_/X _2098_/A vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__a22o_1
X_3085_ _3371_/CLK _3085_/D vssd1 vssd1 vccd1 vccd1 _3085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2036_ _3246_/Q _2031_/X _1965_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _3246_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2938_ _3189_/Q _3437_/Q _3141_/Q _3117_/Q _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2938_/X sky130_fd_sc_hd__mux4_1
X_2869_ _2865_/X _2866_/X _2867_/X _2868_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2869_/X sky130_fd_sc_hd__mux4_2
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2723_ _3048_/Q _3352_/Q _3096_/Q _3072_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2723_/X sky130_fd_sc_hd__mux4_2
X_2654_ _2654_/A0 _2654_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2654_/X sky130_fd_sc_hd__mux2_1
X_2585_ _2585_/A0 _2585_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__mux2_1
X_1605_ _1609_/A _2948_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__and2_1
X_1536_ _2683_/S input3/X input2/X vssd1 vssd1 vccd1 vccd1 _1678_/D sky130_fd_sc_hd__or3_1
XFILLER_86_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _3279_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3137_ _3433_/CLK _3137_/D vssd1 vssd1 vccd1 vccd1 _3137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3068_ _3392_/CLK _3068_/D vssd1 vssd1 vccd1 vccd1 _3068_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2019_ _3256_/Q _1817_/X _1929_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _3256_/D sky130_fd_sc_hd__a22o_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2370_ _3038_/Q _2367_/X _2330_/X _2368_/X vssd1 vssd1 vccd1 vccd1 _3038_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _3316_/Q _3300_/Q _3164_/Q _3332_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2706_/X sky130_fd_sc_hd__mux4_1
X_2637_ _2853_/X _2854_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2637_/X sky130_fd_sc_hd__mux2_1
X_2568_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__clkbuf_1
X_2499_ _2522_/A _2499_/B vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__and2_1
XINSDIODE2_5 _3467_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput298 _2557_/X vssd1 vssd1 vccd1 vccd1 io_b_adr_i[1] sky130_fd_sc_hd__clkbuf_2
X_1519_ _1515_/X _3512_/Q _1516_/X _2737_/X _1510_/X vssd1 vssd1 vccd1 vccd1 _3512_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_39_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3303_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1870_ _3346_/Q _1864_/X _1824_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3471_ _3482_/CLK _3471_/D vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfxtp_1
X_2422_ _2429_/A _2422_/B vssd1 vssd1 vccd1 vccd1 _2422_/X sky130_fd_sc_hd__and2_1
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2353_ _3051_/Q _2351_/X _2327_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3051_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ _3094_/Q _2282_/X _2247_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _3094_/D sky130_fd_sc_hd__a22o_1
XFILLER_64_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1999_ _3272_/Q _1996_/X _1959_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2971_ _2967_/X _2968_/X _2969_/X _2970_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2971_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1922_ _1943_/A vssd1 vssd1 vccd1 vccd1 _1922_/X sky130_fd_sc_hd__clkbuf_2
X_1853_ _3359_/Q _1849_/X _1634_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__a22o_1
X_1784_ _2064_/A vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3454_ _3455_/CLK _3454_/D vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfxtp_1
X_2405_ _3009_/Q _2397_/A _1947_/A _2398_/A vssd1 vssd1 vccd1 vccd1 _3009_/D sky130_fd_sc_hd__a22o_1
X_3385_ _3392_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
X_2336_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2336_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2267_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2198_ _3148_/Q _2191_/X _2134_/X _2193_/X vssd1 vssd1 vccd1 vccd1 _3148_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_54_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3502_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3170_ _3504_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
X_2121_ _3191_/Q _2115_/X _2050_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2052_ _2052_/A vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2954_ _3420_/Q _3376_/Q _3392_/Q _3388_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2954_/X sky130_fd_sc_hd__mux4_2
X_2885_ _2881_/X _2882_/X _2883_/X _2884_/X _2660_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2885_/X sky130_fd_sc_hd__mux4_1
X_1905_ _3324_/Q _1898_/X _1641_/X _1900_/X vssd1 vssd1 vccd1 vccd1 _3324_/D sky130_fd_sc_hd__a22o_1
X_1836_ _3368_/Q _1829_/X _1654_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__a22o_1
X_1767_ _3397_/Q _1761_/X _1730_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__a22o_1
X_3506_ _3506_/CLK _3506_/D vssd1 vssd1 vccd1 vccd1 _3506_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _3426_/Q _1693_/X _1668_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__a22o_1
X_3437_ _3437_/CLK _3437_/D vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfxtp_1
X_3368_ _3371_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
X_2319_ _3069_/Q _2316_/X _2250_/X _2317_/X vssd1 vssd1 vccd1 vccd1 _3069_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3299_ _3331_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater373 _2847_/X vssd1 vssd1 vccd1 vccd1 _2751_/S1 sky130_fd_sc_hd__buf_8
Xrepeater384 input8/X vssd1 vssd1 vccd1 vccd1 _2992_/S1 sky130_fd_sc_hd__buf_6
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater395 _1700_/B vssd1 vssd1 vccd1 vccd1 _2944_/S1 sky130_fd_sc_hd__buf_8
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput110 io_b_dat_o_5[10] vssd1 vssd1 vccd1 vccd1 _2879_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput143 io_b_dat_o_7[11] vssd1 vssd1 vccd1 vccd1 _2871_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput154 io_b_dat_o_7[7] vssd1 vssd1 vccd1 vccd1 _2908_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput121 io_b_dat_o_5[6] vssd1 vssd1 vccd1 vccd1 _2921_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput132 io_b_dat_o_6[1] vssd1 vssd1 vccd1 vccd1 _2986_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput176 io_b_dat_o_9[12] vssd1 vssd1 vccd1 vccd1 _2585_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput187 io_b_dat_o_9[8] vssd1 vssd1 vccd1 vccd1 _2594_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput165 io_b_dat_o_8[2] vssd1 vssd1 vccd1 vccd1 _2606_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput198 io_dat_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__buf_1
XFILLER_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _2670_/A0 _2670_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2670_/X sky130_fd_sc_hd__mux2_4
X_1621_ input8/X vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__inv_2
X_1552_ _2565_/A vssd1 vssd1 vccd1 vccd1 _1939_/A sky130_fd_sc_hd__buf_2
X_1483_ _3518_/Q _1483_/B vssd1 vssd1 vccd1 vccd1 _1484_/A sky130_fd_sc_hd__nand2_1
X_3222_ _3294_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
X_3153_ _3501_/CLK _3153_/D vssd1 vssd1 vccd1 vccd1 _3153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2104_ _3202_/Q _2097_/A _2053_/X _2098_/A vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _3109_/CLK _3084_/D vssd1 vssd1 vccd1 vccd1 _3084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2035_ _3247_/Q _2031_/X _1963_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2937_ _3285_/Q _3261_/Q _3237_/Q _3213_/Q _1700_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2937_/X sky130_fd_sc_hd__mux4_2
X_2868_ _3024_/Q _3016_/Q _3008_/Q _3280_/Q _2982_/S0 _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2868_/X sky130_fd_sc_hd__mux4_1
X_2799_ _3183_/Q _3159_/Q _3135_/Q _3111_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2799_/X sky130_fd_sc_hd__mux4_1
X_1819_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2021_/A sky130_fd_sc_hd__inv_2
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2722_ _2718_/X _2719_/X _2720_/X _2721_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2722_/X sky130_fd_sc_hd__mux4_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2653_ _3497_/Q _2901_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__mux2_1
X_1604_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1609_/A sky130_fd_sc_hd__buf_1
X_2584_ _2584_/A0 _2584_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__mux2_1
X_1535_ _2540_/A _1678_/B _2557_/A vssd1 vssd1 vccd1 vccd1 _1626_/D sky130_fd_sc_hd__or3_1
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3205_ _3279_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_1
X_3136_ _3500_/CLK _3136_/D vssd1 vssd1 vccd1 vccd1 _3136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3067_ _3392_/CLK _3067_/D vssd1 vssd1 vccd1 vccd1 _3067_/Q sky130_fd_sc_hd__dfxtp_1
X_2018_ _3257_/Q _2011_/A _1955_/X _2012_/A vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__a22o_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_9_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3420_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2705_ _3236_/Q _3212_/Q _3284_/Q _3260_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2705_/X sky130_fd_sc_hd__mux4_2
X_2636_ _2636_/A0 _2636_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__mux2_2
X_2567_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_6 _1610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2498_ _2509_/A _2584_/X vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__and2_1
X_1518_ _1515_/X _3513_/Q _1516_/X _2742_/X _1510_/X vssd1 vssd1 vccd1 vccd1 _3513_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput299 _2553_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_0 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3119_ _3439_/CLK _3119_/D vssd1 vssd1 vccd1 vccd1 _3119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ _3482_/CLK _3470_/D vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfxtp_1
X_2421_ _2430_/A _2609_/X vssd1 vssd1 vccd1 vccd1 _2421_/X sky130_fd_sc_hd__and2_1
X_2352_ _2359_/A vssd1 vssd1 vccd1 vccd1 _2352_/X sky130_fd_sc_hd__clkbuf_2
X_2283_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1998_ _2012_/A vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__clkbuf_2
X_2619_ _2529_/X _2827_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2970_ _3407_/Q _3403_/Q _3411_/Q _3383_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2970_/X sky130_fd_sc_hd__mux4_1
X_1921_ _1995_/A _2550_/A vssd1 vssd1 vccd1 vccd1 _1943_/A sky130_fd_sc_hd__or2_4
X_1852_ _3360_/Q _1849_/X _1630_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1783_ _2063_/A vssd1 vssd1 vccd1 vccd1 _2064_/A sky130_fd_sc_hd__inv_2
X_3453_ _3456_/CLK _3453_/D vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfxtp_1
X_2404_ _3010_/Q _2397_/A _1944_/A _2398_/A vssd1 vssd1 vccd1 vccd1 _3010_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3384_ _3409_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2335_ _3060_/Q _2326_/X _2334_/X _2328_/X vssd1 vssd1 vccd1 vccd1 _3060_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2266_ _2342_/A _2342_/B _2266_/C _2300_/D vssd1 vssd1 vccd1 vccd1 _2282_/A sky130_fd_sc_hd__or4_4
X_2197_ _3149_/Q _2191_/X _2162_/X _2193_/X vssd1 vssd1 vccd1 vccd1 _3149_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _3192_/Q _2115_/X _2048_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__a22o_1
X_2051_ _3239_/Q _2040_/X _2050_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _2949_/X _2950_/X _2951_/X _2952_/X input7/X input8/X vssd1 vssd1 vccd1 vccd1
+ _2953_/X sky130_fd_sc_hd__mux4_2
X_1904_ _3325_/Q _1898_/X _1638_/X _1900_/X vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__a22o_1
X_2884_ _3022_/Q _3014_/Q _3006_/Q _3278_/Q _2644_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2884_/X sky130_fd_sc_hd__mux4_1
X_1835_ _3369_/Q _1829_/X _1652_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__a22o_1
X_1766_ _3398_/Q _1761_/X _1728_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__a22o_1
X_3505_ _3506_/CLK _3505_/D vssd1 vssd1 vccd1 vccd1 _3505_/Q sky130_fd_sc_hd__dfxtp_1
X_1697_ _3427_/Q _1693_/X _1666_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__a22o_1
X_3436_ _3437_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
X_3367_ _3367_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
X_2318_ _3070_/Q _2316_/X _2247_/X _2317_/X vssd1 vssd1 vccd1 vccd1 _3070_/D sky130_fd_sc_hd__a22o_1
X_3298_ _3331_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater385 _2660_/S vssd1 vssd1 vccd1 vccd1 _2684_/S sky130_fd_sc_hd__buf_8
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater374 _2847_/X vssd1 vssd1 vccd1 vccd1 _2716_/S1 sky130_fd_sc_hd__buf_8
X_2249_ _3118_/Q _2246_/X _2247_/X _2248_/X vssd1 vssd1 vccd1 vccd1 _3118_/D sky130_fd_sc_hd__a22o_1
Xrepeater396 _1700_/B vssd1 vssd1 vccd1 vccd1 _2991_/S1 sky130_fd_sc_hd__buf_6
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput111 io_b_dat_o_5[11] vssd1 vssd1 vccd1 vccd1 _2871_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput100 io_b_dat_o_4[1] vssd1 vssd1 vccd1 vccd1 _2986_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput144 io_b_dat_o_7[12] vssd1 vssd1 vccd1 vccd1 _2863_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput133 io_b_dat_o_6[2] vssd1 vssd1 vccd1 vccd1 _2973_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput122 io_b_dat_o_5[7] vssd1 vssd1 vccd1 vccd1 _2908_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput166 io_b_dat_o_8[3] vssd1 vssd1 vccd1 vccd1 _2604_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput177 io_b_dat_o_9[13] vssd1 vssd1 vccd1 vccd1 _2582_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput155 io_b_dat_o_7[8] vssd1 vssd1 vccd1 vccd1 _2895_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput188 io_b_dat_o_9[9] vssd1 vssd1 vccd1 vccd1 _2592_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput199 io_dat_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__buf_1
XFILLER_44_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1620_ _1815_/A vssd1 vssd1 vccd1 vccd1 _2224_/A sky130_fd_sc_hd__clkbuf_2
X_1551_ _3498_/Q _1539_/X _1728_/A _1541_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _3498_/D
+ sky130_fd_sc_hd__o221a_1
X_1482_ _1482_/A _1482_/B vssd1 vssd1 vccd1 vccd1 _1483_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3221_ _3294_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3152_ _3447_/CLK _3152_/D vssd1 vssd1 vccd1 vccd1 _3152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2103_ _3203_/Q _2097_/X _2050_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__a22o_1
X_3083_ _3275_/CLK _3083_/D vssd1 vssd1 vccd1 vccd1 _3083_/Q sky130_fd_sc_hd__dfxtp_1
X_2034_ _3248_/Q _2031_/X _1959_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _3248_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2936_ _3165_/Q _3333_/Q _3317_/Q _3301_/Q _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2936_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2867_ _3088_/Q _3372_/Q _3040_/Q _3032_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2867_/X sky130_fd_sc_hd__mux4_1
X_1818_ _2561_/A vssd1 vssd1 vccd1 vccd1 _1818_/X sky130_fd_sc_hd__clkbuf_2
X_2798_ _3063_/Q _3255_/Q _3231_/Q _3207_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2798_/X sky130_fd_sc_hd__mux4_2
X_1749_ _3406_/Q _1744_/X _1728_/X _1746_/X vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3419_ _3423_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ _3319_/Q _3303_/Q _3167_/Q _3335_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2721_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2894_/X _2895_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2583_ _2582_/X _2499_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__mux2_1
X_1603_ _1603_/A _2935_/X vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__and2_1
X_1534_ _2574_/A vssd1 vssd1 vccd1 vccd1 _1678_/B sky130_fd_sc_hd__inv_2
XFILLER_87_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3204_ _3279_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_1
X_3135_ _3456_/CLK _3135_/D vssd1 vssd1 vccd1 vccd1 _3135_/Q sky130_fd_sc_hd__dfxtp_1
X_3066_ _3346_/CLK _3066_/D vssd1 vssd1 vccd1 vccd1 _3066_/Q sky130_fd_sc_hd__dfxtp_1
X_2017_ _3258_/Q _2011_/X _1953_/X _2012_/X vssd1 vssd1 vccd1 vccd1 _3258_/D sky130_fd_sc_hd__a22o_1
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
X_2919_ _2915_/X _2916_/X _2917_/X _2918_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2919_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _3140_/Q _3116_/Q _3188_/Q _3436_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2704_/X sky130_fd_sc_hd__mux4_2
X_2635_ _2635_/A0 _2635_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2635_/X sky130_fd_sc_hd__mux2_1
X_2566_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_7 _2487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2497_ _2509_/A _2767_/X vssd1 vssd1 vccd1 vccd1 _2497_/X sky130_fd_sc_hd__and2_1
X_1517_ _1515_/X _3514_/Q _1516_/X _2747_/X _1510_/X vssd1 vssd1 vccd1 vccd1 _3514_/D
+ sky130_fd_sc_hd__o221a_1
X_3118_ _3438_/CLK _3118_/D vssd1 vssd1 vccd1 vccd1 _3118_/Q sky130_fd_sc_hd__dfxtp_1
X_3049_ _3353_/CLK _3049_/D vssd1 vssd1 vccd1 vccd1 _3049_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3447_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2420_ _2487_/A vssd1 vssd1 vccd1 vccd1 _2430_/A sky130_fd_sc_hd__buf_1
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2351_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__clkbuf_2
X_2282_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2282_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1997_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2012_/A sky130_fd_sc_hd__inv_2
X_2618_ _2530_/X _2822_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2618_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2549_ _2549_/A _2552_/B vssd1 vssd1 vccd1 vccd1 _2549_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1920_ _3313_/Q _1913_/A _1826_/X _1914_/A vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__a22o_1
X_1851_ _1865_/A vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__buf_2
X_1782_ _2063_/A vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__clkbuf_2
X_3452_ _3456_/CLK _3452_/D vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2403_ _3011_/Q _2397_/X _1941_/A _2398_/X vssd1 vssd1 vccd1 vccd1 _3011_/D sky130_fd_sc_hd__a22o_1
X_3383_ _3409_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
X_2334_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2334_/X sky130_fd_sc_hd__clkbuf_2
X_2265_ _3105_/Q _2257_/A _2250_/X _2258_/A vssd1 vssd1 vccd1 vccd1 _3105_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2196_ _3150_/Q _2191_/X _2160_/X _2193_/X vssd1 vssd1 vccd1 vccd1 _3150_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2050_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2050_/X sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_63_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3331_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2952_ _3092_/Q _3068_/Q _3044_/Q _3348_/Q _1676_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2952_/X sky130_fd_sc_hd__mux4_2
X_1903_ _3326_/Q _1898_/X _1636_/X _1900_/X vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__a22o_1
X_2883_ _3086_/Q _3370_/Q _3038_/Q _3030_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2883_/X sky130_fd_sc_hd__mux4_2
X_1834_ _3370_/Q _1829_/X _1649_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__a22o_1
X_1765_ _3399_/Q _1761_/X _1726_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3504_ _3504_/CLK _3504_/D vssd1 vssd1 vccd1 vccd1 _3504_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _3428_/Q _1693_/X _1664_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__a22o_1
X_3435_ _3437_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_3366_ _3367_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
X_3297_ _3297_/CLK _3297_/D vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
X_2317_ _2317_/A vssd1 vssd1 vccd1 vccd1 _2317_/X sky130_fd_sc_hd__clkbuf_2
X_2248_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater375 _2842_/X vssd1 vssd1 vccd1 vccd1 _2752_/S0 sky130_fd_sc_hd__buf_12
Xrepeater386 _2901_/S0 vssd1 vssd1 vccd1 vccd1 _2660_/S sky130_fd_sc_hd__buf_8
XFILLER_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2179_ _3161_/Q _2172_/A _2132_/X _2173_/A vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater397 input6/X vssd1 vssd1 vccd1 vccd1 _1700_/B sky130_fd_sc_hd__buf_8
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput101 io_b_dat_o_4[2] vssd1 vssd1 vccd1 vccd1 _2973_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput145 io_b_dat_o_7[13] vssd1 vssd1 vccd1 vccd1 _2860_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput123 io_b_dat_o_5[8] vssd1 vssd1 vccd1 vccd1 _2895_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput134 io_b_dat_o_6[3] vssd1 vssd1 vccd1 vccd1 _2960_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput112 io_b_dat_o_5[12] vssd1 vssd1 vccd1 vccd1 _2863_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput156 io_b_dat_o_7[9] vssd1 vssd1 vccd1 vccd1 _2887_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput178 io_b_dat_o_9[14] vssd1 vssd1 vccd1 vccd1 _2579_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput167 io_b_dat_o_8[4] vssd1 vssd1 vccd1 vccd1 _2602_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput189 io_cs_i vssd1 vssd1 vccd1 vccd1 _1533_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_91_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _2559_/A vssd1 vssd1 vccd1 vccd1 _1728_/A sky130_fd_sc_hd__buf_2
X_1481_ _3516_/Q vssd1 vssd1 vccd1 vccd1 _1482_/B sky130_fd_sc_hd__inv_2
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3220_ _3297_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
X_3151_ _3447_/CLK _3151_/D vssd1 vssd1 vccd1 vccd1 _3151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2102_ _3204_/Q _2097_/X _2048_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__a22o_1
X_3082_ _3273_/CLK _3082_/D vssd1 vssd1 vccd1 vccd1 _3082_/Q sky130_fd_sc_hd__dfxtp_1
X_2033_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2033_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2935_ _2661_/X _2663_/X _2664_/X _2430_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2935_/X sky130_fd_sc_hd__mux4_2
X_2866_ _3184_/Q _3160_/Q _3136_/Q _3112_/Q _2982_/S0 _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2866_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1817_ _2020_/A vssd1 vssd1 vccd1 vccd1 _1817_/X sky130_fd_sc_hd__clkbuf_2
X_2797_ _2793_/X _2794_/X _2795_/X _2796_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2797_/X sky130_fd_sc_hd__mux4_2
X_1748_ _3407_/Q _1744_/X _1726_/X _1746_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1679_ _1798_/D vssd1 vssd1 vccd1 vccd1 _1816_/A sky130_fd_sc_hd__buf_1
X_3418_ _3420_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
X_3349_ _3437_/CLK _3349_/D vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _3239_/Q _3215_/Q _3287_/Q _3263_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2720_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2651_ _2893_/X _2650_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2651_/X sky130_fd_sc_hd__mux2_2
X_1602_ _1603_/A _2922_/X vssd1 vssd1 vccd1 vccd1 _3463_/D sky130_fd_sc_hd__and2_1
X_2582_ _2582_/A0 _2582_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1533_ _1533_/A vssd1 vssd1 vccd1 vccd1 _2540_/A sky130_fd_sc_hd__inv_2
XFILLER_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3203_ _3371_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_1
X_3134_ _3456_/CLK _3134_/D vssd1 vssd1 vccd1 vccd1 _3134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3065_ _3502_/CLK _3065_/D vssd1 vssd1 vccd1 vccd1 _3065_/Q sky130_fd_sc_hd__dfxtp_1
X_2016_ _3259_/Q _2011_/X _1951_/X _2012_/X vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2918_ _3019_/Q _3011_/Q _3003_/Q _3275_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2918_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2849_ _3377_/Q _3413_/Q _3429_/Q _3425_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2849_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2703_ _3044_/Q _3348_/Q _3092_/Q _3068_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2703_/X sky130_fd_sc_hd__mux4_2
X_2634_ _2634_/A0 _2634_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__mux2_1
X_2565_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__clkbuf_1
X_1516_ _1524_/A vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__buf_1
XFILLER_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2496_ _3395_/Q vssd1 vssd1 vccd1 vccd1 _2496_/Y sky130_fd_sc_hd__inv_2
XINSDIODE2_8 _2697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3117_ _3437_/CLK _3117_/D vssd1 vssd1 vccd1 vccd1 _3117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3048_ _3371_/CLK _3048_/D vssd1 vssd1 vccd1 vccd1 _3048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3518_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2350_ _3052_/Q _2343_/X _2324_/X _2345_/X vssd1 vssd1 vccd1 vccd1 _3052_/D sky130_fd_sc_hd__a22o_1
X_2281_ _3095_/Q _2275_/X _2244_/X _2276_/X vssd1 vssd1 vccd1 vccd1 _3095_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _2011_/A vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__clkbuf_2
X_2617_ _2531_/X _2817_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2617_/X sky130_fd_sc_hd__mux2_1
X_2548_ _2548_/A _2552_/B vssd1 vssd1 vccd1 vccd1 _2548_/Y sky130_fd_sc_hd__nor2_1
X_2479_ _2479_/A _2479_/B vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__and2_1
XFILLER_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1850_ _1864_/A vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__inv_2
X_1781_ _1816_/A _2551_/A vssd1 vssd1 vccd1 vccd1 _2063_/A sky130_fd_sc_hd__or2_4
X_3451_ _3519_/CLK _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfxtp_1
X_3382_ _3424_/CLK _3382_/D vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfxtp_1
X_2402_ _3012_/Q _2397_/X _1939_/A _2398_/X vssd1 vssd1 vccd1 vccd1 _3012_/D sky130_fd_sc_hd__a22o_1
X_2333_ _3061_/Q _2326_/X _2332_/X _2328_/X vssd1 vssd1 vccd1 vccd1 _3061_/D sky130_fd_sc_hd__a22o_1
X_2264_ _3106_/Q _2257_/A _2247_/X _2258_/A vssd1 vssd1 vccd1 vccd1 _3106_/D sky130_fd_sc_hd__a22o_1
X_2195_ _3151_/Q _2191_/X _2158_/X _2193_/X vssd1 vssd1 vccd1 vccd1 _3151_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1979_ _3286_/Q _1977_/X _1944_/X _1978_/X vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2951_ _3188_/Q _3436_/Q _3140_/Q _3116_/Q _1676_/A _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2951_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1902_ _3327_/Q _1898_/X _1634_/X _1900_/X vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2882_ _3182_/Q _3158_/Q _3134_/Q _3110_/Q _2644_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2882_/X sky130_fd_sc_hd__mux4_2
X_1833_ _3371_/Q _1829_/X _1645_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__a22o_1
X_1764_ _3400_/Q _1761_/X _1722_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3503_ _3504_/CLK _3503_/D vssd1 vssd1 vccd1 vccd1 _3503_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _2258_/A vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__clkbuf_2
X_3434_ _3437_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
X_3365_ _3372_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
X_3296_ _3296_/CLK _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
X_2316_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2316_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2247_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2247_/X sky130_fd_sc_hd__buf_2
Xrepeater376 _2750_/S0 vssd1 vssd1 vccd1 vccd1 _2751_/S0 sky130_fd_sc_hd__buf_12
Xrepeater387 _2992_/S0 vssd1 vssd1 vccd1 vccd1 _2901_/S0 sky130_fd_sc_hd__buf_4
X_2178_ _3162_/Q _2172_/X _2130_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__a22o_1
Xrepeater398 _1700_/A vssd1 vssd1 vccd1 vccd1 _2991_/S0 sky130_fd_sc_hd__buf_8
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput102 io_b_dat_o_4[3] vssd1 vssd1 vccd1 vccd1 _2960_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput135 io_b_dat_o_6[4] vssd1 vssd1 vccd1 vccd1 _2947_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput113 io_b_dat_o_5[13] vssd1 vssd1 vccd1 vccd1 _2860_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput124 io_b_dat_o_5[9] vssd1 vssd1 vccd1 vccd1 _2887_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput146 io_b_dat_o_7[14] vssd1 vssd1 vccd1 vccd1 _2857_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput168 io_b_dat_o_8[5] vssd1 vssd1 vccd1 vccd1 _2600_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput157 io_b_dat_o_8[0] vssd1 vssd1 vccd1 vccd1 _2610_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput179 io_b_dat_o_9[15] vssd1 vssd1 vccd1 vccd1 _2576_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _3517_/Q vssd1 vssd1 vccd1 vccd1 _1482_/A sky130_fd_sc_hd__inv_2
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3150_ _3506_/CLK _3150_/D vssd1 vssd1 vccd1 vccd1 _3150_/Q sky130_fd_sc_hd__dfxtp_1
X_2101_ _3205_/Q _2097_/X _2046_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__a22o_1
X_3081_ _3273_/CLK _3081_/D vssd1 vssd1 vccd1 vccd1 _3081_/Q sky130_fd_sc_hd__dfxtp_1
X_2032_ _2052_/A vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__inv_2
XFILLER_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2934_ _2934_/A0 _2934_/A1 _2934_/A2 _2934_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2934_/X sky130_fd_sc_hd__mux4_1
X_2865_ _3064_/Q _3256_/Q _3232_/Q _3208_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2865_/X sky130_fd_sc_hd__mux4_2
X_1816_ _1816_/A _2552_/A vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__or2_4
X_2796_ _3024_/Q _3016_/Q _3008_/Q _3280_/Q _2851_/S0 _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2796_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1747_ _3408_/Q _1744_/X _1722_/X _1746_/X vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__a22o_1
X_1678_ _2540_/A _1678_/B _1678_/C _1678_/D vssd1 vssd1 vccd1 vccd1 _1798_/D sky130_fd_sc_hd__or4_4
X_3417_ _3423_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
X_3348_ _3392_/CLK _3348_/D vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3279_ _3279_/CLK _3279_/D vssd1 vssd1 vccd1 vccd1 _3279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A0 _2650_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2650_/X sky130_fd_sc_hd__mux2_1
X_1601_ _1603_/A _2909_/X vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__and2_1
X_2581_ _2581_/A0 _2581_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__mux2_1
X_1532_ _1515_/A _3503_/Q _1524_/A _2692_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _3503_/D
+ sky130_fd_sc_hd__o221a_1
X_3202_ _3372_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_1
X_3133_ _3180_/CLK _3133_/D vssd1 vssd1 vccd1 vccd1 _3133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3064_ _3398_/CLK _3064_/D vssd1 vssd1 vccd1 vccd1 _3064_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2015_ _3260_/Q _2011_/X _1949_/X _2012_/X vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2917_ _3083_/Q _3367_/Q _3035_/Q _3027_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2917_/X sky130_fd_sc_hd__mux4_1
X_2848_ _3417_/Q _3373_/Q _3389_/Q _3385_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2848_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2779_ _3291_/Q _3267_/Q _3243_/Q _3219_/Q _2682_/S _2911_/S1 vssd1 vssd1 vccd1 vccd1
+ _2779_/X sky130_fd_sc_hd__mux4_2
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2702_ _2698_/X _2699_/X _2700_/X _2701_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2702_/X sky130_fd_sc_hd__mux4_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2633_ _2633_/A0 _2633_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__mux2_1
X_2564_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__clkbuf_1
X_1515_ _1515_/A vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__buf_1
X_2495_ _3431_/Q vssd1 vssd1 vccd1 vccd1 _2495_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_9 _2707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3116_ _3333_/CLK _3116_/D vssd1 vssd1 vccd1 vccd1 _3116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3047_ _3351_/CLK _3047_/D vssd1 vssd1 vccd1 vccd1 _3047_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_57_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3297_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2280_ _3096_/Q _2275_/X _2242_/X _2276_/X vssd1 vssd1 vccd1 vccd1 _3096_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1995_ _1995_/A _2548_/A vssd1 vssd1 vccd1 vccd1 _2011_/A sky130_fd_sc_hd__or2_4
X_2616_ _2533_/X _2812_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2616_/X sky130_fd_sc_hd__mux2_1
X_2547_ _2553_/B vssd1 vssd1 vccd1 vccd1 _2552_/B sky130_fd_sc_hd__buf_1
X_2478_ _3427_/Q vssd1 vssd1 vccd1 vccd1 _2478_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _1815_/A _1780_/B _2342_/C vssd1 vssd1 vccd1 vccd1 _2551_/A sky130_fd_sc_hd__or3_4
X_3450_ _3519_/CLK _3450_/D vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2401_ _3013_/Q _2397_/X _2046_/A _2398_/X vssd1 vssd1 vccd1 vccd1 _3013_/D sky130_fd_sc_hd__a22o_1
X_3381_ _3409_/CLK _3381_/D vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2332_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2263_ _3107_/Q _2257_/X _2244_/X _2258_/X vssd1 vssd1 vccd1 vccd1 _3107_/D sky130_fd_sc_hd__a22o_1
X_2194_ _3152_/Q _2191_/X _2154_/X _2193_/X vssd1 vssd1 vccd1 vccd1 _3152_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1978_ _1978_/A vssd1 vssd1 vccd1 vccd1 _1978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_2_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3392_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2950_ _3284_/Q _3260_/Q _3236_/Q _3212_/Q _1700_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2950_/X sky130_fd_sc_hd__mux4_2
X_1901_ _3328_/Q _1898_/X _1630_/X _1900_/X vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__a22o_1
X_2881_ _3062_/Q _3254_/Q _3230_/Q _3206_/Q _2682_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2881_/X sky130_fd_sc_hd__mux4_2
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ _3372_/Q _1829_/X _1641_/X _1831_/X vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1763_ _2368_/A vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__clkbuf_2
X_1694_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2258_/A sky130_fd_sc_hd__inv_2
X_3502_ _3502_/CLK _3502_/D vssd1 vssd1 vccd1 vccd1 _3502_/Q sky130_fd_sc_hd__dfxtp_2
X_3433_ _3433_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
X_3364_ _3420_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
X_3295_ _3295_/CLK _3295_/D vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dfxtp_1
X_2315_ _3071_/Q _2309_/X _2244_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _3071_/D sky130_fd_sc_hd__a22o_1
X_2246_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2246_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater377 _2716_/S0 vssd1 vssd1 vccd1 vccd1 _2750_/S0 sky130_fd_sc_hd__buf_12
XFILLER_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2177_ _3163_/Q _2172_/X _2128_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__a22o_1
Xrepeater388 input7/X vssd1 vssd1 vccd1 vccd1 _2992_/S0 sky130_fd_sc_hd__clkbuf_8
Xrepeater399 _2996_/S0 vssd1 vssd1 vccd1 vccd1 _2982_/S0 sky130_fd_sc_hd__buf_8
XFILLER_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 io_b_dat_o_4[4] vssd1 vssd1 vccd1 vccd1 _2947_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput114 io_b_dat_o_5[14] vssd1 vssd1 vccd1 vccd1 _2857_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput136 io_b_dat_o_6[5] vssd1 vssd1 vccd1 vccd1 _2934_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput125 io_b_dat_o_6[0] vssd1 vssd1 vccd1 vccd1 _2999_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput147 io_b_dat_o_7[15] vssd1 vssd1 vccd1 vccd1 _2854_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput158 io_b_dat_o_8[10] vssd1 vssd1 vccd1 vccd1 _2590_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput169 io_b_dat_o_8[6] vssd1 vssd1 vccd1 vccd1 _2598_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _3448_/CLK _3080_/D vssd1 vssd1 vccd1 vccd1 _3080_/Q sky130_fd_sc_hd__dfxtp_1
X_2100_ _3206_/Q _2097_/X _2044_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__a22o_1
X_2031_ _2052_/A vssd1 vssd1 vccd1 vccd1 _2031_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2933_ input24/X input56/X input72/X input88/X _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2933_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2864_ _2490_/X _2492_/X _2640_/X _2494_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2864_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1815_ _1815_/A input8/X _2300_/C vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__or3_4
X_2795_ _3088_/Q _3372_/Q _3040_/Q _3032_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2795_/X sky130_fd_sc_hd__mux4_2
X_1746_ _2388_/A vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__clkbuf_2
X_1677_ _1846_/A _1780_/B _2342_/C vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__or3_4
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3416_ _3500_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3347_ _3392_/CLK _3347_/D vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3278_ _3279_/CLK _3278_/D vssd1 vssd1 vccd1 vccd1 _3278_/Q sky130_fd_sc_hd__dfxtp_1
X_2229_ _3127_/Q _2225_/X _2158_/X _2227_/X vssd1 vssd1 vccd1 vccd1 _3127_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1600_ _1603_/A _2896_/X vssd1 vssd1 vccd1 vccd1 _3465_/D sky130_fd_sc_hd__and2_1
X_2580_ _2579_/X _2511_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__mux2_1
X_1531_ _1515_/A _3504_/Q _1524_/A _2697_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _3504_/D
+ sky130_fd_sc_hd__o221a_1
X_3201_ _3372_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_1
X_3132_ _3180_/CLK _3132_/D vssd1 vssd1 vccd1 vccd1 _3132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3063_ _3279_/CLK _3063_/D vssd1 vssd1 vccd1 vccd1 _3063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2014_ _3261_/Q _2011_/X _1947_/X _2012_/X vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2916_ _3179_/Q _3155_/Q _3131_/Q _3107_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2916_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2847_ _2843_/X _2844_/X _2845_/X _2846_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2847_/X sky130_fd_sc_hd__mux4_2
X_2778_ _3171_/Q _3339_/Q _3323_/Q _3307_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2778_/X sky130_fd_sc_hd__mux4_2
X_1729_ _3414_/Q _1721_/X _1728_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2701_ _3315_/Q _3299_/Q _3163_/Q _3331_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2701_/X sky130_fd_sc_hd__mux4_1
X_2632_ _2632_/A0 _2632_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2632_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2563_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__clkbuf_1
X_1514_ _3515_/Q _1515_/A _2752_/X _1524_/A _1510_/X vssd1 vssd1 vccd1 vccd1 _3515_/D
+ sky130_fd_sc_hd__o221a_1
X_2494_ _2523_/A _2586_/X vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__and2_1
XFILLER_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3115_ _3346_/CLK _3115_/D vssd1 vssd1 vccd1 vccd1 _3115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3046_ _3350_/CLK _3046_/D vssd1 vssd1 vccd1 vccd1 _3046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3497_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1994_ _3273_/Q _1986_/A _1947_/X _1987_/A vssd1 vssd1 vccd1 vccd1 _3273_/D sky130_fd_sc_hd__a22o_1
X_2615_ _2535_/X _2807_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__mux2_1
X_2546_ _2546_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__nor2_1
X_2477_ _3387_/Q vssd1 vssd1 vccd1 vccd1 _2477_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3029_ _3371_/CLK _3029_/D vssd1 vssd1 vccd1 vccd1 _3029_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2400_ _3014_/Q _2397_/X _2044_/A _2398_/X vssd1 vssd1 vccd1 vccd1 _3014_/D sky130_fd_sc_hd__a22o_1
X_3380_ _3429_/CLK _3380_/D vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfxtp_1
X_2331_ _3062_/Q _2326_/X _2330_/X _2328_/X vssd1 vssd1 vccd1 vccd1 _3062_/D sky130_fd_sc_hd__a22o_1
X_2262_ _3108_/Q _2257_/X _2242_/X _2258_/X vssd1 vssd1 vccd1 vccd1 _3108_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2193_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2193_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1977_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1977_/X sky130_fd_sc_hd__clkbuf_2
X_2529_ _3449_/Q _3450_/Q _2526_/B vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__a21bo_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2880_ _2475_/X _2645_/X _2646_/X _2480_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2880_/X sky130_fd_sc_hd__mux4_2
X_1900_ _1914_/A vssd1 vssd1 vccd1 vccd1 _1900_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1831_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1831_/X sky130_fd_sc_hd__buf_2
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1762_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2368_/A sky130_fd_sc_hd__inv_2
X_3501_ _3501_/CLK _3501_/D vssd1 vssd1 vccd1 vccd1 _3501_/Q sky130_fd_sc_hd__dfxtp_1
X_1693_ _2257_/A vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__clkbuf_2
X_3432_ _3493_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3515_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3363_ _3420_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
X_3294_ _3294_/CLK _3294_/D vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfxtp_1
X_2314_ _3072_/Q _2309_/X _2242_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _3072_/D sky130_fd_sc_hd__a22o_1
X_2245_ _3119_/Q _2234_/X _2244_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _3119_/D sky130_fd_sc_hd__a22o_1
Xrepeater378 _2710_/S0 vssd1 vssd1 vccd1 vccd1 _2716_/S0 sky130_fd_sc_hd__buf_6
X_2176_ _3164_/Q _2172_/X _2126_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater389 _2911_/S1 vssd1 vssd1 vccd1 vccd1 _2913_/S1 sky130_fd_sc_hd__buf_6
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput126 io_b_dat_o_6[10] vssd1 vssd1 vccd1 vccd1 _2879_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput115 io_b_dat_o_5[15] vssd1 vssd1 vccd1 vccd1 _2854_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput104 io_b_dat_o_4[5] vssd1 vssd1 vccd1 vccd1 _2934_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput159 io_b_dat_o_8[11] vssd1 vssd1 vccd1 vccd1 _2588_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput148 io_b_dat_o_7[1] vssd1 vssd1 vccd1 vccd1 _2986_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput137 io_b_dat_o_6[6] vssd1 vssd1 vccd1 vccd1 _2921_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2030_ _2190_/A _2546_/A vssd1 vssd1 vccd1 vccd1 _2052_/A sky130_fd_sc_hd__or2_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2932_ _2928_/X _2929_/X _2930_/X _2931_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2932_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2863_ input96/X _2863_/A1 _2863_/A2 _2863_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2863_/X sky130_fd_sc_hd__mux4_1
X_1814_ _3377_/Q _1808_/X _1778_/X _1810_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__a22o_1
X_2794_ _3184_/Q _3160_/Q _3136_/Q _3112_/Q _2851_/S0 _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2794_/X sky130_fd_sc_hd__mux4_1
XFILLER_7_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1745_ _2387_/A vssd1 vssd1 vccd1 vccd1 _2388_/A sky130_fd_sc_hd__inv_2
X_1676_ _1676_/A _1689_/B vssd1 vssd1 vccd1 vccd1 _2342_/C sky130_fd_sc_hd__or2_2
X_3415_ _3482_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3346_/CLK _3346_/D vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3277_ _3277_/CLK _3277_/D vssd1 vssd1 vccd1 vccd1 _3277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2228_ _3128_/Q _2225_/X _2154_/X _2227_/X vssd1 vssd1 vccd1 vccd1 _3128_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _3175_/Q _2153_/X _2158_/X _2156_/X vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1530_ _1523_/X _3505_/Q _1524_/X _2702_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _3505_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200_ _3294_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_1
X_3131_ _3497_/CLK _3131_/D vssd1 vssd1 vccd1 vccd1 _3131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3062_ _3279_/CLK _3062_/D vssd1 vssd1 vccd1 vccd1 _3062_/Q sky130_fd_sc_hd__dfxtp_1
X_2013_ _3262_/Q _2011_/X _1944_/X _2012_/X vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2915_ _3059_/Q _3251_/Q _3227_/Q _3203_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2915_/X sky130_fd_sc_hd__mux4_2
X_2846_ _2452_/Y _2471_/Y _2474_/Y _2453_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2846_/X sky130_fd_sc_hd__mux4_1
X_2777_ _2773_/X _2774_/X _2775_/X _2776_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2777_/X sky130_fd_sc_hd__mux4_2
X_1728_ _1728_/A vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__clkbuf_2
X_1659_ _1944_/A vssd1 vssd1 vccd1 vccd1 _1659_/X sky130_fd_sc_hd__buf_2
X_3329_ _3433_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ _3235_/Q _3211_/Q _3283_/Q _3259_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2700_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2631_ _2631_/A0 _2631_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2631_/X sky130_fd_sc_hd__mux2_1
X_2562_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2562_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1513_ _1513_/A vssd1 vssd1 vccd1 vccd1 _1524_/A sky130_fd_sc_hd__clkbuf_2
X_2493_ _2522_/A _2493_/B vssd1 vssd1 vccd1 vccd1 _2493_/X sky130_fd_sc_hd__and2_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3114_ _3346_/CLK _3114_/D vssd1 vssd1 vccd1 vccd1 _3114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3045_ _3350_/CLK _3045_/D vssd1 vssd1 vccd1 vccd1 _3045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2829_ _3177_/Q _3153_/Q _3129_/Q _3105_/Q _2851_/S0 _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2829_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _3274_/Q _1986_/A _1944_/X _1987_/A vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__a22o_1
X_2614_ _2538_/Y _2802_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2614_/X sky130_fd_sc_hd__mux2_1
X_2545_ _2545_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2545_/Y sky130_fd_sc_hd__nor2_1
X_2476_ _3411_/Q vssd1 vssd1 vccd1 vccd1 _2476_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _3371_/CLK _3028_/D vssd1 vssd1 vccd1 vccd1 _3028_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2330_/X sky130_fd_sc_hd__clkbuf_2
X_2261_ _3109_/Q _2257_/X _2240_/X _2258_/X vssd1 vssd1 vccd1 vccd1 _3109_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2192_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2207_/A sky130_fd_sc_hd__inv_2
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1976_ _3287_/Q _1970_/X _1941_/X _1971_/X vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2528_ _2528_/A _2532_/B vssd1 vssd1 vccd1 vccd1 _2620_/S sky130_fd_sc_hd__nor2_8
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2459_ _2458_/Y _2459_/A2 _1557_/X _2459_/B2 _3496_/Q vssd1 vssd1 vccd1 vccd1 _2459_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _1837_/A vssd1 vssd1 vccd1 vccd1 _1838_/A sky130_fd_sc_hd__inv_2
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ _3500_/CLK _3500_/D vssd1 vssd1 vccd1 vccd1 _3500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1761_ _2367_/A vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__clkbuf_2
X_1692_ _1760_/A _2545_/A vssd1 vssd1 vccd1 vccd1 _2257_/A sky130_fd_sc_hd__or2_4
X_3431_ _3493_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
X_3362_ _3398_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
X_2313_ _3073_/Q _2309_/X _2240_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _3073_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3293_ _3294_/CLK _3293_/D vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2244_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__clkbuf_2
X_2175_ _3165_/Q _2172_/X _2150_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3423_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xrepeater379 _2852_/X vssd1 vssd1 vccd1 vccd1 _2710_/S0 sky130_fd_sc_hd__buf_8
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1959_ _2573_/A vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput105 io_b_dat_o_4[6] vssd1 vssd1 vccd1 vccd1 _2921_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput127 io_b_dat_o_6[11] vssd1 vssd1 vccd1 vccd1 _2871_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput116 io_b_dat_o_5[1] vssd1 vssd1 vccd1 vccd1 _2986_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput149 io_b_dat_o_7[2] vssd1 vssd1 vccd1 vccd1 _2973_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput138 io_b_dat_o_6[7] vssd1 vssd1 vccd1 vccd1 _2908_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2931_ _3018_/Q _3010_/Q _3002_/Q _3274_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2931_/X sky130_fd_sc_hd__mux4_1
X_2862_ input16/X input48/X input64/X input80/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2862_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1813_ _3378_/Q _1808_/X _1776_/X _1810_/X vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__a22o_1
X_2793_ _3064_/Q _3256_/Q _3232_/Q _3208_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2793_/X sky130_fd_sc_hd__mux4_2
X_1744_ _2387_/A vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3414_ _3500_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
X_1675_ _2611_/S vssd1 vssd1 vccd1 vccd1 _1689_/B sky130_fd_sc_hd__inv_2
X_3345_ _3502_/CLK _3345_/D vssd1 vssd1 vccd1 vccd1 _3345_/Q sky130_fd_sc_hd__dfxtp_1
X_3276_ _3279_/CLK _3276_/D vssd1 vssd1 vccd1 vccd1 _3276_/Q sky130_fd_sc_hd__dfxtp_1
X_2227_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2227_/X sky130_fd_sc_hd__buf_2
X_2158_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2089_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3130_ _3497_/CLK _3130_/D vssd1 vssd1 vccd1 vccd1 _3130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3061_ _3353_/CLK _3061_/D vssd1 vssd1 vccd1 vccd1 _3061_/Q sky130_fd_sc_hd__dfxtp_1
X_2012_ _2012_/A vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__buf_2
XFILLER_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2914_ _2910_/X _2911_/X _2912_/X _2913_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2914_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2845_ _2443_/Y _2457_/Y _2454_/Y _2468_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2845_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2776_ _3100_/Q _3076_/Q _3052_/Q _3356_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2776_/X sky130_fd_sc_hd__mux4_2
X_1727_ _3415_/Q _1721_/X _1726_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__a22o_1
X_1658_ _1658_/A vssd1 vssd1 vccd1 vccd1 _1658_/X sky130_fd_sc_hd__clkbuf_2
X_3328_ _3344_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
X_1589_ _3474_/Q vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__inv_2
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _3474_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _2630_/A0 _2630_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2630_/X sky130_fd_sc_hd__mux2_2
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2561_ _2561_/A vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__buf_1
X_2492_ _2509_/A _2587_/X vssd1 vssd1 vccd1 vccd1 _2492_/X sky130_fd_sc_hd__and2_1
X_1512_ _3502_/Q vssd1 vssd1 vccd1 vccd1 _1515_/A sky130_fd_sc_hd__buf_2
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _3433_/CLK _3113_/D vssd1 vssd1 vccd1 vccd1 _3113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3044_ _3392_/CLK _3044_/D vssd1 vssd1 vccd1 vccd1 _3044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2828_ _3057_/Q _3249_/Q _3225_/Q _3201_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2828_/X sky130_fd_sc_hd__mux4_2
X_2759_ _3295_/Q _3271_/Q _3247_/Q _3223_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2759_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1992_ _3275_/Q _1986_/X _1941_/X _1987_/X vssd1 vssd1 vccd1 vccd1 _3275_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_35_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3351_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2613_ _2539_/X _2797_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2613_/X sky130_fd_sc_hd__mux2_1
X_2544_ _2544_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2475_ _2490_/A _2782_/X vssd1 vssd1 vccd1 vccd1 _2475_/X sky130_fd_sc_hd__and2_1
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3027_ _3275_/CLK _3027_/D vssd1 vssd1 vccd1 vccd1 _3027_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2260_ _3110_/Q _2257_/X _2238_/X _2258_/X vssd1 vssd1 vccd1 vccd1 _3110_/D sky130_fd_sc_hd__a22o_1
X_2191_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2191_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _3288_/Q _1970_/X _1939_/X _1971_/X vssd1 vssd1 vccd1 vccd1 _3288_/D sky130_fd_sc_hd__a22o_1
X_2527_ _3452_/Q _2527_/B vssd1 vssd1 vccd1 vccd1 _2532_/B sky130_fd_sc_hd__or2_4
X_2458_ _3495_/Q vssd1 vssd1 vccd1 vccd1 _2458_/Y sky130_fd_sc_hd__inv_2
X_2389_ _3023_/Q _2387_/X _2327_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _3023_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1760_ _1760_/A _2542_/A vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__or2_4
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1691_ _1806_/A _1780_/B _2224_/C vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__or3_4
X_3430_ _3500_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
X_3361_ _3398_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2312_ _3074_/Q _2309_/X _2238_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _3074_/D sky130_fd_sc_hd__a22o_1
X_3292_ _3297_/CLK _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2243_ _3120_/Q _2234_/X _2242_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _3120_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2174_ _3166_/Q _2172_/X _2148_/X _2173_/X vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1958_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1958_/X sky130_fd_sc_hd__clkbuf_2
X_1889_ _1889_/A vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput117 io_b_dat_o_5[2] vssd1 vssd1 vccd1 vccd1 _2973_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput106 io_b_dat_o_4[7] vssd1 vssd1 vccd1 vccd1 _2908_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput128 io_b_dat_o_6[12] vssd1 vssd1 vccd1 vccd1 _2863_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput139 io_b_dat_o_6[8] vssd1 vssd1 vccd1 vccd1 _2895_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2930_ _3082_/Q _3366_/Q _3034_/Q _3026_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2930_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2497_/X _2498_/X _2639_/X _2500_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2861_/X sky130_fd_sc_hd__mux4_2
X_1812_ _3379_/Q _1808_/X _1774_/X _1810_/X vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2792_ _2788_/X _2789_/X _2790_/X _2791_/X _2901_/S0 _2997_/S1 vssd1 vssd1 vccd1
+ vccd1 _2792_/X sky130_fd_sc_hd__mux4_2
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1743_ _2342_/A _1798_/B _2266_/C _1828_/B vssd1 vssd1 vccd1 vccd1 _2387_/A sky130_fd_sc_hd__or4_4
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1674_ input8/X vssd1 vssd1 vccd1 vccd1 _1780_/B sky130_fd_sc_hd__buf_1
X_3413_ _3429_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3344_/CLK _3344_/D vssd1 vssd1 vccd1 vccd1 _3344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3275_ _3275_/CLK _3275_/D vssd1 vssd1 vccd1 vccd1 _3275_/Q sky130_fd_sc_hd__dfxtp_1
X_2226_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2248_/A sky130_fd_sc_hd__inv_2
X_2157_ _3176_/Q _2153_/X _2154_/X _2156_/X vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2088_ _2088_/A vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3060_ _3279_/CLK _3060_/D vssd1 vssd1 vccd1 vccd1 _3060_/Q sky130_fd_sc_hd__dfxtp_1
X_2011_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2011_/X sky130_fd_sc_hd__buf_2
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2913_ _3095_/Q _3071_/Q _3047_/Q _3351_/Q _2913_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2913_/X sky130_fd_sc_hd__mux4_1
X_2844_ _2442_/Y _2440_/Y _2445_/Y _2444_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2844_/X sky130_fd_sc_hd__mux4_2
X_2775_ _3196_/Q _3444_/Q _3148_/Q _3124_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2775_/X sky130_fd_sc_hd__mux4_1
X_1726_ _1726_/A vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__clkbuf_2
X_1657_ _3439_/Q _1643_/X _1656_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__a22o_1
X_1588_ _1590_/A _2540_/A vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3327_ _3344_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
X_3258_ _3331_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2209_ _3141_/Q _2206_/X _2150_/X _2207_/X vssd1 vssd1 vccd1 vccd1 _3141_/D sky130_fd_sc_hd__a22o_1
X_3189_ _3437_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__buf_1
X_1511_ _2687_/S _1508_/Y _3516_/Q _1502_/Y _1510_/X vssd1 vssd1 vccd1 vccd1 _3516_/D
+ sky130_fd_sc_hd__o221a_1
X_2491_ _2520_/A vssd1 vssd1 vccd1 vccd1 _2509_/A sky130_fd_sc_hd__buf_1
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _3501_/CLK _3112_/D vssd1 vssd1 vccd1 vccd1 _3112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3043_ _3392_/CLK _3043_/D vssd1 vssd1 vccd1 vccd1 _3043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2827_ _2823_/X _2824_/X _2825_/X _2826_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2827_/X sky130_fd_sc_hd__mux4_2
X_2758_ _3175_/Q _3343_/Q _3327_/Q _3311_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2758_/X sky130_fd_sc_hd__mux4_2
X_1709_ _3421_/Q _1703_/X _1670_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__a22o_1
X_2689_ _3137_/Q _3113_/Q _3185_/Q _3433_/Q _2716_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2689_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3350_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1991_ _3276_/Q _1986_/X _1939_/X _1987_/X vssd1 vssd1 vccd1 vccd1 _3276_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2612_ _1506_/X _3517_/Q _2687_/S vssd1 vssd1 vccd1 vccd1 _2612_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2543_ _2543_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2543_/Y sky130_fd_sc_hd__nor2_1
X_2474_ _3410_/Q vssd1 vssd1 vccd1 vccd1 _2474_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3026_ _3367_/CLK _3026_/D vssd1 vssd1 vccd1 vccd1 _3026_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2190_ _2190_/A _2542_/A vssd1 vssd1 vccd1 vccd1 _2206_/A sky130_fd_sc_hd__or2_4
XFILLER_1_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _3289_/Q _1970_/X _1937_/X _1971_/X vssd1 vssd1 vccd1 vccd1 _3289_/D sky130_fd_sc_hd__a22o_1
X_2526_ _3451_/Q _2526_/B vssd1 vssd1 vccd1 vccd1 _2527_/B sky130_fd_sc_hd__or2_1
X_2457_ _3362_/Q vssd1 vssd1 vccd1 vccd1 _2457_/Y sky130_fd_sc_hd__inv_2
X_2388_ _2388_/A vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ _3273_/CLK _3009_/D vssd1 vssd1 vccd1 vccd1 _3009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1690_ _1789_/C vssd1 vssd1 vccd1 vccd1 _2224_/C sky130_fd_sc_hd__clkbuf_2
X_3360_ _3448_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_1
X_2311_ _3075_/Q _2309_/X _2235_/X _2310_/X vssd1 vssd1 vccd1 vccd1 _3075_/D sky130_fd_sc_hd__a22o_1
X_3291_ _3303_/CLK _3291_/D vssd1 vssd1 vccd1 vccd1 _3291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2242_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2173_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2173_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1957_ _1995_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__or2_4
X_1888_ _3335_/Q _1882_/X _1656_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__a22o_1
X_2509_ _2509_/A _2581_/X vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__and2_1
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput118 io_b_dat_o_5[3] vssd1 vssd1 vccd1 vccd1 _2960_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput107 io_b_dat_o_4[8] vssd1 vssd1 vccd1 vccd1 _2895_/A0 sky130_fd_sc_hd__clkbuf_1
X_3489_ _3518_/CLK _3489_/D vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfxtp_1
Xinput129 io_b_dat_o_6[13] vssd1 vssd1 vccd1 vccd1 _2860_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2860_ input97/X _2860_/A1 _2860_/A2 _2860_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2860_/X sky130_fd_sc_hd__mux4_1
X_1811_ _3380_/Q _1808_/X _1770_/X _1810_/X vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__a22o_1
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ _3097_/Q _3073_/Q _3049_/Q _3353_/Q _2913_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2791_/X sky130_fd_sc_hd__mux4_2
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1742_ _3409_/Q _1736_/X _1730_/X _1738_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1673_ _1806_/A vssd1 vssd1 vccd1 vccd1 _1846_/A sky130_fd_sc_hd__buf_1
X_3412_ _3429_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_1
X_3343_ _3344_/CLK _3343_/D vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfxtp_1
X_3274_ _3275_/CLK _3274_/D vssd1 vssd1 vccd1 vccd1 _3274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2225_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__buf_2
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2156_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2156_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2087_ _3215_/Q _2081_/X _2050_/X _2082_/X vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2989_ _3281_/Q _3257_/Q _3233_/Q _3209_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2989_/X sky130_fd_sc_hd__mux4_2
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _3263_/Q _2004_/X _1941_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_29_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2912_ _3191_/Q _3439_/Q _3143_/Q _3119_/Q _2913_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2912_/X sky130_fd_sc_hd__mux4_1
X_2843_ _2433_/Y _2432_/Y _2431_/Y _2428_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2843_/X sky130_fd_sc_hd__mux4_2
X_2774_ _3292_/Q _3268_/Q _3244_/Q _3220_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2774_/X sky130_fd_sc_hd__mux4_2
X_1725_ _3416_/Q _1721_/X _1722_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__a22o_1
X_1656_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__clkbuf_2
X_1587_ _1591_/A _2687_/X vssd1 vssd1 vccd1 vccd1 _3475_/D sky130_fd_sc_hd__and2_1
X_3326_ _3509_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3257_ _3297_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3188_ _3333_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_1
X_2208_ _3142_/Q _2206_/X _2148_/X _2207_/X vssd1 vssd1 vccd1 vccd1 _3142_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2139_ _3183_/Q _2136_/X _2137_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1510_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1510_/X sky130_fd_sc_hd__clkbuf_4
X_2490_ _2490_/A _2772_/X vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__and2_1
XFILLER_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3111_ _3180_/CLK _3111_/D vssd1 vssd1 vccd1 vccd1 _3111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput290 io_dsi_in[4] vssd1 vssd1 vccd1 vccd1 _2463_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_67_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3042_ _3346_/CLK _3042_/D vssd1 vssd1 vccd1 vccd1 _3042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2826_ _3018_/Q _3010_/Q _3002_/Q _3274_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2826_/X sky130_fd_sc_hd__mux4_1
X_2757_ _2753_/X _2754_/X _2755_/X _2756_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2757_/X sky130_fd_sc_hd__mux4_2
X_2688_ _3041_/Q _3345_/Q _3089_/Q _3065_/Q _2716_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2688_/X sky130_fd_sc_hd__mux4_2
X_1708_ _3422_/Q _1703_/X _1668_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__a22o_1
X_1639_ _3445_/Q _1629_/X _1638_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__a22o_1
XFILLER_86_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3309_ _3340_/CLK _3309_/D vssd1 vssd1 vccd1 vccd1 _3309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _3277_/Q _1986_/X _1937_/X _1987_/X vssd1 vssd1 vccd1 vccd1 _3277_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2611_ _2610_/X _2422_/X _2611_/S vssd1 vssd1 vccd1 vccd1 _2611_/X sky130_fd_sc_hd__mux2_1
X_2542_ _2542_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__nor2_1
X_2473_ _2480_/A _2593_/X vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__and2_1
XFILLER_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3509_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3025_ _3273_/CLK _3025_/D vssd1 vssd1 vccd1 vccd1 _3025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2809_ _3181_/Q _3157_/Q _3133_/Q _3109_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2809_/X sky130_fd_sc_hd__mux4_2
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1973_ _3290_/Q _1970_/X _1935_/X _1971_/X vssd1 vssd1 vccd1 vccd1 _3290_/D sky130_fd_sc_hd__a22o_1
X_2525_ _3449_/Q _3450_/Q vssd1 vssd1 vccd1 vccd1 _2526_/B sky130_fd_sc_hd__or2_1
X_2456_ _2480_/A _2595_/X vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__and2_1
XFILLER_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2387_ _2387_/A vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3008_ _3410_/CLK _3008_/D vssd1 vssd1 vccd1 vccd1 _3008_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3290_ _3515_/CLK _3290_/D vssd1 vssd1 vccd1 vccd1 _3290_/Q sky130_fd_sc_hd__dfxtp_1
X_2310_ _2317_/A vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__clkbuf_2
X_2241_ _3121_/Q _2234_/X _2240_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _3121_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2172_ _2172_/A vssd1 vssd1 vccd1 vccd1 _2172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1956_ _3297_/Q _1943_/A _1955_/X _1945_/A vssd1 vssd1 vccd1 vccd1 _3297_/D sky130_fd_sc_hd__a22o_1
X_1887_ _3336_/Q _1882_/X _1654_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__a22o_1
X_2508_ _2509_/A _2762_/X vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__and2_1
Xinput108 io_b_dat_o_4[9] vssd1 vssd1 vccd1 vccd1 _2887_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3488_ _3518_/CLK _3488_/D vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfxtp_1
Xinput119 io_b_dat_o_5[4] vssd1 vssd1 vccd1 vccd1 _2947_/A1 sky130_fd_sc_hd__clkbuf_1
X_2439_ _2480_/A _2599_/X vssd1 vssd1 vccd1 vccd1 _2439_/X sky130_fd_sc_hd__and2_1
XFILLER_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _2138_/A vssd1 vssd1 vccd1 vccd1 _1810_/X sky130_fd_sc_hd__clkbuf_2
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2790_ _3193_/Q _3441_/Q _3145_/Q _3121_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2790_/X sky130_fd_sc_hd__mux4_1
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1741_ _3410_/Q _1736_/X _1728_/X _1738_/X vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1672_ input7/X vssd1 vssd1 vccd1 vccd1 _1806_/A sky130_fd_sc_hd__inv_2
X_3411_ _3429_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3342_ _3344_/CLK _3342_/D vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfxtp_1
X_3273_ _3273_/CLK _3273_/D vssd1 vssd1 vccd1 vccd1 _3273_/Q sky130_fd_sc_hd__dfxtp_1
X_2224_ _2224_/A _2342_/B _2224_/C _2300_/D vssd1 vssd1 vccd1 vccd1 _2246_/A sky130_fd_sc_hd__or4_4
X_2155_ _2172_/A vssd1 vssd1 vccd1 vccd1 _2173_/A sky130_fd_sc_hd__inv_2
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ _3216_/Q _2081_/X _2048_/X _2082_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2988_ _3161_/Q _3329_/Q _3313_/Q _3297_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2988_/X sky130_fd_sc_hd__mux4_2
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ _1939_/A vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__clkbuf_2
Xinput90 io_b_dat_o_3[7] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2911_ _3287_/Q _3263_/Q _3239_/Q _3215_/Q _2682_/S _2911_/S1 vssd1 vssd1 vccd1 vccd1
+ _2911_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2842_ _2838_/X _2839_/X _2840_/X _2841_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2842_/X sky130_fd_sc_hd__mux4_2
X_2773_ _3172_/Q _3340_/Q _3324_/Q _3308_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2773_/X sky130_fd_sc_hd__mux4_2
X_1724_ _2182_/A vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__clkbuf_2
X_1655_ _3440_/Q _1643_/X _1654_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__a22o_1
X_1586_ _1591_/A _2612_/X vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__and2_1
X_3325_ _3509_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3256_ _3398_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
X_2207_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2207_/X sky130_fd_sc_hd__buf_2
X_3187_ _3333_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
X_2138_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2069_ _3227_/Q _2063_/X _2050_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3110_ _3180_/CLK _3110_/D vssd1 vssd1 vccd1 vccd1 _3110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput280 io_dataLastBlock[62] vssd1 vssd1 vccd1 vccd1 _2622_/A1 sky130_fd_sc_hd__clkbuf_1
X_3041_ _3502_/CLK _3041_/D vssd1 vssd1 vccd1 vccd1 _3041_/Q sky130_fd_sc_hd__dfxtp_1
Xinput291 io_dsi_in[5] vssd1 vssd1 vccd1 vccd1 _2463_/B2 sky130_fd_sc_hd__buf_2
XFILLER_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2825_ _3082_/Q _3366_/Q _3034_/Q _3026_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2825_/X sky130_fd_sc_hd__mux4_2
X_2756_ _3104_/Q _3080_/Q _3056_/Q _3360_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2756_/X sky130_fd_sc_hd__mux4_1
X_2687_ _1508_/Y _3516_/Q _2687_/S vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__mux2_1
X_1707_ _3423_/Q _1703_/X _1666_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__a22o_1
X_1638_ _2570_/A vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1569_ _1569_/A _2625_/X vssd1 vssd1 vccd1 vccd1 _3490_/D sky130_fd_sc_hd__nor2b_1
X_3308_ _3515_/CLK _3308_/D vssd1 vssd1 vccd1 vccd1 _3308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3239_ _3303_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2610_ _2610_/A0 _2610_/A1 _2610_/S vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__mux2_1
X_2541_ _2553_/B vssd1 vssd1 vccd1 vccd1 _2546_/B sky130_fd_sc_hd__buf_1
X_2472_ _2479_/A _2472_/B vssd1 vssd1 vccd1 vccd1 _2472_/X sky130_fd_sc_hd__and2_1
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3024_ _3410_/CLK _3024_/D vssd1 vssd1 vccd1 vccd1 _3024_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2808_ _3061_/Q _3253_/Q _3229_/Q _3205_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2808_/X sky130_fd_sc_hd__mux4_2
X_2739_ _3147_/Q _3123_/Q _3195_/Q _3443_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2739_/X sky130_fd_sc_hd__mux4_1
XFILLER_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1972_ _3291_/Q _1970_/X _1932_/X _1971_/X vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2524_ _3420_/Q vssd1 vssd1 vccd1 vccd1 _2524_/Y sky130_fd_sc_hd__inv_2
X_2455_ _2479_/A _2455_/B vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__and2_1
X_2386_ _3024_/Q _1744_/X _2324_/X _1746_/X vssd1 vssd1 vccd1 vccd1 _3024_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3007_ _3277_/CLK _3007_/D vssd1 vssd1 vccd1 vccd1 _3007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput370 _3510_/Q vssd1 vssd1 vccd1 vccd1 io_vout[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2240_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _3167_/Q _2165_/X _2146_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ _2558_/A vssd1 vssd1 vccd1 vccd1 _1955_/X sky130_fd_sc_hd__clkbuf_2
X_1886_ _3337_/Q _1882_/X _1652_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__a22o_1
X_2507_ _3399_/Q vssd1 vssd1 vccd1 vccd1 _2507_/Y sky130_fd_sc_hd__inv_2
Xinput109 io_b_dat_o_5[0] vssd1 vssd1 vccd1 vccd1 _2999_/A1 sky130_fd_sc_hd__clkbuf_1
X_3487_ _3518_/CLK _3487_/D vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfxtp_1
X_2438_ _2487_/A vssd1 vssd1 vccd1 vccd1 _2480_/A sky130_fd_sc_hd__buf_1
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2369_ _3039_/Q _2367_/X _2327_/X _2368_/X vssd1 vssd1 vccd1 vccd1 _3039_/D sky130_fd_sc_hd__a22o_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _3411_/Q _1736_/X _1726_/X _1738_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__a22o_1
X_1671_ _3433_/Q _1658_/A _1670_/X _1660_/A vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__a22o_1
X_3410_ _3410_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
X_3341_ _3509_/CLK _3341_/D vssd1 vssd1 vccd1 vccd1 _3341_/Q sky130_fd_sc_hd__dfxtp_1
X_3272_ _3301_/CLK _3272_/D vssd1 vssd1 vccd1 vccd1 _3272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2223_ _3129_/Q _2215_/A _2150_/X _2216_/A vssd1 vssd1 vccd1 vccd1 _3129_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2154_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _3217_/Q _2081_/X _2046_/X _2082_/X vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2987_ _2677_/X _2679_/X _2680_/X _2421_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2987_/X sky130_fd_sc_hd__mux4_1
X_1938_ _3305_/Q _1931_/X _1937_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _3305_/D sky130_fd_sc_hd__a22o_1
X_1869_ _3347_/Q _1864_/X _1822_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__a22o_1
Xinput80 io_b_dat_o_3[12] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_1
Xinput91 io_b_dat_o_3[8] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2910_ _3167_/Q _3335_/Q _3319_/Q _3303_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2910_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2841_ _2506_/Y _2484_/Y _2476_/Y _2449_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2841_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2772_ _2768_/X _2769_/X _2770_/X _2771_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2772_/X sky130_fd_sc_hd__mux4_2
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1723_ _2181_/A vssd1 vssd1 vccd1 vccd1 _2182_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_38_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3355_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1654_ _1939_/A vssd1 vssd1 vccd1 vccd1 _1654_/X sky130_fd_sc_hd__clkbuf_2
X_1585_ _1591_/A _2685_/X vssd1 vssd1 vccd1 vccd1 _3477_/D sky130_fd_sc_hd__and2_1
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3324_ _3515_/CLK _3324_/D vssd1 vssd1 vccd1 vccd1 _3324_/Q sky130_fd_sc_hd__dfxtp_1
X_3255_ _3279_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
X_2206_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3186_ _3346_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2137_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2137_/X sky130_fd_sc_hd__buf_2
X_2068_ _3228_/Q _2063_/X _2048_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _3228_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput281 io_dataLastBlock[63] vssd1 vssd1 vccd1 vccd1 _2621_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput270 io_dataLastBlock[53] vssd1 vssd1 vccd1 vccd1 _2631_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ _3398_/CLK _3040_/D vssd1 vssd1 vccd1 vccd1 _3040_/Q sky130_fd_sc_hd__dfxtp_1
Xinput292 io_dsi_in[6] vssd1 vssd1 vccd1 vccd1 _2464_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2824_ _3178_/Q _3154_/Q _3130_/Q _3106_/Q _2851_/S0 _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2824_/X sky130_fd_sc_hd__mux4_2
X_2755_ _3200_/Q _3448_/Q _3152_/Q _3128_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2755_/X sky130_fd_sc_hd__mux4_1
X_2686_ _1491_/X _3519_/Q _2687_/S vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__mux2_1
X_1706_ _3424_/Q _1703_/X _1664_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__a22o_1
X_1637_ _3446_/Q _1629_/X _1636_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__a22o_1
X_1568_ _1569_/A _2624_/X vssd1 vssd1 vccd1 vccd1 _3491_/D sky130_fd_sc_hd__nor2b_1
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3307_ _3307_/CLK _3307_/D vssd1 vssd1 vccd1 vccd1 _3307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1499_ _1513_/A _1499_/B vssd1 vssd1 vccd1 vccd1 _1502_/A sky130_fd_sc_hd__or2_2
X_3238_ _3296_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
X_3169_ _3335_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2540_ _2540_/A input3/X input2/X vssd1 vssd1 vccd1 vccd1 _2553_/B sky130_fd_sc_hd__or3b_4
X_2471_ _3402_/Q vssd1 vssd1 vccd1 vccd1 _2471_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3023_ _3277_/CLK _3023_/D vssd1 vssd1 vccd1 vccd1 _3023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2807_ _2803_/X _2804_/X _2805_/X _2806_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2807_/X sky130_fd_sc_hd__mux4_2
X_2738_ _3051_/Q _3355_/Q _3099_/Q _3075_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2738_/X sky130_fd_sc_hd__mux4_2
X_2669_ _3500_/Q _2953_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1971_ _1978_/A vssd1 vssd1 vccd1 vccd1 _1971_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2523_ _2523_/A _2577_/X vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__and2_1
X_2454_ _3398_/Q vssd1 vssd1 vccd1 vccd1 _2454_/Y sky130_fd_sc_hd__inv_2
X_2385_ _3025_/Q _2377_/A _2340_/X _2378_/A vssd1 vssd1 vccd1 vccd1 _3025_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 io_adr_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3006_ _3277_/CLK _3006_/D vssd1 vssd1 vccd1 vccd1 _3006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput371 _3511_/Q vssd1 vssd1 vccd1 vccd1 io_vout[8] sky130_fd_sc_hd__clkbuf_2
Xoutput360 _3514_/Q vssd1 vssd1 vccd1 vccd1 io_irq sky130_fd_sc_hd__clkbuf_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_0 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2170_ _3168_/Q _2165_/X _2144_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1954_ _3298_/Q _1943_/X _1953_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__a22o_1
X_1885_ _3338_/Q _1882_/X _1649_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__a22o_1
X_3486_ _3518_/CLK _3486_/D vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfxtp_1
X_2506_ _3407_/Q vssd1 vssd1 vccd1 vccd1 _2506_/Y sky130_fd_sc_hd__inv_2
X_2437_ _2479_/A _2437_/B vssd1 vssd1 vccd1 vccd1 _2437_/X sky130_fd_sc_hd__and2_1
X_2368_ _2368_/A vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__clkbuf_2
X_2299_ _3081_/Q _2291_/A _2250_/X _2292_/A vssd1 vssd1 vccd1 vccd1 _3081_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1670_ _1730_/A vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__clkbuf_4
X_3340_ _3340_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3271_ _3295_/CLK _3271_/D vssd1 vssd1 vccd1 vccd1 _3271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2222_ _3130_/Q _2215_/A _2148_/X _2216_/A vssd1 vssd1 vccd1 vccd1 _3130_/D sky130_fd_sc_hd__a22o_1
X_2153_ _2172_/A vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _3218_/Q _2081_/X _2044_/X _2082_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__a22o_1
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2986_ _2986_/A0 _2986_/A1 _2986_/A2 _2986_/A3 _2610_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2986_/X sky130_fd_sc_hd__mux4_1
X_1937_ _2046_/A vssd1 vssd1 vccd1 vccd1 _1937_/X sky130_fd_sc_hd__clkbuf_2
X_1868_ _3348_/Q _1864_/X _1818_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__a22o_1
Xinput81 io_b_dat_o_3[13] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_1
Xinput70 io_b_dat_o_2[3] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
Xinput92 io_b_dat_o_3[9] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_1
X_1799_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3469_ _3482_/CLK _3469_/D vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3424_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2840_ _2503_/Y _2441_/Y _2507_/Y _2496_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2840_/X sky130_fd_sc_hd__mux4_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _3101_/Q _3077_/Q _3053_/Q _3357_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2771_/X sky130_fd_sc_hd__mux4_2
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1722_ _1722_/A vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__clkbuf_2
X_1653_ _3441_/Q _1643_/X _1652_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__a22o_1
X_1584_ _1591_/A _2686_/X vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__and2_1
X_3323_ _3443_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
X_3254_ _3279_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
X_2205_ _3143_/Q _2199_/X _2146_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _3143_/D sky130_fd_sc_hd__a22o_1
X_3185_ _3433_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2136_ _2136_/A vssd1 vssd1 vccd1 vccd1 _2136_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2067_ _3229_/Q _2063_/X _2046_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _3423_/Q _3363_/Q _3399_/Q _3395_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2969_/X sky130_fd_sc_hd__mux4_2
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput271 io_dataLastBlock[54] vssd1 vssd1 vccd1 vccd1 _2630_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput260 io_dataLastBlock[44] vssd1 vssd1 vccd1 vccd1 _2587_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput282 io_dataLastBlock[6] vssd1 vssd1 vccd1 vccd1 _2658_/A0 sky130_fd_sc_hd__buf_1
Xinput293 io_dsi_in[7] vssd1 vssd1 vccd1 vccd1 _2464_/B2 sky130_fd_sc_hd__buf_2
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2823_ _3058_/Q _3250_/Q _3226_/Q _3202_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2823_/X sky130_fd_sc_hd__mux4_2
X_2754_ _3296_/Q _3272_/Q _3248_/Q _3224_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2754_/X sky130_fd_sc_hd__mux4_2
X_1705_ _2292_/A vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__clkbuf_2
X_2685_ _1501_/X _3518_/Q _2687_/S vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__mux2_1
X_1636_ _2571_/A vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__clkbuf_2
X_1567_ _1569_/A _2623_/X vssd1 vssd1 vccd1 vccd1 _3492_/D sky130_fd_sc_hd__nor2b_1
X_3306_ _3515_/CLK _3306_/D vssd1 vssd1 vccd1 vccd1 _3306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1498_ _1493_/X _1494_/X _2528_/A _1497_/X vssd1 vssd1 vccd1 vccd1 _1499_/B sky130_fd_sc_hd__o22a_1
X_3237_ _3301_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3168_ _3439_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_1
X_2119_ _3193_/Q _2115_/X _2046_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3099_ _3371_/CLK _3099_/D vssd1 vssd1 vccd1 vccd1 _3099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2470_ _3419_/Q vssd1 vssd1 vccd1 vccd1 _2470_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3022_ _3277_/CLK _3022_/D vssd1 vssd1 vccd1 vccd1 _3022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2806_ _3022_/Q _3014_/Q _3006_/Q _3278_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2806_/X sky130_fd_sc_hd__mux4_2
X_2737_ _2733_/X _2734_/X _2735_/X _2736_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2737_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_22_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3275_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2668_ _2946_/X _2947_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__mux2_1
X_1619_ input7/X vssd1 vssd1 vccd1 vccd1 _1815_/A sky130_fd_sc_hd__buf_1
X_2599_ _2598_/X _2437_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2599_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1970_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2522_ _2522_/A _2522_/B vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__and2_1
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2453_ _3382_/Q vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2384_ _3026_/Q _2377_/A _2338_/X _2378_/A vssd1 vssd1 vccd1 vccd1 _3026_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_adr_i[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3005_ _3277_/CLK _3005_/D vssd1 vssd1 vccd1 vccd1 _3005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput350 _3493_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput361 _3515_/Q vssd1 vssd1 vccd1 vccd1 io_sync_out sky130_fd_sc_hd__clkbuf_2
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput372 _3512_/Q vssd1 vssd1 vccd1 vccd1 io_vout[9] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_1 _2896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1953_ _2559_/A vssd1 vssd1 vccd1 vccd1 _1953_/X sky130_fd_sc_hd__clkbuf_2
X_1884_ _3339_/Q _1882_/X _1645_/X _1883_/X vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__a22o_1
X_3485_ _3485_/CLK _3485_/D vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfxtp_1
X_2505_ _3384_/Q vssd1 vssd1 vccd1 vccd1 _2505_/Y sky130_fd_sc_hd__inv_2
X_2436_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2479_/A sky130_fd_sc_hd__buf_1
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2367_ _2367_/A vssd1 vssd1 vccd1 vccd1 _2367_/X sky130_fd_sc_hd__clkbuf_2
X_2298_ _3082_/Q _2291_/A _2247_/X _2292_/A vssd1 vssd1 vccd1 vccd1 _3082_/D sky130_fd_sc_hd__a22o_1
XFILLER_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3270_ _3294_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3270_/Q sky130_fd_sc_hd__dfxtp_1
X_2221_ _3131_/Q _2215_/X _2146_/X _2216_/X vssd1 vssd1 vccd1 vccd1 _3131_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2152_ _2190_/A _2553_/A vssd1 vssd1 vccd1 vccd1 _2172_/A sky130_fd_sc_hd__or2_4
X_2083_ _3219_/Q _2081_/X _2041_/X _2082_/X vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2985_ input20/X input52/X input68/X input84/X _2610_/S _2611_/S vssd1 vssd1 vccd1
+ vccd1 _2985_/X sky130_fd_sc_hd__mux4_1
X_1936_ _3306_/Q _1931_/X _1935_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _3306_/D sky130_fd_sc_hd__a22o_1
X_1867_ _3349_/Q _1864_/X _1662_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__a22o_1
Xinput82 io_b_dat_o_3[14] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput60 io_b_dat_o_1[9] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 io_b_dat_o_2[4] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
X_1798_ _1846_/A _1798_/B _2224_/C _1798_/D vssd1 vssd1 vccd1 vccd1 _1986_/A sky130_fd_sc_hd__or4_4
Xinput93 io_b_dat_o_4[0] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_1
X_3468_ _3482_/CLK _3468_/D vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ _2429_/A _2419_/B vssd1 vssd1 vccd1 vccd1 _2419_/X sky130_fd_sc_hd__and2_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3399_ _3409_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _3197_/Q _3445_/Q _3149_/Q _3125_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2770_/X sky130_fd_sc_hd__mux4_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _2181_/A vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__clkbuf_2
X_1652_ _2046_/A vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__clkbuf_2
X_1583_ _1592_/A vssd1 vssd1 vccd1 vccd1 _1591_/A sky130_fd_sc_hd__buf_1
X_3322_ _3445_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3253_ _3353_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3184_ _3410_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2204_ _3144_/Q _2199_/X _2144_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _3144_/D sky130_fd_sc_hd__a22o_1
X_2135_ _3184_/Q _1808_/X _2134_/X _1810_/X vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2066_ _3230_/Q _2063_/X _2044_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _3230_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2968_ _3379_/Q _3415_/Q _3431_/Q _3427_/Q _2610_/S _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2968_/X sky130_fd_sc_hd__mux4_2
X_1919_ _3314_/Q _1913_/X _1824_/X _1914_/X vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__a22o_1
X_2899_ _3192_/Q _3440_/Q _3144_/Q _3120_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2899_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput272 io_dataLastBlock[55] vssd1 vssd1 vccd1 vccd1 _2629_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput261 io_dataLastBlock[45] vssd1 vssd1 vccd1 vccd1 _2584_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput250 io_dataLastBlock[35] vssd1 vssd1 vccd1 vccd1 _2670_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput283 io_dataLastBlock[7] vssd1 vssd1 vccd1 vccd1 _2654_/A0 sky130_fd_sc_hd__buf_1
Xinput294 io_we_i vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__buf_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2822_ _2818_/X _2819_/X _2820_/X _2821_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2822_/X sky130_fd_sc_hd__mux4_2
X_2753_ _3176_/Q _3344_/Q _3328_/Q _3312_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2753_/X sky130_fd_sc_hd__mux4_2
X_1704_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2292_/A sky130_fd_sc_hd__inv_2
X_2684_ _2998_/X _2999_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__mux2_1
X_1635_ _3447_/Q _1629_/X _1634_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__a22o_1
X_1566_ _1569_/A _2622_/X vssd1 vssd1 vccd1 vccd1 _3493_/D sky130_fd_sc_hd__nor2b_2
X_3305_ _3307_/CLK _3305_/D vssd1 vssd1 vccd1 vccd1 _3305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1497_ _1497_/A _3450_/Q _3452_/Q _3451_/Q vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__or4_4
X_3236_ _3301_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167_ _3439_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2118_ _3194_/Q _2115_/X _2044_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__a22o_1
X_3098_ _3335_/CLK _3098_/D vssd1 vssd1 vccd1 vccd1 _3098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2049_ _3240_/Q _2040_/X _2048_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _3240_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3021_ _3087_/CLK _3021_/D vssd1 vssd1 vccd1 vccd1 _3021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2805_ _3086_/Q _3370_/Q _3038_/Q _3030_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2805_/X sky130_fd_sc_hd__mux4_2
X_2736_ _3322_/Q _3306_/Q _3170_/Q _3338_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2736_/X sky130_fd_sc_hd__mux4_1
X_2667_ _2945_/X _2666_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__mux2_2
X_1618_ _1618_/A _2620_/X vssd1 vssd1 vccd1 vccd1 _3449_/D sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_62_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3474_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2598_ _2598_/A0 _2598_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__mux2_1
X_1549_ _3499_/Q _1539_/X _1726_/A _1541_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _3499_/D
+ sky130_fd_sc_hd__o221a_1
X_3219_ _3303_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2521_ _3416_/Q vssd1 vssd1 vccd1 vccd1 _2521_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2452_ _3406_/Q vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__inv_2
X_2383_ _3027_/Q _2377_/X _2336_/X _2378_/X vssd1 vssd1 vccd1 vccd1 _3027_/D sky130_fd_sc_hd__a22o_1
X_3004_ _3277_/CLK _3004_/D vssd1 vssd1 vccd1 vccd1 _3004_/Q sky130_fd_sc_hd__dfxtp_1
Xinput3 io_adr_i[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2719_ _3143_/Q _3119_/Q _3191_/Q _3439_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2719_/X sky130_fd_sc_hd__mux4_1
Xoutput351 _3494_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput340 _3484_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput362 _3503_/Q vssd1 vssd1 vccd1 vccd1 io_vout[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_2 _2630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1952_ _3299_/Q _1943_/X _1951_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__a22o_1
X_1883_ _1890_/A vssd1 vssd1 vccd1 vccd1 _1883_/X sky130_fd_sc_hd__clkbuf_2
X_3484_ _3485_/CLK _3484_/D vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfxtp_1
X_2504_ _3412_/Q vssd1 vssd1 vccd1 vccd1 _2504_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _3392_/Q vssd1 vssd1 vccd1 vccd1 _2435_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2366_ _3040_/Q _1761_/X _2324_/X _1763_/X vssd1 vssd1 vccd1 vccd1 _3040_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2297_ _3083_/Q _2291_/X _2244_/X _2292_/X vssd1 vssd1 vccd1 vccd1 _3083_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2220_ _3132_/Q _2215_/X _2144_/X _2216_/X vssd1 vssd1 vccd1 vccd1 _3132_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2151_ _3177_/Q _2136_/A _2150_/X _2138_/A vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__a22o_1
X_2082_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2984_ _2980_/X _2981_/X _2982_/X _2983_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2984_/X sky130_fd_sc_hd__mux4_1
X_1935_ _2044_/A vssd1 vssd1 vccd1 vccd1 _1935_/X sky130_fd_sc_hd__buf_2
X_1866_ _3350_/Q _1864_/X _1659_/X _1865_/X vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__a22o_1
Xinput50 io_b_dat_o_1[14] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput72 io_b_dat_o_2[5] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_1
Xinput61 io_b_dat_o_2[0] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
X_1797_ _3385_/Q _1791_/X _1778_/X _1793_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__a22o_1
Xinput83 io_b_dat_o_3[15] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
Xinput94 io_b_dat_o_4[10] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3467_ _3482_/CLK _3467_/D vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2418_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2429_/A sky130_fd_sc_hd__buf_1
X_3398_ _3398_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2349_ _3053_/Q _2343_/X _2570_/A _2345_/X vssd1 vssd1 vccd1 vccd1 _3053_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _1760_/A _2548_/A vssd1 vssd1 vccd1 vccd1 _2181_/A sky130_fd_sc_hd__or2_4
X_1651_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2046_/A sky130_fd_sc_hd__clkbuf_2
X_1582_ _1582_/A _2636_/X vssd1 vssd1 vccd1 vccd1 _3479_/D sky130_fd_sc_hd__nor2b_1
X_3321_ _3443_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
X_3252_ _3279_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
X_3183_ _3456_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
X_2203_ _3145_/Q _2199_/X _2142_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _3145_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2134_ _2569_/A vssd1 vssd1 vccd1 vccd1 _2134_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2065_ _3231_/Q _2063_/X _2041_/X _2064_/X vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3500_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2967_ _3419_/Q _3375_/Q _3391_/Q _3387_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2967_/X sky130_fd_sc_hd__mux4_2
X_1918_ _3315_/Q _1913_/X _1822_/X _1914_/X vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__a22o_1
X_2898_ _3288_/Q _3264_/Q _3240_/Q _3216_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2898_/X sky130_fd_sc_hd__mux4_2
X_1849_ _1864_/A vssd1 vssd1 vccd1 vccd1 _1849_/X sky130_fd_sc_hd__buf_2
X_3519_ _3519_/CLK _3519_/D vssd1 vssd1 vccd1 vccd1 _3519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput262 io_dataLastBlock[46] vssd1 vssd1 vccd1 vccd1 _2581_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput240 io_dataLastBlock[26] vssd1 vssd1 vccd1 vccd1 _2626_/A0 sky130_fd_sc_hd__buf_1
XFILLER_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput251 io_dataLastBlock[36] vssd1 vssd1 vccd1 vccd1 _2666_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput295 wb_rst_i vssd1 vssd1 vccd1 vccd1 _1590_/A sky130_fd_sc_hd__buf_4
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput273 io_dataLastBlock[56] vssd1 vssd1 vccd1 vccd1 _2628_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput284 io_dataLastBlock[8] vssd1 vssd1 vccd1 vccd1 _2650_/A0 sky130_fd_sc_hd__buf_1
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2821_ _3019_/Q _3011_/Q _3003_/Q _3275_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2821_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2752_ _2748_/X _2749_/X _2750_/X _2751_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2752_/X sky130_fd_sc_hd__mux4_2
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1703_ _2291_/A vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__clkbuf_2
X_2683_ _2997_/X _2682_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2683_/X sky130_fd_sc_hd__mux2_1
X_1634_ _2572_/A vssd1 vssd1 vccd1 vccd1 _1634_/X sky130_fd_sc_hd__clkbuf_2
X_1565_ _1569_/A _2621_/X vssd1 vssd1 vccd1 vccd1 _3494_/D sky130_fd_sc_hd__nor2b_1
X_3304_ _3515_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1496_ _3449_/Q vssd1 vssd1 vccd1 vccd1 _1497_/A sky130_fd_sc_hd__inv_2
X_3235_ _3474_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3166_ _3433_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2117_ _3195_/Q _2115_/X _2041_/X _2116_/X vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__a22o_1
X_3097_ _3371_/CLK _3097_/D vssd1 vssd1 vccd1 vccd1 _3097_/Q sky130_fd_sc_hd__dfxtp_1
X_2048_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__buf_2
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_3020_ _3277_/CLK _3020_/D vssd1 vssd1 vccd1 vccd1 _3020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2804_ _3182_/Q _3158_/Q _3134_/Q _3110_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2804_/X sky130_fd_sc_hd__mux4_1
X_2735_ _3242_/Q _3218_/Q _3290_/Q _3266_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2735_/X sky130_fd_sc_hd__mux4_2
X_2666_ _2666_/A0 _2666_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__mux2_2
X_1617_ _1618_/A _2619_/X vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__and2_1
X_2597_ _2596_/X _2446_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__mux2_1
X_1548_ _2560_/A vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__buf_2
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3218_ _3514_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3279_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3445_/CLK _3149_/D vssd1 vssd1 vccd1 vccd1 _3149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2520_ _2520_/A _2578_/X vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__and2_1
X_2451_ _2490_/A _2792_/X vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__and2_1
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2382_ _3028_/Q _2377_/X _2334_/X _2378_/X vssd1 vssd1 vccd1 vccd1 _3028_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3003_ _3019_/CLK _3003_/D vssd1 vssd1 vccd1 vccd1 _3003_/Q sky130_fd_sc_hd__dfxtp_1
Xinput4 io_adr_i[1] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2718_ _3047_/Q _3351_/Q _3095_/Q _3071_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2718_/X sky130_fd_sc_hd__mux4_2
X_2649_ _2886_/X _2887_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2649_/X sky130_fd_sc_hd__mux2_1
Xoutput341 _3485_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput330 _3469_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput352 _3460_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput363 _3513_/Q vssd1 vssd1 vccd1 vccd1 io_vout[10] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_3 _2621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1951_ _2560_/A vssd1 vssd1 vccd1 vccd1 _1951_/X sky130_fd_sc_hd__clkbuf_2
X_1882_ _1889_/A vssd1 vssd1 vccd1 vccd1 _1882_/X sky130_fd_sc_hd__clkbuf_2
X_2503_ _3423_/Q vssd1 vssd1 vccd1 vccd1 _2503_/Y sky130_fd_sc_hd__inv_2
X_3483_ _3485_/CLK _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfxtp_1
X_2434_ _3388_/Q vssd1 vssd1 vccd1 vccd1 _2434_/Y sky130_fd_sc_hd__inv_2
X_2365_ _3041_/Q _2358_/A _1730_/A _2359_/A vssd1 vssd1 vccd1 vccd1 _3041_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2296_ _3084_/Q _2291_/X _2242_/X _2292_/X vssd1 vssd1 vccd1 vccd1 _3084_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2150_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2150_/X sky130_fd_sc_hd__buf_2
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2081_ _2088_/A vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2983_ _3406_/Q _3402_/Q _3410_/Q _3382_/Q _2610_/S _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2983_/X sky130_fd_sc_hd__mux4_1
X_1934_ _3307_/Q _1931_/X _1932_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _3307_/D sky130_fd_sc_hd__a22o_1
Xinput40 io_b_dat_o_10[5] vssd1 vssd1 vccd1 vccd1 _2429_/B sky130_fd_sc_hd__clkbuf_1
X_1865_ _1865_/A vssd1 vssd1 vccd1 vccd1 _1865_/X sky130_fd_sc_hd__clkbuf_2
Xinput51 io_b_dat_o_1[15] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 io_b_dat_o_2[10] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
Xinput73 io_b_dat_o_2[6] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
X_1796_ _3386_/Q _1791_/X _1776_/X _1793_/X vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__a22o_1
Xinput95 io_b_dat_o_4[11] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_1
Xinput84 io_b_dat_o_3[1] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
X_3466_ _3485_/CLK _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2417_ _2607_/X _2487_/A vssd1 vssd1 vccd1 vccd1 _2417_/X sky130_fd_sc_hd__and2_1
X_3397_ _3420_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
X_2348_ _3054_/Q _2343_/X _2571_/A _2345_/X vssd1 vssd1 vccd1 vccd1 _3054_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2279_ _3097_/Q _2275_/X _2240_/X _2276_/X vssd1 vssd1 vccd1 vccd1 _3097_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650_ _3442_/Q _1643_/X _1649_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__a22o_1
X_1581_ _1581_/A _2635_/X vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__nor2b_4
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3320_ _3336_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
X_3251_ _3371_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3182_ _3456_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2202_ _3146_/Q _2199_/X _2140_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _3146_/D sky130_fd_sc_hd__a22o_1
X_2133_ _3185_/Q _2122_/A _2132_/X _2123_/A vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2064_ _2064_/A vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__buf_2
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3334_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2966_ _2962_/X _2963_/X _2964_/X _2965_/X input7/X input8/X vssd1 vssd1 vccd1 vccd1
+ _2966_/X sky130_fd_sc_hd__mux4_2
X_1917_ _3316_/Q _1913_/X _1818_/X _1914_/X vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__a22o_1
X_2897_ _3168_/Q _3336_/Q _3320_/Q _3304_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2897_/X sky130_fd_sc_hd__mux4_1
X_1848_ _2487_/A _2342_/B _2224_/C _2300_/D vssd1 vssd1 vccd1 vccd1 _1864_/A sky130_fd_sc_hd__or4_4
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1779_ _3393_/Q _1769_/X _1778_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__a22o_1
X_3518_ _3518_/CLK _3518_/D vssd1 vssd1 vccd1 vccd1 _3518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3449_ _3519_/CLK _3449_/D vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput263 io_dataLastBlock[47] vssd1 vssd1 vccd1 vccd1 _2578_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput230 io_dataLastBlock[17] vssd1 vssd1 vccd1 vccd1 _2635_/A0 sky130_fd_sc_hd__buf_1
Xinput241 io_dataLastBlock[27] vssd1 vssd1 vccd1 vccd1 _2625_/A0 sky130_fd_sc_hd__buf_1
Xinput252 io_dataLastBlock[37] vssd1 vssd1 vccd1 vccd1 _2662_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput274 io_dataLastBlock[57] vssd1 vssd1 vccd1 vccd1 _2627_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput285 io_dataLastBlock[9] vssd1 vssd1 vccd1 vccd1 _2647_/A0 sky130_fd_sc_hd__buf_1
XFILLER_48_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2820_ _3083_/Q _3367_/Q _3035_/Q _3027_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2820_/X sky130_fd_sc_hd__mux4_1
X_2751_ _3325_/Q _3309_/Q _3173_/Q _3341_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2751_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2682_ _2682_/A0 _2682_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2682_/X sky130_fd_sc_hd__mux2_4
X_1702_ _1760_/A _2544_/A vssd1 vssd1 vccd1 vccd1 _2291_/A sky130_fd_sc_hd__or2_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1633_ _3448_/Q _1629_/X _1630_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__a22o_1
X_1564_ _1582_/A vssd1 vssd1 vccd1 vccd1 _1569_/A sky130_fd_sc_hd__clkbuf_2
X_1495_ _3454_/Q _3455_/Q _3453_/Q _3456_/Q vssd1 vssd1 vccd1 vccd1 _2528_/A sky130_fd_sc_hd__or4_4
X_3303_ _3303_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
X_3234_ _3331_/CLK _3234_/D vssd1 vssd1 vccd1 vccd1 _3234_/Q sky130_fd_sc_hd__dfxtp_1
X_3165_ _3438_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_1
X_2116_ _2123_/A vssd1 vssd1 vccd1 vccd1 _2116_/X sky130_fd_sc_hd__buf_2
X_3096_ _3351_/CLK _3096_/D vssd1 vssd1 vccd1 vccd1 _3096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2047_ _3241_/Q _2040_/X _2046_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2949_ _3164_/Q _3332_/Q _3316_/Q _3300_/Q _1700_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2949_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_1_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3346_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2803_ _3062_/Q _3254_/Q _3230_/Q _3206_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2803_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2734_ _3146_/Q _3122_/Q _3194_/Q _3442_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2734_/X sky130_fd_sc_hd__mux4_2
X_2665_ _3501_/Q _2940_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__mux2_1
X_2596_ _2596_/A0 _2596_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__mux2_1
X_1616_ _1618_/A _2618_/X vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__and2_1
X_1547_ _3500_/Q _1539_/X _1722_/A _1541_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _3500_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3217_ _3307_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3148_ _3336_/CLK _3148_/D vssd1 vssd1 vccd1 vccd1 _3148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3079_ _3448_/CLK _3079_/D vssd1 vssd1 vccd1 vccd1 _3079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2450_ _2520_/A vssd1 vssd1 vccd1 vccd1 _2490_/A sky130_fd_sc_hd__buf_1
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2381_ _3029_/Q _2377_/X _2332_/X _2378_/X vssd1 vssd1 vccd1 vccd1 _3029_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3002_ _3019_/CLK _3002_/D vssd1 vssd1 vccd1 vccd1 _3002_/Q sky130_fd_sc_hd__dfxtp_1
Xinput5 io_adr_i[2] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2717_ _2713_/X _2714_/X _2715_/X _2716_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2717_/X sky130_fd_sc_hd__mux4_2
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput342 _3486_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput331 _3470_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[13] sky130_fd_sc_hd__clkbuf_2
X_2648_ _2885_/X _2647_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2648_/X sky130_fd_sc_hd__mux2_2
Xoutput320 _2562_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[4] sky130_fd_sc_hd__clkbuf_2
Xoutput353 _3461_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[4] sky130_fd_sc_hd__clkbuf_2
X_2579_ _2579_/A0 _2579_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2579_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput364 _3504_/Q vssd1 vssd1 vccd1 vccd1 io_vout[1] sky130_fd_sc_hd__clkbuf_2
XINSDIODE3_4 _2670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _3300_/Q _1943_/X _1949_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__a22o_1
X_1881_ _3340_/Q _1874_/X _1641_/X _1876_/X vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__a22o_1
X_2502_ _3404_/Q vssd1 vssd1 vccd1 vccd1 _2502_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3482_ _3482_/CLK _3482_/D vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfxtp_1
X_2433_ _3418_/Q vssd1 vssd1 vccd1 vccd1 _2433_/Y sky130_fd_sc_hd__inv_2
X_2364_ _3042_/Q _2358_/X _1728_/A _2359_/X vssd1 vssd1 vccd1 vccd1 _3042_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2295_ _3085_/Q _2291_/X _2240_/X _2292_/X vssd1 vssd1 vccd1 vccd1 _3085_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2080_ _3220_/Q _2073_/X _2038_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _3422_/Q _3362_/Q _3398_/Q _3394_/Q _2982_/S0 _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2982_/X sky130_fd_sc_hd__mux4_1
X_1933_ _1945_/A vssd1 vssd1 vccd1 vccd1 _1933_/X sky130_fd_sc_hd__clkbuf_2
Xinput30 io_b_dat_o_10[10] vssd1 vssd1 vccd1 vccd1 _2479_/B sky130_fd_sc_hd__clkbuf_1
X_1864_ _1864_/A vssd1 vssd1 vccd1 vccd1 _1864_/X sky130_fd_sc_hd__clkbuf_2
Xinput63 io_b_dat_o_2[11] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
Xinput41 io_b_dat_o_10[6] vssd1 vssd1 vccd1 vccd1 _2437_/B sky130_fd_sc_hd__clkbuf_1
Xinput52 io_b_dat_o_1[1] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
X_1795_ _3387_/Q _1791_/X _1774_/X _1793_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__a22o_1
Xinput74 io_b_dat_o_2[7] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
Xinput96 io_b_dat_o_4[12] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_1
Xinput85 io_b_dat_o_3[2] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
X_3465_ _3493_/CLK _3465_/D vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfxtp_1
X_2416_ _2416_/A _2485_/A vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__and2_1
X_3396_ _3420_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
X_2347_ _3055_/Q _2343_/X _2572_/A _2345_/X vssd1 vssd1 vccd1 vccd1 _3055_/D sky130_fd_sc_hd__a22o_1
X_2278_ _3098_/Q _2275_/X _2238_/X _2276_/X vssd1 vssd1 vccd1 vccd1 _3098_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _1581_/A _2634_/X vssd1 vssd1 vccd1 vccd1 _3481_/D sky130_fd_sc_hd__nor2b_4
XFILLER_22_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3250_ _3367_/CLK _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/Q sky130_fd_sc_hd__dfxtp_1
X_3181_ _3456_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
X_2201_ _3147_/Q _2199_/X _2137_/X _2200_/X vssd1 vssd1 vccd1 vccd1 _3147_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2132_ _2558_/A vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2063_ _2063_/A vssd1 vssd1 vccd1 vccd1 _2063_/X sky130_fd_sc_hd__buf_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2965_ _3091_/Q _3067_/Q _3043_/Q _3347_/Q _1676_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2965_/X sky130_fd_sc_hd__mux4_1
X_2896_ _2451_/X _2651_/X _2652_/X _2456_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2896_/X sky130_fd_sc_hd__mux4_2
X_1916_ _3317_/Q _1913_/X _1662_/X _1914_/X vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1847_ _1847_/A vssd1 vssd1 vccd1 vccd1 _2342_/B sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3180_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3517_ _3518_/CLK _3517_/D vssd1 vssd1 vccd1 vccd1 _3517_/Q sky130_fd_sc_hd__dfxtp_1
X_1778_ _2558_/A vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__clkbuf_2
X_3448_ _3448_/CLK _3448_/D vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfxtp_1
X_3379_ _3482_/CLK _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput220 io_dat_i[8] vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput231 io_dataLastBlock[18] vssd1 vssd1 vccd1 vccd1 _2634_/A0 sky130_fd_sc_hd__buf_1
Xinput242 io_dataLastBlock[28] vssd1 vssd1 vccd1 vccd1 _2624_/A0 sky130_fd_sc_hd__buf_1
Xinput253 io_dataLastBlock[38] vssd1 vssd1 vccd1 vccd1 _2658_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput275 io_dataLastBlock[58] vssd1 vssd1 vccd1 vccd1 _2626_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput286 io_dsi_in[0] vssd1 vssd1 vccd1 vccd1 _2459_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput264 io_dataLastBlock[48] vssd1 vssd1 vccd1 vccd1 _2636_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _3245_/Q _3221_/Q _3293_/Q _3269_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2750_/X sky130_fd_sc_hd__mux4_2
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2681_ _3502_/Q _2992_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__mux2_4
X_1701_ _2224_/A _1847_/A _2266_/C vssd1 vssd1 vccd1 vccd1 _2544_/A sky130_fd_sc_hd__or3_4
X_1632_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__buf_2
X_1563_ _1626_/A _2575_/S _1590_/A _1678_/C vssd1 vssd1 vccd1 vccd1 _1582_/A sky130_fd_sc_hd__or4_4
X_1494_ _2797_/X _2802_/X _2807_/X _2812_/X vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__or4_4
X_3302_ _3334_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
X_3233_ _3297_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3164_ _3333_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2115_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2115_/X sky130_fd_sc_hd__buf_2
X_3095_ _3351_/CLK _3095_/D vssd1 vssd1 vccd1 vccd1 _3095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2046_ _2046_/A vssd1 vssd1 vccd1 vccd1 _2046_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2948_ _2665_/X _2667_/X _2668_/X _2427_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2948_/X sky130_fd_sc_hd__mux4_2
X_2879_ input94/X _2879_/A1 _2879_/A2 _2879_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2879_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_10 _2573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2802_ _2798_/X _2799_/X _2800_/X _2801_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2802_/X sky130_fd_sc_hd__mux4_2
X_2733_ _3050_/Q _3354_/Q _3098_/Q _3074_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2733_/X sky130_fd_sc_hd__mux4_2
X_2664_ _2933_/X _2934_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__mux2_1
X_2595_ _2594_/X _2455_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__mux2_1
X_1615_ _1615_/A _2617_/X vssd1 vssd1 vccd1 vccd1 _3452_/D sky130_fd_sc_hd__and2_1
X_1546_ _2561_/A vssd1 vssd1 vccd1 vccd1 _1722_/A sky130_fd_sc_hd__buf_2
XFILLER_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3216_ _3307_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3147_ _3335_/CLK _3147_/D vssd1 vssd1 vccd1 vccd1 _3147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3078_ _3447_/CLK _3078_/D vssd1 vssd1 vccd1 vccd1 _3078_/Q sky130_fd_sc_hd__dfxtp_1
X_2029_ _2342_/D vssd1 vssd1 vccd1 vccd1 _2190_/A sky130_fd_sc_hd__buf_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3307_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2380_ _3030_/Q _2377_/X _2330_/X _2378_/X vssd1 vssd1 vccd1 vccd1 _3030_/D sky130_fd_sc_hd__a22o_1
X_3001_ _3501_/CLK _3001_/D vssd1 vssd1 vccd1 vccd1 _3001_/Q sky130_fd_sc_hd__dfxtp_1
Xinput6 io_adr_i[3] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2716_ _3318_/Q _3302_/Q _3166_/Q _3334_/Q _2716_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2716_/X sky130_fd_sc_hd__mux4_1
Xoutput310 _2558_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[0] sky130_fd_sc_hd__clkbuf_2
X_2647_ _2647_/A0 _2647_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__mux2_1
Xoutput343 _3487_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput332 _3471_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput321 _2563_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2578_ _2578_/A0 _2578_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2578_/X sky130_fd_sc_hd__mux2_1
Xoutput354 _3462_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput365 _3505_/Q vssd1 vssd1 vccd1 vccd1 io_vout[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE3_5 _3480_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1529_ _1523_/X _3506_/Q _1524_/X _2707_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _3506_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1880_ _3341_/Q _1874_/X _1638_/X _1876_/X vssd1 vssd1 vccd1 vccd1 _3341_/D sky130_fd_sc_hd__a22o_1
X_2501_ _3408_/Q vssd1 vssd1 vccd1 vccd1 _2501_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3481_ _3482_/CLK _3481_/D vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2432_ _3374_/Q vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__inv_2
X_2363_ _3043_/Q _2358_/X _1726_/A _2359_/X vssd1 vssd1 vccd1 vccd1 _3043_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2294_ _3086_/Q _2291_/X _2238_/X _2292_/X vssd1 vssd1 vccd1 vccd1 _3086_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2981_ _3378_/Q _3414_/Q _3430_/Q _3426_/Q _2610_/S _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2981_/X sky130_fd_sc_hd__mux4_2
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1932_ _2041_/A vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__clkbuf_2
X_1863_ _3351_/Q _1857_/X _1656_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__a22o_1
Xinput31 io_b_dat_o_10[11] vssd1 vssd1 vccd1 vccd1 _2486_/B sky130_fd_sc_hd__clkbuf_1
Xinput20 io_b_dat_o_0[1] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
Xinput42 io_b_dat_o_10[7] vssd1 vssd1 vccd1 vccd1 _2446_/B sky130_fd_sc_hd__clkbuf_1
Xinput53 io_b_dat_o_1[2] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 io_b_dat_o_2[12] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
X_1794_ _3388_/Q _1791_/X _1770_/X _1793_/X vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__a22o_1
Xinput75 io_b_dat_o_2[8] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
Xinput86 io_b_dat_o_3[3] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_1
Xinput97 io_b_dat_o_4[13] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_1
X_3464_ _3493_/CLK _3464_/D vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2415_ _3001_/Q _2407_/A _1947_/A _2408_/A vssd1 vssd1 vccd1 vccd1 _3001_/D sky130_fd_sc_hd__a22o_1
X_3395_ _3423_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
X_2346_ _3056_/Q _2343_/X _2573_/A _2345_/X vssd1 vssd1 vccd1 vccd1 _3056_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2277_ _3099_/Q _2275_/X _2235_/X _2276_/X vssd1 vssd1 vccd1 vccd1 _3099_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2200_ _2207_/A vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__clkbuf_2
X_3180_ _3180_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_1
X_2131_ _3186_/Q _2122_/X _2130_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2062_ _3232_/Q _1782_/X _2038_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _3232_/D sky130_fd_sc_hd__a22o_1
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2964_ _3187_/Q _3435_/Q _3139_/Q _3115_/Q _1676_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2964_/X sky130_fd_sc_hd__mux4_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1915_ _3318_/Q _1913_/X _1659_/X _1914_/X vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__a22o_1
X_2895_ _2895_/A0 _2895_/A1 _2895_/A2 _2895_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2895_/X sky130_fd_sc_hd__mux4_1
X_1846_ _1846_/A vssd1 vssd1 vccd1 vccd1 _2487_/A sky130_fd_sc_hd__clkbuf_4
X_1777_ _3394_/Q _1769_/X _1776_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__a22o_1
X_3516_ _3519_/CLK _3516_/D vssd1 vssd1 vccd1 vccd1 _3516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3447_ _3447_/CLK _3447_/D vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3378_ _3500_/CLK _3378_/D vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2329_ _3063_/Q _2326_/X _2327_/X _2328_/X vssd1 vssd1 vccd1 vccd1 _3063_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput210 io_dat_i[28] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__buf_1
XFILLER_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput221 io_dat_i[9] vssd1 vssd1 vccd1 vccd1 _2567_/A sky130_fd_sc_hd__clkbuf_4
Xinput232 io_dataLastBlock[19] vssd1 vssd1 vccd1 vccd1 _2633_/A0 sky130_fd_sc_hd__buf_1
Xinput243 io_dataLastBlock[29] vssd1 vssd1 vccd1 vccd1 _2623_/A0 sky130_fd_sc_hd__buf_1
Xinput254 io_dataLastBlock[39] vssd1 vssd1 vccd1 vccd1 _2654_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput276 io_dataLastBlock[59] vssd1 vssd1 vccd1 vccd1 _2625_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput287 io_dsi_in[1] vssd1 vssd1 vccd1 vccd1 _2459_/B2 sky130_fd_sc_hd__clkbuf_1
Xinput265 io_dataLastBlock[49] vssd1 vssd1 vccd1 vccd1 _2635_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_90_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _2985_/X _2986_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1700_ _1700_/A _1700_/B vssd1 vssd1 vccd1 vccd1 _2266_/C sky130_fd_sc_hd__or2_2
X_1631_ _1658_/A vssd1 vssd1 vccd1 vccd1 _1660_/A sky130_fd_sc_hd__inv_2
X_1562_ _2557_/A vssd1 vssd1 vccd1 vccd1 _1678_/C sky130_fd_sc_hd__inv_2
X_3301_ _3301_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
X_1493_ _2817_/X _2822_/X _2827_/X _2832_/X vssd1 vssd1 vccd1 vccd1 _1493_/X sky130_fd_sc_hd__or4_4
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3232_ _3372_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
X_3163_ _3333_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_1
X_2114_ _3196_/Q _2107_/X _2038_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__a22o_1
X_3094_ _3350_/CLK _3094_/D vssd1 vssd1 vccd1 vccd1 _3094_/Q sky130_fd_sc_hd__dfxtp_1
X_2045_ _3242_/Q _2040_/X _2044_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _3242_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2947_ _2947_/A0 _2947_/A1 _2947_/A2 _2947_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2947_/X sky130_fd_sc_hd__mux4_1
X_2878_ input14/X input46/X input62/X input78/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2878_/X sky130_fd_sc_hd__mux4_1
X_1829_ _1837_/A vssd1 vssd1 vccd1 vccd1 _1829_/X sky130_fd_sc_hd__buf_2
XFILLER_2_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_11 _2463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2801_ _3023_/Q _3015_/Q _3007_/Q _3279_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2801_/X sky130_fd_sc_hd__mux4_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2732_ _2728_/X _2729_/X _2730_/X _2731_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2732_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _2932_/X _2662_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2663_/X sky130_fd_sc_hd__mux2_2
X_2594_ _2594_/A0 _2594_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__mux2_1
X_1614_ _1615_/A _2616_/X vssd1 vssd1 vccd1 vccd1 _3453_/D sky130_fd_sc_hd__and2_1
X_1545_ _3501_/Q _1539_/X _1947_/A _1541_/X _1544_/X vssd1 vssd1 vccd1 vccd1 _3501_/D
+ sky130_fd_sc_hd__o221a_1
X_3215_ _3303_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3146_ _3443_/CLK _3146_/D vssd1 vssd1 vccd1 vccd1 _3146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _3336_/CLK _3077_/D vssd1 vssd1 vccd1 vccd1 _3077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2028_ _3249_/Q _2020_/A _1947_/X _2021_/A vssd1 vssd1 vccd1 vccd1 _3249_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _2681_/X _2683_/X _2684_/X _2423_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _3000_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 io_adr_i[4] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2715_ _3238_/Q _3214_/Q _3286_/Q _3262_/Q _2716_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2715_/X sky130_fd_sc_hd__mux4_2
X_2646_ _2878_/X _2879_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2646_/X sky130_fd_sc_hd__mux2_1
Xoutput300 _2552_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_1 sky130_fd_sc_hd__clkbuf_2
Xoutput344 _3488_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput333 _3472_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput322 _2564_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[6] sky130_fd_sc_hd__clkbuf_2
Xoutput311 _2568_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[10] sky130_fd_sc_hd__clkbuf_2
X_2577_ _2576_/X _2522_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__mux2_1
Xoutput355 _3463_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput366 _3506_/Q vssd1 vssd1 vccd1 vccd1 io_vout[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE3_6 _3481_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1528_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__clkbuf_4
X_3129_ _3501_/CLK _3129_/D vssd1 vssd1 vccd1 vccd1 _3129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2500_ _2523_/A _2583_/X vssd1 vssd1 vccd1 vccd1 _2500_/X sky130_fd_sc_hd__and2_1
X_3480_ _3482_/CLK _3480_/D vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2431_ _3390_/Q vssd1 vssd1 vccd1 vccd1 _2431_/Y sky130_fd_sc_hd__inv_2
X_2362_ _3044_/Q _2358_/X _1722_/A _2359_/X vssd1 vssd1 vccd1 vccd1 _3044_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2293_ _3087_/Q _2291_/X _2235_/X _2292_/X vssd1 vssd1 vccd1 vccd1 _3087_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2629_ _2629_/A0 _2629_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2629_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _3418_/Q _3374_/Q _3390_/Q _3386_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2980_/X sky130_fd_sc_hd__mux4_2
X_1931_ _1943_/A vssd1 vssd1 vccd1 vccd1 _1931_/X sky130_fd_sc_hd__clkbuf_2
X_1862_ _3352_/Q _1857_/X _1654_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__a22o_1
Xinput21 io_b_dat_o_0[2] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_1
Xinput10 io_adr_i[7] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput32 io_b_dat_o_10[12] vssd1 vssd1 vccd1 vccd1 _2493_/B sky130_fd_sc_hd__clkbuf_1
Xinput43 io_b_dat_o_10[8] vssd1 vssd1 vccd1 vccd1 _2455_/B sky130_fd_sc_hd__clkbuf_1
Xinput54 io_b_dat_o_1[3] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
X_1793_ _2098_/A vssd1 vssd1 vccd1 vccd1 _1793_/X sky130_fd_sc_hd__clkbuf_2
Xinput65 io_b_dat_o_2[13] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
Xinput87 io_b_dat_o_3[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput98 io_b_dat_o_4[14] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_1
Xinput76 io_b_dat_o_2[9] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
X_3463_ _3500_/CLK _3463_/D vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfxtp_1
X_2414_ _3002_/Q _2407_/A _1944_/A _2408_/A vssd1 vssd1 vccd1 vccd1 _3002_/D sky130_fd_sc_hd__a22o_1
X_3394_ _3424_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
X_2345_ _2359_/A vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__clkbuf_2
X_2276_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2276_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2130_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2061_ _3233_/Q _2052_/A _1955_/X _2054_/A vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ _3283_/Q _3259_/Q _3235_/Q _3211_/Q input5/X input6/X vssd1 vssd1 vccd1 vccd1
+ _2963_/X sky130_fd_sc_hd__mux4_2
X_1914_ _1914_/A vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__clkbuf_2
X_2894_ input27/X input59/X input75/X input91/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2894_/X sky130_fd_sc_hd__mux4_1
X_1845_ _3361_/Q _1837_/A _1826_/X _1838_/A vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__a22o_1
X_1776_ _2559_/A vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__clkbuf_2
X_3515_ _3515_/CLK _3515_/D vssd1 vssd1 vccd1 vccd1 _3515_/Q sky130_fd_sc_hd__dfxtp_1
X_3446_ _3506_/CLK _3446_/D vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfxtp_1
X_3377_ _3429_/CLK _3377_/D vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2328_ _2328_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2259_ _3111_/Q _2257_/X _2235_/X _2258_/X vssd1 vssd1 vccd1 vccd1 _3111_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3371_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput200 io_dat_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__buf_1
Xinput211 io_dat_i[29] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput233 io_dataLastBlock[1] vssd1 vssd1 vccd1 vccd1 _2678_/A0 sky130_fd_sc_hd__buf_1
Xinput244 io_dataLastBlock[2] vssd1 vssd1 vccd1 vccd1 _2674_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput222 io_dataLastBlock[0] vssd1 vssd1 vccd1 vccd1 _2682_/A0 sky130_fd_sc_hd__buf_1
Xinput288 io_dsi_in[2] vssd1 vssd1 vccd1 vccd1 _2461_/A2 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput277 io_dataLastBlock[5] vssd1 vssd1 vccd1 vccd1 _2662_/A0 sky130_fd_sc_hd__buf_1
Xinput255 io_dataLastBlock[3] vssd1 vssd1 vccd1 vccd1 _2670_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput266 io_dataLastBlock[4] vssd1 vssd1 vccd1 vccd1 _2666_/A0 sky130_fd_sc_hd__buf_1
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1630_ _2573_/A vssd1 vssd1 vccd1 vccd1 _1630_/X sky130_fd_sc_hd__clkbuf_2
X_1561_ _2520_/A vssd1 vssd1 vccd1 vccd1 _1626_/A sky130_fd_sc_hd__inv_2
X_3300_ _3333_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_1
X_1492_ _3502_/Q vssd1 vssd1 vccd1 vccd1 _1513_/A sky130_fd_sc_hd__inv_2
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3231_ _3279_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
X_3162_ _3333_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_1
X_2113_ _3197_/Q _2107_/X _1967_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__a22o_1
X_3093_ _3350_/CLK _3093_/D vssd1 vssd1 vccd1 vccd1 _3093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2044_ _2044_/A vssd1 vssd1 vccd1 vccd1 _2044_/X sky130_fd_sc_hd__buf_2
X_2946_ input23/X input55/X input71/X input87/X _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2946_/X sky130_fd_sc_hd__mux4_1
X_2877_ _2873_/X _2874_/X _2875_/X _2876_/X _2660_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2877_/X sky130_fd_sc_hd__mux4_1
X_1828_ _2543_/A _1828_/B vssd1 vssd1 vccd1 vccd1 _1837_/A sky130_fd_sc_hd__or2_2
X_1759_ _1815_/A _1847_/A _2342_/C vssd1 vssd1 vccd1 vccd1 _2542_/A sky130_fd_sc_hd__or3_4
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _3429_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2800_ _3087_/Q _3371_/Q _3039_/Q _3031_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2800_/X sky130_fd_sc_hd__mux4_1
X_2731_ _3321_/Q _3305_/Q _3169_/Q _3337_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2731_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2662_ _2662_/A0 _2662_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2662_/X sky130_fd_sc_hd__mux2_2
X_2593_ _2592_/X _2472_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__mux2_1
X_1613_ _1615_/A _2615_/X vssd1 vssd1 vccd1 vccd1 _3454_/D sky130_fd_sc_hd__and2_1
X_1544_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3214_ _3296_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145_ _3335_/CLK _3145_/D vssd1 vssd1 vccd1 vccd1 _3145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3076_ _3439_/CLK _3076_/D vssd1 vssd1 vccd1 vccd1 _3076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2027_ _3250_/Q _2020_/A _1944_/X _2021_/A vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2929_ _3178_/Q _3154_/Q _3130_/Q _3106_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2929_/X sky130_fd_sc_hd__mux4_2
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput8 io_adr_i[5] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _3142_/Q _3118_/Q _3190_/Q _3438_/Q _2716_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2714_/X sky130_fd_sc_hd__mux4_2
X_2645_ _2877_/X _2644_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput301 _2542_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_10 sky130_fd_sc_hd__clkbuf_2
Xoutput334 _3479_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput323 _2565_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[7] sky130_fd_sc_hd__clkbuf_2
Xoutput312 _2569_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[11] sky130_fd_sc_hd__clkbuf_2
X_2576_ _2576_/A0 _2576_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__mux2_1
Xoutput345 _3489_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput356 _3464_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput367 _3507_/Q vssd1 vssd1 vccd1 vccd1 io_vout[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE3_7 _3484_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1527_ _1523_/X _3507_/Q _1524_/X _2712_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _3507_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3128_ _3447_/CLK _3128_/D vssd1 vssd1 vccd1 vccd1 _3128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3059_ _3367_/CLK _3059_/D vssd1 vssd1 vccd1 vccd1 _3059_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2430_ _2430_/A _2601_/X vssd1 vssd1 vccd1 vccd1 _2430_/X sky130_fd_sc_hd__and2_1
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2361_ _3045_/Q _2358_/X _2340_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _3045_/D sky130_fd_sc_hd__a22o_1
X_2292_ _2292_/A vssd1 vssd1 vccd1 vccd1 _2292_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_59_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2628_ _2628_/A0 _2628_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2628_/X sky130_fd_sc_hd__mux2_2
XFILLER_87_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2559_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1930_ _3308_/Q _1922_/X _1929_/X _1924_/X vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1861_ _3353_/Q _1857_/X _1652_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__a22o_1
Xinput22 io_b_dat_o_0[3] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_1
Xinput11 io_adr_i[8] vssd1 vssd1 vccd1 vccd1 _2683_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 io_b_dat_o_10[13] vssd1 vssd1 vccd1 vccd1 _2499_/B sky130_fd_sc_hd__clkbuf_1
Xinput44 io_b_dat_o_10[9] vssd1 vssd1 vccd1 vccd1 _2472_/B sky130_fd_sc_hd__clkbuf_1
Xinput55 io_b_dat_o_1[4] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
X_1792_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2098_/A sky130_fd_sc_hd__inv_2
Xinput66 io_b_dat_o_2[14] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
Xinput88 io_b_dat_o_3[5] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput77 io_b_dat_o_3[0] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
Xinput99 io_b_dat_o_4[15] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_1
X_3462_ _3493_/CLK _3462_/D vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfxtp_1
X_2413_ _3003_/Q _2407_/X _1941_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _3003_/D sky130_fd_sc_hd__a22o_1
X_3393_ _3423_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
X_2344_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2359_/A sky130_fd_sc_hd__inv_2
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2275_ _2282_/A vssd1 vssd1 vccd1 vccd1 _2275_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3438_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2060_ _3234_/Q _2052_/X _1953_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _3234_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2962_ _3163_/Q _3331_/Q _3315_/Q _3299_/Q _1700_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2962_/X sky130_fd_sc_hd__mux4_2
X_1913_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2893_ _2889_/X _2890_/X _2891_/X _2892_/X _2901_/S0 _2997_/S1 vssd1 vssd1 vccd1
+ vccd1 _2893_/X sky130_fd_sc_hd__mux4_1
X_1844_ _3362_/Q _1837_/A _1824_/X _1838_/A vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__a22o_1
X_1775_ _3395_/Q _1769_/X _1774_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__a22o_1
X_3514_ _3514_/CLK _3514_/D vssd1 vssd1 vccd1 vccd1 _3514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3445_ _3445_/CLK _3445_/D vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3376_ _3420_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2327_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2258_ _2258_/A vssd1 vssd1 vccd1 vccd1 _2258_/X sky130_fd_sc_hd__clkbuf_2
X_2189_ _3153_/Q _2181_/A _2150_/X _2182_/A vssd1 vssd1 vccd1 vccd1 _3153_/D sky130_fd_sc_hd__a22o_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput201 io_dat_i[1] vssd1 vssd1 vccd1 vccd1 _2559_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput223 io_dataLastBlock[10] vssd1 vssd1 vccd1 vccd1 _2644_/A0 sky130_fd_sc_hd__buf_1
Xinput212 io_dat_i[2] vssd1 vssd1 vccd1 vccd1 _2560_/A sky130_fd_sc_hd__buf_2
Xinput234 io_dataLastBlock[20] vssd1 vssd1 vccd1 vccd1 _2632_/A0 sky130_fd_sc_hd__buf_1
Xinput245 io_dataLastBlock[30] vssd1 vssd1 vccd1 vccd1 _2622_/A0 sky130_fd_sc_hd__buf_1
Xinput278 io_dataLastBlock[60] vssd1 vssd1 vccd1 vccd1 _2624_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput267 io_dataLastBlock[50] vssd1 vssd1 vccd1 vccd1 _2634_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput256 io_dataLastBlock[40] vssd1 vssd1 vccd1 vccd1 _2650_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput289 io_dsi_in[3] vssd1 vssd1 vccd1 vccd1 _2461_/B2 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1560_ _2669_/S vssd1 vssd1 vccd1 vccd1 _2520_/A sky130_fd_sc_hd__buf_1
X_1491_ _3519_/Q _1484_/Y _1485_/Y _1484_/A _1508_/B vssd1 vssd1 vccd1 vccd1 _1491_/X
+ sky130_fd_sc_hd__o221a_1
X_3230_ _3279_/CLK _3230_/D vssd1 vssd1 vccd1 vccd1 _3230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3161_ _3433_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2112_ _3198_/Q _2107_/X _1965_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _3437_/CLK _3092_/D vssd1 vssd1 vccd1 vccd1 _3092_/Q sky130_fd_sc_hd__dfxtp_1
X_2043_ _3243_/Q _2040_/X _2041_/X _2042_/X vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2945_ _2941_/X _2942_/X _2943_/X _2944_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2945_/X sky130_fd_sc_hd__mux4_1
X_2876_ _3023_/Q _3015_/Q _3007_/Q _3279_/Q _2644_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2876_/X sky130_fd_sc_hd__mux4_1
X_1827_ _3373_/Q _1817_/X _1826_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__a22o_1
X_1758_ _3401_/Q _1752_/X _1730_/X _1754_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__a22o_1
X_1689_ _1689_/A _1689_/B vssd1 vssd1 vccd1 vccd1 _1789_/C sky130_fd_sc_hd__or2_1
X_3428_ _3493_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
X_3359_ _3447_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2730_ _3241_/Q _3217_/Q _3289_/Q _3265_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2730_/X sky130_fd_sc_hd__mux4_2
X_2661_ _3495_/Q _2927_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__mux2_1
X_1612_ _1615_/A _2614_/X vssd1 vssd1 vccd1 vccd1 _3455_/D sky130_fd_sc_hd__and2_1
X_2592_ _2592_/A0 _2592_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2592_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1543_ _2562_/A vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _3301_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3144_ _3439_/CLK _3144_/D vssd1 vssd1 vccd1 vccd1 _3144_/Q sky130_fd_sc_hd__dfxtp_1
X_3075_ _3335_/CLK _3075_/D vssd1 vssd1 vccd1 vccd1 _3075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2026_ _3251_/Q _2020_/X _1941_/X _2021_/X vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _3058_/Q _3250_/Q _3226_/Q _3202_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2928_/X sky130_fd_sc_hd__mux4_2
X_2859_ input17/X input49/X input65/X input81/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2859_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 io_adr_i[6] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2713_ _3046_/Q _3350_/Q _3094_/Q _3070_/Q _2716_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2713_/X sky130_fd_sc_hd__mux4_2
X_2644_ _2644_/A0 _2644_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__mux2_1
Xoutput335 _3480_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[17] sky130_fd_sc_hd__clkbuf_2
X_2575_ _2557_/A _2997_/S1 _2575_/S vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__mux2_2
Xoutput302 _2551_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_2 sky130_fd_sc_hd__clkbuf_2
Xoutput324 _2566_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[8] sky130_fd_sc_hd__clkbuf_2
Xoutput313 _2570_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[12] sky130_fd_sc_hd__clkbuf_2
Xoutput346 _3490_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput357 _3465_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[8] sky130_fd_sc_hd__clkbuf_2
X_1526_ _1523_/X _3508_/Q _1524_/X _2717_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _3508_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput368 _3508_/Q vssd1 vssd1 vccd1 vccd1 io_vout[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3127_ _3447_/CLK _3127_/D vssd1 vssd1 vccd1 vccd1 _3127_/Q sky130_fd_sc_hd__dfxtp_1
X_3058_ _3367_/CLK _3058_/D vssd1 vssd1 vccd1 vccd1 _3058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2009_ _3264_/Q _2004_/X _1939_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__a22o_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2360_ _3046_/Q _2358_/X _2338_/X _2359_/X vssd1 vssd1 vccd1 vccd1 _3046_/D sky130_fd_sc_hd__a22o_1
X_2291_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2627_ _2627_/A0 _2627_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2627_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3456_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2558_ _2558_/A vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__clkbuf_1
X_1509_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1610_/A sky130_fd_sc_hd__buf_4
X_2489_ _3391_/Q vssd1 vssd1 vccd1 vccd1 _2489_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1860_ _3354_/Q _1857_/X _1649_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__a22o_1
Xinput12 io_adr_i[9] vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__clkbuf_4
X_1791_ _2097_/A vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__clkbuf_2
Xinput34 io_b_dat_o_10[14] vssd1 vssd1 vccd1 vccd1 _2511_/B sky130_fd_sc_hd__clkbuf_1
Xinput23 io_b_dat_o_0[4] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput45 io_b_dat_o_1[0] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput67 io_b_dat_o_2[15] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
Xinput89 io_b_dat_o_3[6] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput56 io_b_dat_o_1[5] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput78 io_b_dat_o_3[10] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
X_3461_ _3485_/CLK _3461_/D vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2412_ _3004_/Q _2407_/X _1939_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _3004_/D sky130_fd_sc_hd__a22o_1
X_3392_ _3392_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
X_2343_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2343_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2274_ _3100_/Q _2267_/X _2232_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _3100_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1989_ _3278_/Q _1986_/X _1935_/X _1987_/X vssd1 vssd1 vccd1 vccd1 _3278_/D sky130_fd_sc_hd__a22o_1
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _2669_/X _2671_/X _2672_/X _2425_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2961_/X sky130_fd_sc_hd__mux4_2
X_1912_ _3319_/Q _1906_/X _1656_/X _1907_/X vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__a22o_1
X_2892_ _3021_/Q _3013_/Q _3005_/Q _3277_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2892_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1843_ _3363_/Q _1837_/X _1822_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__a22o_1
X_1774_ _2560_/A vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__clkbuf_2
X_3513_ _3514_/CLK _3513_/D vssd1 vssd1 vccd1 vccd1 _3513_/Q sky130_fd_sc_hd__dfxtp_1
X_3444_ _3444_/CLK _3444_/D vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3375_ _3420_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater410 _1676_/A vssd1 vssd1 vccd1 vccd1 _2996_/S0 sky130_fd_sc_hd__buf_8
X_2326_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2257_ _2257_/A vssd1 vssd1 vccd1 vccd1 _2257_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2188_ _3154_/Q _2181_/A _2148_/X _2182_/A vssd1 vssd1 vccd1 vccd1 _3154_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_43_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput202 io_dat_i[20] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_1
Xinput224 io_dataLastBlock[11] vssd1 vssd1 vccd1 vccd1 _2641_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput235 io_dataLastBlock[21] vssd1 vssd1 vccd1 vccd1 _2631_/A0 sky130_fd_sc_hd__buf_1
Xinput213 io_dat_i[30] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_1
Xinput279 io_dataLastBlock[61] vssd1 vssd1 vccd1 vccd1 _2623_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput268 io_dataLastBlock[51] vssd1 vssd1 vccd1 vccd1 _2633_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput246 io_dataLastBlock[31] vssd1 vssd1 vccd1 vccd1 _2621_/A0 sky130_fd_sc_hd__buf_1
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput257 io_dataLastBlock[41] vssd1 vssd1 vccd1 vccd1 _2647_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1490_ _1490_/A _1490_/B _1490_/C _1490_/D vssd1 vssd1 vccd1 vccd1 _1508_/B sky130_fd_sc_hd__or4_4
X_3160_ _3410_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_1
X_2111_ _3199_/Q _2107_/X _1963_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__a22o_1
X_3091_ _3392_/CLK _3091_/D vssd1 vssd1 vccd1 vccd1 _3091_/Q sky130_fd_sc_hd__dfxtp_1
X_2042_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2944_ _3017_/Q _3009_/Q _3001_/Q _3273_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2944_/X sky130_fd_sc_hd__mux4_1
X_2875_ _3087_/Q _3371_/Q _3039_/Q _3031_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2875_/X sky130_fd_sc_hd__mux4_1
X_1826_ _2558_/A vssd1 vssd1 vccd1 vccd1 _1826_/X sky130_fd_sc_hd__buf_2
X_1757_ _3402_/Q _1752_/X _1728_/X _1754_/X vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__a22o_1
X_1688_ _1798_/D vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__buf_1
X_3427_ _3493_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
X_3358_ _3506_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2309_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2309_/X sky130_fd_sc_hd__clkbuf_2
X_3289_ _3303_/CLK _3289_/D vssd1 vssd1 vccd1 vccd1 _3289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2660_ _2920_/X _2921_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__mux2_1
X_1611_ _1615_/A _2613_/X vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__and2_1
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2591_ _2590_/X _2479_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2591_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1542_ _1515_/A _1539_/X _1730_/A _1541_/X _1528_/X vssd1 vssd1 vccd1 vccd1 _3502_/D
+ sky130_fd_sc_hd__o221a_1
X_3212_ _3295_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3143_ _3439_/CLK _3143_/D vssd1 vssd1 vccd1 vccd1 _3143_/Q sky130_fd_sc_hd__dfxtp_1
X_3074_ _3335_/CLK _3074_/D vssd1 vssd1 vccd1 vccd1 _3074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _3252_/Q _2020_/X _1939_/X _2021_/X vssd1 vssd1 vccd1 vccd1 _3252_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2927_ _2923_/X _2924_/X _2925_/X _2926_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2927_/X sky130_fd_sc_hd__mux4_2
X_2858_ _2508_/X _2509_/X _2638_/X _2512_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2858_/X sky130_fd_sc_hd__mux4_2
X_1809_ _2136_/A vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__inv_2
X_2789_ _3289_/Q _3265_/Q _3241_/Q _3217_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2789_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2708_/X _2709_/X _2710_/X _2711_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2712_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2643_ _2870_/X _2871_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2643_/X sky130_fd_sc_hd__mux2_1
X_2574_ _2574_/A vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__clkbuf_1
Xoutput303 _2550_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_3 sky130_fd_sc_hd__clkbuf_2
Xoutput325 _2567_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[9] sky130_fd_sc_hd__clkbuf_2
Xoutput314 _2571_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[13] sky130_fd_sc_hd__clkbuf_2
Xoutput347 _3491_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput336 _3481_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput358 _3466_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[9] sky130_fd_sc_hd__clkbuf_2
X_1525_ _1523_/X _3509_/Q _1524_/X _2722_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _3509_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput369 _3509_/Q vssd1 vssd1 vccd1 vccd1 io_vout[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3126_ _3506_/CLK _3126_/D vssd1 vssd1 vccd1 vccd1 _3126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3057_ _3372_/CLK _3057_/D vssd1 vssd1 vccd1 vccd1 _3057_/Q sky130_fd_sc_hd__dfxtp_1
X_2008_ _3265_/Q _2004_/X _1937_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__a22o_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2290_ _3088_/Q _1703_/X _2232_/X _1705_/X vssd1 vssd1 vccd1 vccd1 _3088_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2626_ _2626_/A0 _2626_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2626_/X sky130_fd_sc_hd__mux2_2
X_2557_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__clkbuf_1
X_2488_ _2523_/A _2589_/X vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__and2_1
XFILLER_87_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1508_ _3516_/Q _1508_/B vssd1 vssd1 vccd1 vccd1 _1508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3109_ _3109_/CLK _3109_/D vssd1 vssd1 vccd1 vccd1 _3109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 io_b_dat_o_0[0] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
X_1790_ _1816_/A _2550_/A vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__or2_4
Xinput35 io_b_dat_o_10[15] vssd1 vssd1 vccd1 vccd1 _2522_/B sky130_fd_sc_hd__clkbuf_1
Xinput46 io_b_dat_o_1[10] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
Xinput24 io_b_dat_o_0[5] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput79 io_b_dat_o_3[11] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_1
Xinput57 io_b_dat_o_1[6] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 io_b_dat_o_2[1] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_3460_ _3485_/CLK _3460_/D vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfxtp_1
X_2411_ _3005_/Q _2407_/X _2046_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _3005_/D sky130_fd_sc_hd__a22o_1
X_3391_ _3423_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2342_ _2342_/A _2342_/B _2342_/C _2342_/D vssd1 vssd1 vccd1 vccd1 _2358_/A sky130_fd_sc_hd__or4_4
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2273_ _3101_/Q _2267_/X _2162_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _3101_/D sky130_fd_sc_hd__a22o_1
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1988_ _3279_/Q _1986_/X _1932_/X _1987_/X vssd1 vssd1 vccd1 vccd1 _3279_/D sky130_fd_sc_hd__a22o_1
X_2609_ _2608_/X _2419_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2960_ _2960_/A0 _2960_/A1 _2960_/A2 _2960_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2960_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1911_ _3320_/Q _1906_/X _1654_/X _1907_/X vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2891_ _3085_/Q _3369_/Q _3037_/Q _3029_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2891_/X sky130_fd_sc_hd__mux4_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1842_ _3364_/Q _1837_/X _1818_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__a22o_1
X_1773_ _3396_/Q _1769_/X _1770_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__a22o_1
X_3512_ _3515_/CLK _3512_/D vssd1 vssd1 vccd1 vccd1 _3512_/Q sky130_fd_sc_hd__dfxtp_1
X_3443_ _3443_/CLK _3443_/D vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3374_ _3420_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater411 _1700_/A vssd1 vssd1 vccd1 vccd1 _1676_/A sky130_fd_sc_hd__buf_4
X_2325_ _3064_/Q _1712_/X _2324_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _3064_/D sky130_fd_sc_hd__a22o_1
Xrepeater400 _2644_/S vssd1 vssd1 vccd1 vccd1 _2682_/S sky130_fd_sc_hd__buf_8
X_2256_ _3112_/Q _1693_/X _2232_/X _1695_/X vssd1 vssd1 vccd1 vccd1 _3112_/D sky130_fd_sc_hd__a22o_1
X_2187_ _3155_/Q _2181_/X _2146_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _3155_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3429_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput225 io_dataLastBlock[12] vssd1 vssd1 vccd1 vccd1 _2587_/A0 sky130_fd_sc_hd__buf_1
Xinput236 io_dataLastBlock[22] vssd1 vssd1 vccd1 vccd1 _2630_/A0 sky130_fd_sc_hd__buf_1
Xinput203 io_dat_i[21] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__buf_1
Xinput214 io_dat_i[31] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__buf_1
Xinput269 io_dataLastBlock[52] vssd1 vssd1 vccd1 vccd1 _2632_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput258 io_dataLastBlock[42] vssd1 vssd1 vccd1 vccd1 _2644_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput247 io_dataLastBlock[32] vssd1 vssd1 vccd1 vccd1 _2682_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2110_ _3200_/Q _2107_/X _1959_/X _2109_/X vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__a22o_1
X_3090_ _3346_/CLK _3090_/D vssd1 vssd1 vccd1 vccd1 _3090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2041_ _2041_/A vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2943_ _3081_/Q _3365_/Q _3033_/Q _3025_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2943_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2874_ _3183_/Q _3159_/Q _3135_/Q _3111_/Q _2644_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2874_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1825_ _3374_/Q _1817_/X _1824_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__a22o_1
X_1756_ _3403_/Q _1752_/X _1726_/X _1754_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1687_ _3429_/Q _1681_/X _1670_/X _1683_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__a22o_1
X_3426_ _3500_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
X_3357_ _3444_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
X_2308_ _3076_/Q _2301_/X _2232_/X _2303_/X vssd1 vssd1 vccd1 vccd1 _3076_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3288_ _3307_/CLK _3288_/D vssd1 vssd1 vccd1 vccd1 _3288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2239_ _3122_/Q _2234_/X _2238_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _3122_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1610_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1615_/A sky130_fd_sc_hd__buf_1
XFILLER_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2590_ _2590_/A0 _2590_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1541_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__buf_2
XFILLER_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3211_ _3295_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_1
X_3142_ _3433_/CLK _3142_/D vssd1 vssd1 vccd1 vccd1 _3142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3073_ _3335_/CLK _3073_/D vssd1 vssd1 vccd1 vccd1 _3073_/Q sky130_fd_sc_hd__dfxtp_1
X_2024_ _3253_/Q _2020_/X _1937_/X _2021_/X vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__a22o_1
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2926_ _3094_/Q _3070_/Q _3046_/Q _3350_/Q _1700_/A _2991_/S1 vssd1 vssd1 vccd1 vccd1
+ _2926_/X sky130_fd_sc_hd__mux4_2
X_2857_ input98/X _2857_/A1 _2857_/A2 _2857_/A3 _2632_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2857_/X sky130_fd_sc_hd__mux4_1
X_1808_ _2136_/A vssd1 vssd1 vccd1 vccd1 _1808_/X sky130_fd_sc_hd__clkbuf_2
X_2788_ _3169_/Q _3337_/Q _3321_/Q _3305_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2788_/X sky130_fd_sc_hd__mux4_1
X_1739_ _3412_/Q _1736_/X _1722_/X _1738_/X vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3409_ _3409_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _3317_/Q _3301_/Q _3165_/Q _3333_/Q _2716_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2711_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2642_ _2869_/X _2641_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__mux2_1
X_2573_ _2573_/A vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__clkbuf_1
Xoutput326 _2574_/X vssd1 vssd1 vccd1 vccd1 io_b_we_i sky130_fd_sc_hd__clkbuf_2
Xoutput304 _2549_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_4 sky130_fd_sc_hd__clkbuf_2
Xoutput315 _2572_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[14] sky130_fd_sc_hd__clkbuf_2
Xoutput348 _3492_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput337 _3482_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[19] sky130_fd_sc_hd__clkbuf_2
X_1524_ _1524_/A vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__buf_1
Xoutput359 _2466_/X vssd1 vssd1 vccd1 vccd1 io_dsi_o sky130_fd_sc_hd__clkbuf_2
XFILLER_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3445_/CLK _3125_/D vssd1 vssd1 vccd1 vccd1 _3125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3056_ _3444_/CLK _3056_/D vssd1 vssd1 vccd1 vccd1 _3056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2007_ _3266_/Q _2004_/X _1935_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2909_ _2653_/X _2655_/X _2656_/X _2447_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2909_/X sky130_fd_sc_hd__mux4_2
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2625_ _2625_/A0 _2625_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__mux2_2
X_2556_ _2683_/S vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__clkbuf_1
X_2487_ _2487_/A vssd1 vssd1 vccd1 vccd1 _2523_/A sky130_fd_sc_hd__buf_1
XFILLER_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1507_ _2687_/S _1506_/X _3517_/Q _1502_/Y _1618_/A vssd1 vssd1 vccd1 vccd1 _3517_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3108_ _3180_/CLK _3108_/D vssd1 vssd1 vccd1 vccd1 _3108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3039_ _3277_/CLK _3039_/D vssd1 vssd1 vccd1 vccd1 _3039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3443_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_b_dat_o_0[10] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 io_b_dat_o_0[6] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 io_b_dat_o_10[1] vssd1 vssd1 vccd1 vccd1 _2419_/B sky130_fd_sc_hd__clkbuf_1
Xinput47 io_b_dat_o_1[11] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 io_b_dat_o_1[7] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_1
Xinput69 io_b_dat_o_2[2] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
X_2410_ _3006_/Q _2407_/X _2044_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _3006_/D sky130_fd_sc_hd__a22o_1
X_3390_ _3420_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2341_ _3057_/Q _2326_/A _2340_/X _2328_/A vssd1 vssd1 vccd1 vccd1 _3057_/D sky130_fd_sc_hd__a22o_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2272_ _3102_/Q _2267_/X _2160_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _3102_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1987_ _1987_/A vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__clkbuf_2
X_2608_ _2608_/A0 _2608_/A1 _2610_/S vssd1 vssd1 vccd1 vccd1 _2608_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2539_ _3456_/Q _2537_/Y _2620_/S vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2890_ _3181_/Q _3157_/Q _3133_/Q _3109_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2890_/X sky130_fd_sc_hd__mux4_2
X_1910_ _3321_/Q _1906_/X _1652_/X _1907_/X vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__a22o_1
XFILLER_42_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1841_ _3365_/Q _1837_/X _1662_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__a22o_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1772_ _2378_/A vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__clkbuf_2
X_3511_ _3514_/CLK _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/Q sky130_fd_sc_hd__dfxtp_1
X_3442_ _3443_/CLK _3442_/D vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfxtp_1
X_3373_ _3420_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_1
X_2324_ _2569_/A vssd1 vssd1 vccd1 vccd1 _2324_/X sky130_fd_sc_hd__buf_2
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater401 _2785_/S0 vssd1 vssd1 vccd1 vccd1 _2910_/S0 sky130_fd_sc_hd__buf_8
XFILLER_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater412 input5/X vssd1 vssd1 vccd1 vccd1 _1700_/A sky130_fd_sc_hd__buf_8
X_2255_ _3113_/Q _2246_/A _2132_/X _2248_/A vssd1 vssd1 vccd1 vccd1 _3113_/D sky130_fd_sc_hd__a22o_1
X_2186_ _3156_/Q _2181_/X _2144_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput226 io_dataLastBlock[13] vssd1 vssd1 vccd1 vccd1 _2584_/A0 sky130_fd_sc_hd__buf_1
Xinput215 io_dat_i[3] vssd1 vssd1 vccd1 vccd1 _2561_/A sky130_fd_sc_hd__buf_2
Xinput204 io_dat_i[22] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__buf_1
Xinput259 io_dataLastBlock[43] vssd1 vssd1 vccd1 vccd1 _2641_/A1 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3504_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput237 io_dataLastBlock[23] vssd1 vssd1 vccd1 vccd1 _2629_/A0 sky130_fd_sc_hd__buf_1
Xinput248 io_dataLastBlock[33] vssd1 vssd1 vccd1 vccd1 _2678_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2040_ _2052_/A vssd1 vssd1 vccd1 vccd1 _2040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _3177_/Q _3153_/Q _3129_/Q _3105_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2942_/X sky130_fd_sc_hd__mux4_2
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2873_ _3063_/Q _3255_/Q _3231_/Q _3207_/Q _2682_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2873_/X sky130_fd_sc_hd__mux4_2
X_1824_ _2559_/A vssd1 vssd1 vccd1 vccd1 _1824_/X sky130_fd_sc_hd__buf_2
X_1755_ _3404_/Q _1752_/X _1722_/X _1754_/X vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__a22o_1
X_1686_ _3430_/Q _1681_/X _1668_/X _1683_/X vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__a22o_1
X_3425_ _3429_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _3439_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2307_ _3077_/Q _2301_/X _2162_/X _2303_/X vssd1 vssd1 vccd1 vccd1 _3077_/D sky130_fd_sc_hd__a22o_1
X_3287_ _3303_/CLK _3287_/D vssd1 vssd1 vccd1 vccd1 _3287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2238_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2238_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2169_ _3169_/Q _2165_/X _2142_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1540_ _2558_/A vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__clkbuf_2
X_3210_ _3474_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3141_ _3438_/CLK _3141_/D vssd1 vssd1 vccd1 vccd1 _3141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _3351_/CLK _3072_/D vssd1 vssd1 vccd1 vccd1 _3072_/Q sky130_fd_sc_hd__dfxtp_1
X_2023_ _3254_/Q _2020_/X _1935_/X _2021_/X vssd1 vssd1 vccd1 vccd1 _3254_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2925_ _3190_/Q _3438_/Q _3142_/Q _3118_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2925_/X sky130_fd_sc_hd__mux4_1
X_2856_ input18/X input50/X input66/X input82/X _2632_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2856_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1807_ _1816_/A _2549_/A vssd1 vssd1 vccd1 vccd1 _2136_/A sky130_fd_sc_hd__or2_4
X_2787_ _2783_/X _2784_/X _2785_/X _2786_/X _2901_/S0 _2997_/S1 vssd1 vssd1 vccd1
+ vccd1 _2787_/X sky130_fd_sc_hd__mux4_2
X_1738_ _2408_/A vssd1 vssd1 vccd1 vccd1 _1738_/X sky130_fd_sc_hd__clkbuf_2
X_1669_ _3434_/Q _1658_/X _1668_/X _1660_/X vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__a22o_1
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3408_ _3409_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3339_ _3443_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2710_ _3237_/Q _3213_/Q _3285_/Q _3261_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2710_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2641_ _2641_/A0 _2641_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__mux2_1
Xoutput305 _2548_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_5 sky130_fd_sc_hd__clkbuf_2
Xoutput316 _2573_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[15] sky130_fd_sc_hd__clkbuf_2
X_2572_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1523_ _3502_/Q vssd1 vssd1 vccd1 vccd1 _1523_/X sky130_fd_sc_hd__buf_1
Xoutput327 _3457_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput349 _3459_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput338 _3458_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3124_ _3336_/CLK _3124_/D vssd1 vssd1 vccd1 vccd1 _3124_/Q sky130_fd_sc_hd__dfxtp_1
X_3055_ _3444_/CLK _3055_/D vssd1 vssd1 vccd1 vccd1 _3055_/Q sky130_fd_sc_hd__dfxtp_1
X_2006_ _3267_/Q _2004_/X _1932_/X _2005_/X vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__a22o_1
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2908_ _2908_/A0 _2908_/A1 _2908_/A2 _2908_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2908_/X sky130_fd_sc_hd__mux4_1
X_2839_ _2483_/Y _2482_/Y _2495_/Y _2478_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2839_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_7_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3398_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2624_ _2624_/A0 _2624_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2624_/X sky130_fd_sc_hd__mux2_2
X_2555_ _1491_/X _2687_/S _3519_/Q _1502_/Y _1592_/A vssd1 vssd1 vccd1 vccd1 _3519_/D
+ sky130_fd_sc_hd__o221a_1
X_2486_ _2522_/A _2486_/B vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__and2_1
X_1506_ _1482_/A _1482_/B _3517_/Q _3516_/Q _1508_/B vssd1 vssd1 vccd1 vccd1 _1506_/X
+ sky130_fd_sc_hd__o221a_1
X_3107_ _3180_/CLK _3107_/D vssd1 vssd1 vccd1 vccd1 _3107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3038_ _3087_/CLK _3038_/D vssd1 vssd1 vccd1 vccd1 _3038_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 io_b_dat_o_0[11] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput26 io_b_dat_o_0[7] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
Xinput37 io_b_dat_o_10[2] vssd1 vssd1 vccd1 vccd1 _2416_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput48 io_b_dat_o_1[12] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput59 io_b_dat_o_1[8] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2340_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__clkbuf_2
X_2271_ _3103_/Q _2267_/X _2158_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _3103_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1986_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1986_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2607_ _2606_/X _2416_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2607_/X sky130_fd_sc_hd__mux2_1
X_2538_ _2537_/A _2537_/B _2537_/Y vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2469_ _3375_/Q vssd1 vssd1 vccd1 vccd1 _2469_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1840_ _3366_/Q _1837_/X _1659_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__a22o_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3510_ _3514_/CLK _3510_/D vssd1 vssd1 vccd1 vccd1 _3510_/Q sky130_fd_sc_hd__dfxtp_1
X_1771_ _2377_/A vssd1 vssd1 vccd1 vccd1 _2378_/A sky130_fd_sc_hd__inv_2
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _3443_/CLK _3441_/D vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfxtp_1
X_3372_ _3372_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2323_ _3065_/Q _2316_/A _1730_/A _2317_/A vssd1 vssd1 vccd1 vccd1 _3065_/D sky130_fd_sc_hd__a22o_1
Xrepeater402 _2913_/S0 vssd1 vssd1 vccd1 vccd1 _2785_/S0 sky130_fd_sc_hd__buf_6
Xrepeater413 input2/X vssd1 vssd1 vccd1 vccd1 _2575_/S sky130_fd_sc_hd__buf_8
X_2254_ _3114_/Q _2246_/X _2130_/X _2248_/X vssd1 vssd1 vccd1 vccd1 _3114_/D sky130_fd_sc_hd__a22o_1
X_2185_ _3157_/Q _2181_/X _2142_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _3157_/D sky130_fd_sc_hd__a22o_1
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1969_ _3292_/Q _1958_/X _1929_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput227 io_dataLastBlock[14] vssd1 vssd1 vccd1 vccd1 _2581_/A0 sky130_fd_sc_hd__buf_1
Xinput216 io_dat_i[4] vssd1 vssd1 vccd1 vccd1 _2562_/A sky130_fd_sc_hd__clkbuf_4
Xinput205 io_dat_i[23] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__buf_1
Xinput238 io_dataLastBlock[24] vssd1 vssd1 vccd1 vccd1 _2628_/A0 sky130_fd_sc_hd__buf_1
Xinput249 io_dataLastBlock[34] vssd1 vssd1 vccd1 vccd1 _2674_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3367_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _3057_/Q _3249_/Q _3225_/Q _3201_/Q _2982_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2941_/X sky130_fd_sc_hd__mux4_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2872_ _2481_/X _2642_/X _2643_/X _2488_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2872_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1823_ _3375_/Q _1817_/X _1822_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__a22o_1
X_1754_ _2398_/A vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1685_ _3431_/Q _1681_/X _1666_/X _1683_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__a22o_1
X_3424_ _3424_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
X_3355_ _3355_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3286_ _3296_/CLK _3286_/D vssd1 vssd1 vccd1 vccd1 _3286_/Q sky130_fd_sc_hd__dfxtp_1
X_2306_ _3078_/Q _2301_/X _2160_/X _2303_/X vssd1 vssd1 vccd1 vccd1 _3078_/D sky130_fd_sc_hd__a22o_1
X_2237_ _3123_/Q _2234_/X _2235_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _3123_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _3170_/Q _2165_/X _2140_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2099_ _3207_/Q _2097_/X _2041_/X _2098_/X vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__a22o_1
XFILLER_70_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3140_ _3333_/CLK _3140_/D vssd1 vssd1 vccd1 vccd1 _3140_/Q sky130_fd_sc_hd__dfxtp_1
X_3071_ _3502_/CLK _3071_/D vssd1 vssd1 vccd1 vccd1 _3071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2022_ _3255_/Q _2020_/X _1932_/X _2021_/X vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__a22o_1
X_2924_ _3286_/Q _3262_/Q _3238_/Q _3214_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2924_/X sky130_fd_sc_hd__mux4_2
X_2855_ _2519_/X _2520_/X _2637_/X _2523_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2855_/X sky130_fd_sc_hd__mux4_2
X_1806_ _1806_/A input8/X _2266_/C vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__or3_4
X_2786_ _3098_/Q _3074_/Q _3050_/Q _3354_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2786_/X sky130_fd_sc_hd__mux4_2
X_1737_ _2407_/A vssd1 vssd1 vccd1 vccd1 _2408_/A sky130_fd_sc_hd__inv_2
X_1668_ _1728_/A vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__buf_2
X_3407_ _3409_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
X_1599_ _1603_/A _2888_/X vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__and2_1
X_3338_ _3445_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3269_ _3294_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ _2862_/X _2863_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2640_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput306 _2546_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_6 sky130_fd_sc_hd__clkbuf_2
Xoutput317 _2559_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[1] sky130_fd_sc_hd__clkbuf_2
X_2571_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2571_/X sky130_fd_sc_hd__clkbuf_1
Xoutput339 _3483_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput328 _3467_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[10] sky130_fd_sc_hd__clkbuf_2
X_1522_ _1515_/X _3510_/Q _1516_/X _2727_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _3510_/D
+ sky130_fd_sc_hd__o221a_1
X_3123_ _3335_/CLK _3123_/D vssd1 vssd1 vccd1 vccd1 _3123_/Q sky130_fd_sc_hd__dfxtp_1
X_3054_ _3336_/CLK _3054_/D vssd1 vssd1 vccd1 vccd1 _3054_/Q sky130_fd_sc_hd__dfxtp_1
X_2005_ _2012_/A vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2907_ input26/X input58/X input74/X input90/X _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2907_/X sky130_fd_sc_hd__mux4_1
X_2838_ _2470_/Y _2469_/Y _2489_/Y _2477_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2838_/X sky130_fd_sc_hd__mux4_2
X_2769_ _3293_/Q _3269_/Q _3245_/Q _3221_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2769_/X sky130_fd_sc_hd__mux4_2
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2623_ _2623_/A0 _2623_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__mux2_2
X_2554_ _2554_/A _3473_/Q vssd1 vssd1 vccd1 vccd1 _2554_/Y sky130_fd_sc_hd__nor2_1
X_1505_ _2687_/S _1501_/X _3518_/Q _1502_/Y _1618_/A vssd1 vssd1 vccd1 vccd1 _3518_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2485_ _2485_/A vssd1 vssd1 vccd1 vccd1 _2522_/A sky130_fd_sc_hd__buf_1
X_3106_ _3497_/CLK _3106_/D vssd1 vssd1 vccd1 vccd1 _3106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3037_ _3353_/CLK _3037_/D vssd1 vssd1 vccd1 vccd1 _3037_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_46_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput16 io_b_dat_o_0[12] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput27 io_b_dat_o_0[8] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
Xinput49 io_b_dat_o_1[13] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 io_b_dat_o_10[3] vssd1 vssd1 vccd1 vccd1 _2424_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2270_ _3104_/Q _2267_/X _2154_/X _2269_/X vssd1 vssd1 vccd1 vccd1 _3104_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1985_ _3280_/Q _1799_/X _1929_/X _1801_/X vssd1 vssd1 vccd1 vccd1 _3280_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2606_ _2606_/A0 _2606_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2606_/X sky130_fd_sc_hd__mux2_1
X_2537_ _2537_/A _2537_/B vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2468_ _3394_/Q vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__inv_2
X_2399_ _3015_/Q _2397_/X _2041_/A _2398_/X vssd1 vssd1 vccd1 vccd1 _3015_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _2561_/A vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _3504_/CLK _3440_/D vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfxtp_1
X_3371_ _3371_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2322_ _3066_/Q _2316_/X _1728_/A _2317_/X vssd1 vssd1 vccd1 vccd1 _3066_/D sky130_fd_sc_hd__a22o_1
XFILLER_85_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater414 _2683_/S vssd1 vssd1 vccd1 vccd1 _2669_/S sky130_fd_sc_hd__buf_8
X_2253_ _3115_/Q _2246_/X _2128_/X _2248_/X vssd1 vssd1 vccd1 vccd1 _3115_/D sky130_fd_sc_hd__a22o_1
Xrepeater403 _2918_/S0 vssd1 vssd1 vccd1 vccd1 _2913_/S0 sky130_fd_sc_hd__buf_8
X_2184_ _3158_/Q _2181_/X _2140_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1968_ _3293_/Q _1958_/X _1967_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _3293_/D sky130_fd_sc_hd__a22o_1
X_1899_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1914_/A sky130_fd_sc_hd__inv_2
XFILLER_88_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput217 io_dat_i[5] vssd1 vssd1 vccd1 vccd1 _2563_/A sky130_fd_sc_hd__clkbuf_4
Xinput206 io_dat_i[24] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__buf_1
XFILLER_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput228 io_dataLastBlock[15] vssd1 vssd1 vccd1 vccd1 _2578_/A0 sky130_fd_sc_hd__buf_1
Xinput239 io_dataLastBlock[25] vssd1 vssd1 vccd1 vccd1 _2627_/A0 sky130_fd_sc_hd__buf_1
XFILLER_84_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3295_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2940_ _2936_/X _2937_/X _2938_/X _2939_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2940_/X sky130_fd_sc_hd__mux4_2
X_2871_ input95/X _2871_/A1 _2871_/A2 _2871_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2871_/X sky130_fd_sc_hd__mux4_1
X_1822_ _2560_/A vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__clkbuf_2
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1753_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2398_/A sky130_fd_sc_hd__inv_2
X_1684_ _3432_/Q _1681_/X _1664_/X _1683_/X vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3423_ _3423_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
X_3354_ _3443_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2305_ _3079_/Q _2301_/X _2158_/X _2303_/X vssd1 vssd1 vccd1 vccd1 _3079_/D sky130_fd_sc_hd__a22o_1
X_3285_ _3301_/CLK _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2236_ _2248_/A vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2167_ _3171_/Q _2165_/X _2137_/X _2166_/X vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2098_ _2098_/A vssd1 vssd1 vccd1 vccd1 _2098_/X sky130_fd_sc_hd__buf_2
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ _3350_/CLK _3070_/D vssd1 vssd1 vccd1 vccd1 _3070_/Q sky130_fd_sc_hd__dfxtp_1
X_2021_ _2021_/A vssd1 vssd1 vccd1 vccd1 _2021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2923_ _3166_/Q _3334_/Q _3318_/Q _3302_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2923_/X sky130_fd_sc_hd__mux4_2
X_2854_ input99/X _2854_/A1 _2854_/A2 _2854_/A3 _2632_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2854_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1805_ _3381_/Q _1799_/X _1778_/X _1801_/X vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__a22o_1
X_2785_ _3194_/Q _3442_/Q _3146_/Q _3122_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2785_/X sky130_fd_sc_hd__mux4_1
X_1736_ _2407_/A vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1667_ _3435_/Q _1658_/X _1666_/X _1660_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__a22o_1
X_1598_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1603_/A sky130_fd_sc_hd__buf_1
X_3406_ _3424_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3337_ _3443_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3268_ _3297_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2219_ _3133_/Q _2215_/X _2142_/X _2216_/X vssd1 vssd1 vccd1 vccd1 _3133_/D sky130_fd_sc_hd__a22o_1
X_3199_ _3448_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput307 _2545_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_7 sky130_fd_sc_hd__clkbuf_2
X_2570_ _2570_/A vssd1 vssd1 vccd1 vccd1 _2570_/X sky130_fd_sc_hd__clkbuf_1
Xoutput329 _3468_/Q vssd1 vssd1 vccd1 vccd1 io_dat_o[11] sky130_fd_sc_hd__clkbuf_2
X_1521_ _1515_/X _3511_/Q _1516_/X _2732_/X _1520_/X vssd1 vssd1 vccd1 vccd1 _3511_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput318 _2560_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3335_/CLK _3122_/D vssd1 vssd1 vccd1 vccd1 _3122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3053_ _3336_/CLK _3053_/D vssd1 vssd1 vccd1 vccd1 _3053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2004_ _2011_/A vssd1 vssd1 vccd1 vccd1 _2004_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2906_ _2902_/X _2903_/X _2904_/X _2905_/X _2660_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2906_/X sky130_fd_sc_hd__mux4_1
X_2837_ _2833_/X _2834_/X _2835_/X _2836_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2837_/X sky130_fd_sc_hd__mux4_2
X_2768_ _3173_/Q _3341_/Q _3325_/Q _3309_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2768_/X sky130_fd_sc_hd__mux4_2
X_2699_ _3139_/Q _3115_/Q _3187_/Q _3435_/Q _2852_/X _2716_/S1 vssd1 vssd1 vccd1 vccd1
+ _2699_/X sky130_fd_sc_hd__mux4_2
X_1719_ _1806_/A _1780_/B _2300_/C vssd1 vssd1 vccd1 vccd1 _2548_/A sky130_fd_sc_hd__or3_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2622_ _2622_/A0 _2622_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2622_/X sky130_fd_sc_hd__mux2_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2553_ _2553_/A _2553_/B vssd1 vssd1 vccd1 vccd1 _2553_/Y sky130_fd_sc_hd__nor2_2
X_1504_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1618_/A sky130_fd_sc_hd__buf_1
X_2484_ _3403_/Q vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3105_ _3501_/CLK _3105_/D vssd1 vssd1 vccd1 vccd1 _3105_/Q sky130_fd_sc_hd__dfxtp_1
X_3036_ _3087_/CLK _3036_/D vssd1 vssd1 vccd1 vccd1 _3036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3493_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 io_b_dat_o_0[13] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 io_b_dat_o_0[9] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 io_b_dat_o_10[4] vssd1 vssd1 vccd1 vccd1 _2426_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1984_ _3281_/Q _1977_/A _1955_/X _1978_/A vssd1 vssd1 vccd1 vccd1 _3281_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2605_ _2604_/X _2424_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2536_ _3455_/Q vssd1 vssd1 vccd1 vccd1 _2537_/A sky130_fd_sc_hd__inv_2
X_2467_ _2490_/A _2787_/X vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__and2_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2398_ _2398_/A vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3019_ _3019_/CLK _3019_/D vssd1 vssd1 vccd1 vccd1 _3019_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ _3371_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_1
X_2321_ _3067_/Q _2316_/X _1726_/A _2317_/X vssd1 vssd1 vccd1 vccd1 _3067_/D sky130_fd_sc_hd__a22o_1
X_2252_ _3116_/Q _2246_/X _2126_/X _2248_/X vssd1 vssd1 vccd1 vccd1 _3116_/D sky130_fd_sc_hd__a22o_1
Xrepeater404 _2644_/S vssd1 vssd1 vccd1 vccd1 _2918_/S0 sky130_fd_sc_hd__buf_8
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2183_ _3159_/Q _2181_/X _2137_/X _2182_/X vssd1 vssd1 vccd1 vccd1 _3159_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _2570_/A vssd1 vssd1 vccd1 vccd1 _1967_/X sky130_fd_sc_hd__clkbuf_2
X_1898_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1898_/X sky130_fd_sc_hd__clkbuf_2
X_2519_ _2520_/A _2757_/X vssd1 vssd1 vccd1 vccd1 _2519_/X sky130_fd_sc_hd__and2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3499_ _3500_/CLK _3499_/D vssd1 vssd1 vccd1 vccd1 _3499_/Q sky130_fd_sc_hd__dfxtp_1
Xinput218 io_dat_i[6] vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__clkbuf_4
Xinput207 io_dat_i[25] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_1
XFILLER_88_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput229 io_dataLastBlock[16] vssd1 vssd1 vccd1 vccd1 _2636_/A0 sky130_fd_sc_hd__buf_1
XFILLER_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3277_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ input15/X input47/X input63/X input79/X _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2870_/X sky130_fd_sc_hd__mux4_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1821_ _3376_/Q _1817_/X _1818_/X _1820_/X vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__a22o_1
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ _2397_/A vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__clkbuf_2
X_1683_ _2216_/A vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__clkbuf_2
X_3422_ _3424_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
X_3353_ _3353_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
X_2304_ _3080_/Q _2301_/X _2154_/X _2303_/X vssd1 vssd1 vccd1 vccd1 _3080_/D sky130_fd_sc_hd__a22o_1
X_3284_ _3295_/CLK _3284_/D vssd1 vssd1 vccd1 vccd1 _3284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2235_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2235_/X sky130_fd_sc_hd__clkbuf_2
X_2166_ _2173_/A vssd1 vssd1 vccd1 vccd1 _2166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2097_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2097_/X sky130_fd_sc_hd__buf_2
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ input93/X _2999_/A1 _2999_/A2 _2999_/A3 _2610_/S _2611_/S vssd1 vssd1 vccd1
+ vccd1 _2999_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2020_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2922_ _2657_/X _2659_/X _2660_/X _2439_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2922_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2853_ input19/X input51/X input67/X input83/X _2632_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2853_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1804_ _3382_/Q _1799_/X _1776_/X _1801_/X vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__a22o_1
X_2784_ _3290_/Q _3266_/Q _3242_/Q _3218_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2784_/X sky130_fd_sc_hd__mux4_2
X_1735_ _2342_/A _1798_/B _2342_/C _1828_/B vssd1 vssd1 vccd1 vccd1 _2407_/A sky130_fd_sc_hd__or4_4
X_1666_ _1726_/A vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__buf_2
X_1597_ _1597_/A _2880_/X vssd1 vssd1 vccd1 vccd1 _3467_/D sky130_fd_sc_hd__and2_1
X_3405_ _3423_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_3336_ _3336_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3267_ _3303_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
X_2218_ _3134_/Q _2215_/X _2140_/X _2216_/X vssd1 vssd1 vccd1 vccd1 _3134_/D sky130_fd_sc_hd__a22o_1
X_3198_ _3294_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_1
X_2149_ _3178_/Q _2136_/A _2148_/X _2138_/A vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput308 _2544_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_8 sky130_fd_sc_hd__clkbuf_2
Xoutput319 _2561_/X vssd1 vssd1 vccd1 vccd1 io_b_dat_i[3] sky130_fd_sc_hd__clkbuf_2
X_1520_ _1610_/A vssd1 vssd1 vccd1 vccd1 _1520_/X sky130_fd_sc_hd__clkbuf_2
X_3121_ _3335_/CLK _3121_/D vssd1 vssd1 vccd1 vccd1 _3121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3052_ _3439_/CLK _3052_/D vssd1 vssd1 vccd1 vccd1 _3052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _3268_/Q _1996_/X _1929_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2905_ _3020_/Q _3012_/Q _3004_/Q _3276_/Q _2644_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2905_/X sky130_fd_sc_hd__mux4_1
X_2836_ _2501_/Y _2502_/Y _2504_/Y _2505_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2836_/X sky130_fd_sc_hd__mux4_2
X_2767_ _2763_/X _2764_/X _2765_/X _2766_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2767_/X sky130_fd_sc_hd__mux4_2
X_2698_ _3043_/Q _3347_/Q _3091_/Q _3067_/Q _2852_/X _2716_/S1 vssd1 vssd1 vccd1 vccd1
+ _2698_/X sky130_fd_sc_hd__mux4_2
X_1718_ _3417_/Q _1712_/X _1670_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__a22o_1
X_1649_ _2044_/A vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3319_ _3504_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2621_ _2621_/A0 _2621_/A1 _2632_/S vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__mux2_2
X_2552_ _2552_/A _2552_/B vssd1 vssd1 vccd1 vccd1 _2552_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1503_ _1590_/A vssd1 vssd1 vccd1 vccd1 _1555_/A sky130_fd_sc_hd__inv_2
X_2483_ _3379_/Q vssd1 vssd1 vccd1 vccd1 _2483_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3104_ _3448_/CLK _3104_/D vssd1 vssd1 vccd1 vccd1 _3104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3035_ _3275_/CLK _3035_/D vssd1 vssd1 vccd1 vccd1 _3035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2819_ _3179_/Q _3155_/Q _3131_/Q _3107_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2819_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_55_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3433_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 io_b_dat_o_0[14] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput29 io_b_dat_o_10[0] vssd1 vssd1 vccd1 vccd1 _2422_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1983_ _3282_/Q _1977_/X _1953_/X _1978_/X vssd1 vssd1 vccd1 vccd1 _3282_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2604_ _2604_/A0 _2604_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__mux2_1
X_2535_ _3454_/Q _2534_/B _2537_/B vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__a21o_1
X_2466_ _2459_/X _2461_/X _2462_/Y _2465_/X vssd1 vssd1 vccd1 vccd1 _2466_/X sky130_fd_sc_hd__a31o_4
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2397_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3018_ _3273_/CLK _3018_/D vssd1 vssd1 vccd1 vccd1 _3018_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2320_ _3068_/Q _2316_/X _1722_/A _2317_/X vssd1 vssd1 vccd1 vccd1 _3068_/D sky130_fd_sc_hd__a22o_1
X_2251_ _3117_/Q _2246_/X _2250_/X _2248_/X vssd1 vssd1 vccd1 vccd1 _3117_/D sky130_fd_sc_hd__a22o_1
Xrepeater405 _2632_/S vssd1 vssd1 vccd1 vccd1 _2644_/S sky130_fd_sc_hd__buf_8
X_2182_ _2182_/A vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3333_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1966_ _3294_/Q _1958_/X _1965_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _3294_/D sky130_fd_sc_hd__a22o_1
X_1897_ _1995_/A _2551_/A vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__or2_4
X_2518_ _3396_/Q vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__inv_2
X_3498_ _3500_/CLK _3498_/D vssd1 vssd1 vccd1 vccd1 _3498_/Q sky130_fd_sc_hd__dfxtp_1
Xinput208 io_dat_i[26] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_1
X_2449_ _3383_/Q vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__inv_2
Xinput219 io_dat_i[7] vssd1 vssd1 vccd1 vccd1 _2565_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1820_ _2021_/A vssd1 vssd1 vccd1 vccd1 _1820_/X sky130_fd_sc_hd__clkbuf_2
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1751_ _1846_/A _1798_/B _2300_/C _1828_/B vssd1 vssd1 vccd1 vccd1 _2397_/A sky130_fd_sc_hd__or4_4
X_1682_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2216_/A sky130_fd_sc_hd__inv_2
X_3421_ _3423_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
X_3352_ _3371_/CLK _3352_/D vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfxtp_1
X_2303_ _2317_/A vssd1 vssd1 vccd1 vccd1 _2303_/X sky130_fd_sc_hd__buf_2
X_3283_ _3474_/CLK _3283_/D vssd1 vssd1 vccd1 vccd1 _3283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2234_ _2246_/A vssd1 vssd1 vccd1 vccd1 _2234_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2165_ _2172_/A vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ _3208_/Q _1791_/X _2038_/X _1793_/X vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2998_ input13/X input45/X input61/X input77/X _2610_/S _2611_/S vssd1 vssd1 vccd1
+ vccd1 _2998_/X sky130_fd_sc_hd__mux4_1
X_1949_ _2561_/A vssd1 vssd1 vccd1 vccd1 _1949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _2921_/A0 _2921_/A1 _2921_/A2 _2921_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2921_/X sky130_fd_sc_hd__mux4_1
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2852_ _2848_/X _2849_/X _2850_/X _2851_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2852_/X sky130_fd_sc_hd__mux4_2
X_1803_ _3383_/Q _1799_/X _1774_/X _1801_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__a22o_1
X_2783_ _3170_/Q _3338_/Q _3322_/Q _3306_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2783_/X sky130_fd_sc_hd__mux4_1
X_1734_ _1798_/D vssd1 vssd1 vccd1 vccd1 _1828_/B sky130_fd_sc_hd__buf_1
X_3404_ _3429_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
X_1665_ _3436_/Q _1658_/X _1664_/X _1660_/X vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__a22o_1
X_1596_ _1597_/A _2872_/X vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__and2_1
X_3335_ _3335_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
X_3266_ _3515_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2217_ _3135_/Q _2215_/X _2137_/X _2216_/X vssd1 vssd1 vccd1 vccd1 _3135_/D sky130_fd_sc_hd__a22o_1
X_3197_ _3297_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2148_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2148_/X sky130_fd_sc_hd__buf_2
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _3221_/Q _2073_/X _1967_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput309 _2543_/Y vssd1 vssd1 vccd1 vccd1 io_b_cs_i_9 sky130_fd_sc_hd__clkbuf_2
X_3120_ _3335_/CLK _3120_/D vssd1 vssd1 vccd1 vccd1 _3120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3353_/CLK _3051_/D vssd1 vssd1 vccd1 vccd1 _3051_/Q sky130_fd_sc_hd__dfxtp_1
X_2002_ _3269_/Q _1996_/X _1967_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2904_ _3084_/Q _3368_/Q _3036_/Q _3028_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2904_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2835_ _2515_/Y _2516_/Y _2517_/Y _2518_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2835_/X sky130_fd_sc_hd__mux4_1
X_2766_ _3102_/Q _3078_/Q _3054_/Q _3358_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2766_/X sky130_fd_sc_hd__mux4_1
X_2697_ _2693_/X _2694_/X _2695_/X _2696_/X _2842_/X _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2697_/X sky130_fd_sc_hd__mux4_2
X_1717_ _3418_/Q _1712_/X _1668_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__a22o_1
X_1648_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__clkbuf_2
X_1579_ _1581_/A _2633_/X vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__nor2b_4
XFILLER_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3318_ _3334_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
X_3249_ _3372_/CLK _3249_/D vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2620_ _1497_/A _2832_/X _2620_/S vssd1 vssd1 vccd1 vccd1 _2620_/X sky130_fd_sc_hd__mux2_1
X_2551_ _2551_/A _2552_/B vssd1 vssd1 vccd1 vccd1 _2551_/Y sky130_fd_sc_hd__nor2_1
X_1502_ _1502_/A vssd1 vssd1 vccd1 vccd1 _1502_/Y sky130_fd_sc_hd__inv_2
X_2482_ _3415_/Q vssd1 vssd1 vccd1 vccd1 _2482_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _3447_/CLK _3103_/D vssd1 vssd1 vccd1 vccd1 _3103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3034_ _3273_/CLK _3034_/D vssd1 vssd1 vccd1 vccd1 _3034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ _3059_/Q _3251_/Q _3227_/Q _3203_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2818_/X sky130_fd_sc_hd__mux4_2
X_2749_ _3149_/Q _3125_/Q _3197_/Q _3445_/Q _2750_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2749_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3109_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 io_b_dat_o_0[15] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _3283_/Q _1977_/X _1951_/X _1978_/X vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__a22o_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2603_ _2602_/X _2426_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__mux2_1
X_2534_ _3454_/Q _2534_/B vssd1 vssd1 vccd1 vccd1 _2537_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2465_ _2465_/A _2465_/B _3497_/Q vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__and3_1
X_2396_ _3016_/Q _1752_/X _2038_/A _1754_/X vssd1 vssd1 vccd1 vccd1 _3016_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3017_ _3410_/CLK _3017_/D vssd1 vssd1 vccd1 vccd1 _3017_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2250_/X sky130_fd_sc_hd__buf_2
Xrepeater406 _2594_/S vssd1 vssd1 vccd1 vccd1 _2632_/S sky130_fd_sc_hd__buf_8
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2181_ _2181_/A vssd1 vssd1 vccd1 vccd1 _2181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1965_ _2571_/A vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__clkbuf_2
X_1896_ _3329_/Q _1889_/A _1826_/X _1890_/A vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__a22o_1
X_3497_ _3497_/CLK _3497_/D vssd1 vssd1 vccd1 vccd1 _3497_/Q sky130_fd_sc_hd__dfxtp_2
X_2517_ _3400_/Q vssd1 vssd1 vccd1 vccd1 _2517_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2448_ _3380_/Q vssd1 vssd1 vccd1 vccd1 _2448_/Y sky130_fd_sc_hd__inv_2
Xinput209 io_dat_i[27] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__buf_1
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2379_ _3031_/Q _2377_/X _2327_/X _2378_/X vssd1 vssd1 vccd1 vccd1 _3031_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _3405_/Q _1744_/X _1730_/X _1746_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__a22o_1
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1681_ _2215_/A vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__clkbuf_2
X_3420_ _3420_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
X_3351_ _3351_/CLK _3351_/D vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2302_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2317_/A sky130_fd_sc_hd__inv_2
X_3282_ _3474_/CLK _3282_/D vssd1 vssd1 vccd1 vccd1 _3282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2233_ _3124_/Q _2225_/X _2232_/X _2227_/X vssd1 vssd1 vccd1 vccd1 _3124_/D sky130_fd_sc_hd__a22o_1
X_2164_ _3172_/Q _2153_/X _2134_/X _2156_/X vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2095_ _3209_/Q _2088_/A _1955_/X _2089_/A vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2997_ _2993_/X _2994_/X _2995_/X _2996_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2997_/X sky130_fd_sc_hd__mux4_1
X_1948_ _3301_/Q _1943_/X _1947_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__a22o_1
X_1879_ _3342_/Q _1874_/X _1636_/X _1876_/X vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2920_ input25/X input57/X input73/X input89/X _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2920_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _3405_/Q _3401_/Q _3409_/Q _3381_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2851_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1802_ _3384_/Q _1799_/X _1770_/X _1801_/X vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__a22o_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2782_ _2778_/X _2779_/X _2780_/X _2781_/X _2901_/S0 _2997_/S1 vssd1 vssd1 vccd1
+ vccd1 _2782_/X sky130_fd_sc_hd__mux4_2
X_1733_ _1847_/A vssd1 vssd1 vccd1 vccd1 _1798_/B sky130_fd_sc_hd__buf_1
X_3403_ _3482_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
X_1664_ _1722_/A vssd1 vssd1 vccd1 vccd1 _1664_/X sky130_fd_sc_hd__buf_2
X_1595_ _1597_/A _2864_/X vssd1 vssd1 vccd1 vccd1 _3469_/D sky130_fd_sc_hd__and2_1
X_3334_ _3334_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
X_3265_ _3303_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
X_2216_ _2216_/A vssd1 vssd1 vccd1 vccd1 _2216_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3196_ _3444_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _3179_/Q _2136_/X _2146_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2078_ _3222_/Q _2073_/X _1965_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3448_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3050_ _3353_/CLK _3050_/D vssd1 vssd1 vccd1 vccd1 _3050_/Q sky130_fd_sc_hd__dfxtp_1
X_2001_ _3270_/Q _1996_/X _1965_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2903_ _3180_/Q _3156_/Q _3132_/Q _3108_/Q _2918_/S0 _2944_/S1 vssd1 vssd1 vccd1
+ vccd1 _2903_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2834_ _2448_/Y _2521_/Y _2513_/Y _2514_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2834_/X sky130_fd_sc_hd__mux4_2
X_2765_ _3198_/Q _3446_/Q _3150_/Q _3126_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2765_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2696_ _3314_/Q _3298_/Q _3162_/Q _3330_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2696_/X sky130_fd_sc_hd__mux4_1
X_1716_ _3419_/Q _1712_/X _1666_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__a22o_1
X_1647_ _3443_/Q _1643_/X _1645_/X _1646_/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__a22o_1
X_1578_ _1581_/A _2632_/X vssd1 vssd1 vccd1 vccd1 _3483_/D sky130_fd_sc_hd__nor2b_4
X_3317_ _3333_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3248_ _3294_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
X_3179_ _3497_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2550_ _2550_/A _2552_/B vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__nor2_1
X_1501_ _3518_/Q _1483_/B _1484_/A _1508_/B vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__o211a_1
X_2481_ _2490_/A _2777_/X vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__and2_1
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3102_ _3447_/CLK _3102_/D vssd1 vssd1 vccd1 vccd1 _3102_/Q sky130_fd_sc_hd__dfxtp_1
X_3033_ _3273_/CLK _3033_/D vssd1 vssd1 vccd1 vccd1 _3033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2817_ _2813_/X _2814_/X _2815_/X _2816_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2817_/X sky130_fd_sc_hd__mux4_2
X_2748_ _3053_/Q _3357_/Q _3101_/Q _3077_/Q _2750_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2748_/X sky130_fd_sc_hd__mux4_2
X_2679_ _2984_/X _2678_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2679_/X sky130_fd_sc_hd__mux2_2
XFILLER_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1981_ _3284_/Q _1977_/X _1949_/X _1978_/X vssd1 vssd1 vccd1 vccd1 _3284_/D sky130_fd_sc_hd__a22o_1
X_2602_ _2602_/A0 _2602_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2533_ _3453_/Q _2532_/B _2534_/B vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__a21bo_1
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _2458_/Y _2464_/A2 _1557_/X _2464_/B2 _2460_/Y vssd1 vssd1 vccd1 vccd1 _2465_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2395_ _3017_/Q _2387_/A _2340_/X _2388_/A vssd1 vssd1 vccd1 vccd1 _3017_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ _3410_/CLK _3016_/D vssd1 vssd1 vccd1 vccd1 _3016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XINSDIODE4_0 _2571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater407 _2606_/S vssd1 vssd1 vccd1 vccd1 _2594_/S sky130_fd_sc_hd__buf_8
X_2180_ _3160_/Q _1721_/X _2134_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__a22o_1
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _3295_/Q _1958_/X _1963_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _3330_/Q _1889_/X _1824_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__a22o_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3497_/CLK _3496_/D vssd1 vssd1 vccd1 vccd1 _3496_/Q sky130_fd_sc_hd__dfxtp_2
X_2516_ _3364_/Q vssd1 vssd1 vccd1 vccd1 _2516_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2447_ _2480_/A _2597_/X vssd1 vssd1 vccd1 vccd1 _2447_/X sky130_fd_sc_hd__and2_1
X_2378_ _2378_/A vssd1 vssd1 vccd1 vccd1 _2378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1680_ _2546_/A _1816_/A vssd1 vssd1 vccd1 vccd1 _2215_/A sky130_fd_sc_hd__or2_4
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3350_ _3350_/CLK _3350_/D vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfxtp_1
X_2301_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2301_/X sky130_fd_sc_hd__buf_2
X_3281_ _3297_/CLK _3281_/D vssd1 vssd1 vccd1 vccd1 _3281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2232_ _2569_/A vssd1 vssd1 vccd1 vccd1 _2232_/X sky130_fd_sc_hd__buf_2
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2163_ _3173_/Q _2153_/X _2162_/X _2156_/X vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__a22o_1
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2094_ _3210_/Q _2088_/X _1953_/X _2089_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _3405_/Q _3401_/Q _3409_/Q _3381_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2996_/X sky130_fd_sc_hd__mux4_1
X_1947_ _1947_/A vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__buf_2
X_1878_ _3343_/Q _1874_/X _1634_/X _1876_/X vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3479_ _3501_/CLK _3479_/D vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2850_ _3421_/Q _3361_/Q _3397_/Q _3393_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2850_/X sky130_fd_sc_hd__mux4_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1801_ _1987_/A vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__clkbuf_2
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _3099_/Q _3075_/Q _3051_/Q _3355_/Q _2913_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2781_/X sky130_fd_sc_hd__mux4_1
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1732_ _1846_/A vssd1 vssd1 vccd1 vccd1 _2342_/A sky130_fd_sc_hd__buf_1
X_1663_ _3437_/Q _1658_/X _1662_/X _1660_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__a22o_1
X_3402_ _3410_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
X_1594_ _1597_/A _2861_/X vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__and2_1
X_3333_ _3333_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
X_3264_ _3307_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2215_ _2215_/A vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3195_ _3355_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2146_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2146_/X sky130_fd_sc_hd__buf_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2077_ _3223_/Q _2073_/X _1963_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _3223_/D sky130_fd_sc_hd__a22o_1
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2979_ _2975_/X _2976_/X _2977_/X _2978_/X input7/X input8/X vssd1 vssd1 vccd1 vccd1
+ _2979_/X sky130_fd_sc_hd__mux4_2
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3501_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _3271_/Q _1996_/X _1963_/X _1998_/X vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__a22o_1
XFILLER_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _3060_/Q _3252_/Q _3228_/Q _3204_/Q _2682_/S _2905_/S1 vssd1 vssd1 vccd1 vccd1
+ _2902_/X sky130_fd_sc_hd__mux4_2
X_2833_ _2524_/Y _2510_/Y _2435_/Y _2434_/Y _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2833_/X sky130_fd_sc_hd__mux4_2
X_2764_ _3294_/Q _3270_/Q _3246_/Q _3222_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2764_/X sky130_fd_sc_hd__mux4_2
X_1715_ _3420_/Q _1712_/X _1664_/X _1714_/X vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__a22o_1
X_2695_ _3234_/Q _3210_/Q _3282_/Q _3258_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2695_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1646_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__clkbuf_2
X_1577_ _1581_/A _2631_/X vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__nor2b_4
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3316_ _3333_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3247_ _3294_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3247_/Q sky130_fd_sc_hd__dfxtp_1
X_3178_ _3501_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2129_ _3187_/Q _2122_/X _2128_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2480_ _2480_/A _2591_/X vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__and2_1
X_1500_ _1502_/A vssd1 vssd1 vccd1 vccd1 _2687_/S sky130_fd_sc_hd__buf_2
XFILLER_68_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3101_ _3445_/CLK _3101_/D vssd1 vssd1 vccd1 vccd1 _3101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput190 io_dat_i[0] vssd1 vssd1 vccd1 vccd1 _2558_/A sky130_fd_sc_hd__buf_4
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3032_ _3398_/CLK _3032_/D vssd1 vssd1 vccd1 vccd1 _3032_/Q sky130_fd_sc_hd__dfxtp_1
X_2816_ _3020_/Q _3012_/Q _3004_/Q _3276_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2816_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2747_ _2743_/X _2744_/X _2745_/X _2746_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2747_/X sky130_fd_sc_hd__mux4_2
X_2678_ _2678_/A0 _2678_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2678_/X sky130_fd_sc_hd__mux2_2
X_1629_ _1658_/A vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__buf_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3087_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _3285_/Q _1977_/X _1947_/X _1978_/X vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__a22o_1
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2601_ _2600_/X _2429_/X _2609_/S vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__mux2_1
X_2532_ _3453_/Q _2532_/B vssd1 vssd1 vccd1 vccd1 _2534_/B sky130_fd_sc_hd__or2_2
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2463_ _2458_/Y _2463_/A2 _1557_/X _2463_/B2 _3496_/Q vssd1 vssd1 vccd1 vccd1 _2465_/A
+ sky130_fd_sc_hd__a221o_1
X_2394_ _3018_/Q _2387_/A _2338_/X _2388_/A vssd1 vssd1 vccd1 vccd1 _3018_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3015_ _3277_/CLK _3015_/D vssd1 vssd1 vccd1 vccd1 _3015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater408 _2610_/S vssd1 vssd1 vccd1 vccd1 _2606_/S sky130_fd_sc_hd__buf_8
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1963_ _2572_/A vssd1 vssd1 vccd1 vccd1 _1963_/X sky130_fd_sc_hd__clkbuf_2
X_1894_ _3331_/Q _1889_/X _1822_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__a22o_1
X_3495_ _3519_/CLK _3495_/D vssd1 vssd1 vccd1 vccd1 _3495_/Q sky130_fd_sc_hd__dfxtp_2
X_2515_ _3424_/Q vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__inv_2
X_2446_ _2479_/A _2446_/B vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__and2_1
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2377_ _2377_/A vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _3410_/CLK _3280_/D vssd1 vssd1 vccd1 vccd1 _3280_/Q sky130_fd_sc_hd__dfxtp_1
X_2300_ _2342_/A _2342_/B _2300_/C _2300_/D vssd1 vssd1 vccd1 vccd1 _2316_/A sky130_fd_sc_hd__or4_4
X_2231_ _3125_/Q _2225_/X _2162_/X _2227_/X vssd1 vssd1 vccd1 vccd1 _3125_/D sky130_fd_sc_hd__a22o_1
XFILLER_78_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2162_ _2570_/A vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2093_ _3211_/Q _2088_/X _1951_/X _2089_/X vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2995_ _3421_/Q _3361_/Q _3397_/Q _3393_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2995_/X sky130_fd_sc_hd__mux4_1
X_1946_ _3302_/Q _1943_/X _1944_/X _1945_/X vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__a22o_1
X_1877_ _3344_/Q _1874_/X _1630_/X _1876_/X vssd1 vssd1 vccd1 vccd1 _3344_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3478_ _3497_/CLK _3478_/D vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2429_ _2429_/A _2429_/B vssd1 vssd1 vccd1 vccd1 _2429_/X sky130_fd_sc_hd__and2_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ _1986_/A vssd1 vssd1 vccd1 vccd1 _1987_/A sky130_fd_sc_hd__inv_2
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _3195_/Q _3443_/Q _3147_/Q _3123_/Q _2913_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2780_/X sky130_fd_sc_hd__mux4_1
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1731_ _3413_/Q _1721_/X _1730_/X _1724_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1662_ _1947_/A vssd1 vssd1 vccd1 vccd1 _1662_/X sky130_fd_sc_hd__buf_2
X_3401_ _3409_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
X_1593_ _1597_/A _2858_/X vssd1 vssd1 vccd1 vccd1 _3471_/D sky130_fd_sc_hd__and2_1
X_3332_ _3333_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
X_3263_ _3303_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2214_ _3136_/Q _1681_/X _2134_/X _1683_/X vssd1 vssd1 vccd1 vccd1 _3136_/D sky130_fd_sc_hd__a22o_1
X_3194_ _3515_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2145_ _3180_/Q _2136_/X _2144_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _3180_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2076_ _3224_/Q _2073_/X _1959_/X _2075_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__a22o_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2978_ _3090_/Q _3066_/Q _3042_/Q _3346_/Q _1676_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2978_/X sky130_fd_sc_hd__mux4_1
X_1929_ _2038_/A vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_58_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3294_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2901_ _2897_/X _2898_/X _2899_/X _2900_/X _2901_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2901_/X sky130_fd_sc_hd__mux4_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2832_ _2828_/X _2829_/X _2830_/X _2831_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2832_/X sky130_fd_sc_hd__mux4_2
X_2763_ _3174_/Q _3342_/Q _3326_/Q _3310_/Q _2785_/S0 _2911_/S1 vssd1 vssd1 vccd1
+ vccd1 _2763_/X sky130_fd_sc_hd__mux4_2
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1714_ _2328_/A vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__buf_2
X_2694_ _3138_/Q _3114_/Q _3186_/Q _3434_/Q _2852_/X _2716_/S1 vssd1 vssd1 vccd1 vccd1
+ _2694_/X sky130_fd_sc_hd__mux4_2
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1645_ _2041_/A vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__clkbuf_2
X_1576_ _1582_/A vssd1 vssd1 vccd1 vccd1 _1581_/A sky130_fd_sc_hd__buf_4
X_3315_ _3331_/CLK _3315_/D vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3246_ _3294_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3177_ _3501_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2128_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2128_/X sky130_fd_sc_hd__clkbuf_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _3235_/Q _2052_/X _1951_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__a22o_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ _3439_/CLK _3100_/D vssd1 vssd1 vccd1 vccd1 _3100_/Q sky130_fd_sc_hd__dfxtp_1
Xinput180 io_b_dat_o_9[1] vssd1 vssd1 vccd1 vccd1 _2608_/A1 sky130_fd_sc_hd__clkbuf_1
X_3031_ _3087_/CLK _3031_/D vssd1 vssd1 vccd1 vccd1 _3031_/Q sky130_fd_sc_hd__dfxtp_1
Xinput191 io_dat_i[10] vssd1 vssd1 vccd1 vccd1 _2568_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3437_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2815_ _3084_/Q _3368_/Q _3036_/Q _3028_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2815_/X sky130_fd_sc_hd__mux4_1
X_2746_ _3324_/Q _3308_/Q _3172_/Q _3340_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2746_/X sky130_fd_sc_hd__mux4_2
X_2677_ _3498_/Q _2979_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2677_/X sky130_fd_sc_hd__mux2_1
X_1628_ _2543_/A _2300_/D vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__or2_4
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1559_ _1557_/X _1539_/A _1944_/A _1541_/A _1592_/A vssd1 vssd1 vccd1 vccd1 _3495_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3229_ _3353_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _2600_/A0 _2600_/A1 _2606_/S vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__mux2_1
X_2531_ _3452_/Q _2527_/B _2532_/B vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__a21bo_1
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2462_ _3497_/Q vssd1 vssd1 vccd1 vccd1 _2462_/Y sky130_fd_sc_hd__inv_2
X_2393_ _3019_/Q _2387_/X _2336_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _3019_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _3277_/CLK _3014_/D vssd1 vssd1 vccd1 vccd1 _3014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2729_ _3145_/Q _3121_/Q _3193_/Q _3441_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2729_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater409 _2996_/S0 vssd1 vssd1 vccd1 vccd1 _2610_/S sky130_fd_sc_hd__buf_8
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1962_ _3296_/Q _1958_/X _1959_/X _1961_/X vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1893_ _3332_/Q _1889_/X _1818_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__a22o_1
X_3494_ _3518_/CLK _3494_/D vssd1 vssd1 vccd1 vccd1 _3494_/Q sky130_fd_sc_hd__dfxtp_1
X_2514_ _3428_/Q vssd1 vssd1 vccd1 vccd1 _2514_/Y sky130_fd_sc_hd__inv_2
X_2445_ _3430_/Q vssd1 vssd1 vccd1 vccd1 _2445_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _3032_/Q _1769_/X _2324_/X _1772_/X vssd1 vssd1 vccd1 vccd1 _3032_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2230_ _3126_/Q _2225_/X _2160_/X _2227_/X vssd1 vssd1 vccd1 vccd1 _3126_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2161_ _3174_/Q _2153_/X _2160_/X _2156_/X vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2092_ _3212_/Q _2088_/X _1949_/X _2089_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _3377_/Q _3413_/Q _3429_/Q _3425_/Q _2610_/S _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2994_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1945_ _1945_/A vssd1 vssd1 vccd1 vccd1 _1945_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1876_ _1890_/A vssd1 vssd1 vccd1 vccd1 _1876_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3477_ _3501_/CLK _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2428_ _3386_/Q vssd1 vssd1 vccd1 vccd1 _2428_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2359_ _2359_/A vssd1 vssd1 vccd1 vccd1 _2359_/X sky130_fd_sc_hd__buf_2
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1730_ _1730_/A vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__buf_2
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1661_ _3438_/Q _1658_/X _1659_/X _1660_/X vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ _3424_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
X_1592_ _1592_/A vssd1 vssd1 vccd1 vccd1 _1597_/A sky130_fd_sc_hd__buf_1
X_3331_ _3331_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
X_3262_ _3296_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2213_ _3137_/Q _2206_/A _2132_/X _2207_/A vssd1 vssd1 vccd1 vccd1 _3137_/D sky130_fd_sc_hd__a22o_1
X_3193_ _3443_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2144_ _2565_/A vssd1 vssd1 vccd1 vccd1 _2144_/X sky130_fd_sc_hd__buf_2
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2075_ _2089_/A vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2977_ _3186_/Q _3434_/Q _3138_/Q _3114_/Q _1676_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2977_/X sky130_fd_sc_hd__mux4_1
X_1928_ _3309_/Q _1922_/X _1638_/X _1924_/X vssd1 vssd1 vccd1 vccd1 _3309_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1859_ _3355_/Q _1857_/X _1645_/X _1858_/X vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3519_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2900_ _3096_/Q _3072_/Q _3048_/Q _3352_/Q _2913_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2900_/X sky130_fd_sc_hd__mux4_2
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _3017_/Q _3009_/Q _3001_/Q _3273_/Q _2851_/S0 _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2831_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2762_ _2758_/X _2759_/X _2760_/X _2761_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2762_/X sky130_fd_sc_hd__mux4_2
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1713_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2328_/A sky130_fd_sc_hd__inv_2
X_2693_ _3042_/Q _3346_/Q _3090_/Q _3066_/Q _2852_/X _2716_/S1 vssd1 vssd1 vccd1 vccd1
+ _2693_/X sky130_fd_sc_hd__mux4_2
X_1644_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2041_/A sky130_fd_sc_hd__clkbuf_2
X_1575_ _1575_/A _2630_/X vssd1 vssd1 vccd1 vccd1 _3485_/D sky130_fd_sc_hd__nor2b_2
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3314_ _3331_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3245_ _3297_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3176_ _3506_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2127_ _3188_/Q _2122_/X _2126_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__a22o_1
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _3236_/Q _2052_/X _1949_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _3236_/D sky130_fd_sc_hd__a22o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput181 io_b_dat_o_9[2] vssd1 vssd1 vccd1 vccd1 _2606_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput170 io_b_dat_o_8[7] vssd1 vssd1 vccd1 vccd1 _2596_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3030_ _3087_/CLK _3030_/D vssd1 vssd1 vccd1 vccd1 _3030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput192 io_dat_i[11] vssd1 vssd1 vccd1 vccd1 _2569_/A sky130_fd_sc_hd__buf_2
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2814_ _3180_/Q _3156_/Q _3132_/Q _3108_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2814_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2745_ _3244_/Q _3220_/Q _3292_/Q _3268_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2745_/X sky130_fd_sc_hd__mux4_2
X_2676_ _2972_/X _2973_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__mux2_1
X_1627_ _2342_/D vssd1 vssd1 vccd1 vccd1 _2300_/D sky130_fd_sc_hd__clkbuf_2
X_1558_ _2563_/A vssd1 vssd1 vccd1 vccd1 _1944_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1489_ _1485_/Y _3501_/Q _1485_/Y _3501_/Q vssd1 vssd1 vccd1 vccd1 _1490_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3228_ _3279_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3456_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3514_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2530_ _3451_/Q _2526_/B _2527_/B vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__a21bo_1
X_2461_ _2458_/Y _2461_/A2 _1557_/X _2461_/B2 _2460_/Y vssd1 vssd1 vccd1 vccd1 _2461_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2392_ _3020_/Q _2387_/X _2334_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _3020_/D sky130_fd_sc_hd__a22o_1
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3013_ _3277_/CLK _3013_/D vssd1 vssd1 vccd1 vccd1 _3013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2728_ _3049_/Q _3353_/Q _3097_/Q _3073_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2728_/X sky130_fd_sc_hd__mux4_2
X_2659_ _2919_/X _2658_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1961_ _1978_/A vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1892_ _3333_/Q _1889_/X _1662_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__a22o_1
X_2513_ _3432_/Q vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__inv_2
X_3493_ _3493_/CLK _3493_/D vssd1 vssd1 vccd1 vccd1 _3493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2444_ _3426_/Q vssd1 vssd1 vccd1 vccd1 _2444_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2375_ _3033_/Q _2367_/A _2340_/X _2368_/A vssd1 vssd1 vccd1 vccd1 _3033_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_0 _2861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2571_/A vssd1 vssd1 vccd1 vccd1 _2160_/X sky130_fd_sc_hd__clkbuf_2
X_2091_ _3213_/Q _2088_/X _2056_/X _2089_/X vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__a22o_1
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _3417_/Q _3373_/Q _3389_/Q _3385_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2993_/X sky130_fd_sc_hd__mux4_2
XFILLER_61_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1944_ _1944_/A vssd1 vssd1 vccd1 vccd1 _1944_/X sky130_fd_sc_hd__buf_2
X_1875_ _1889_/A vssd1 vssd1 vccd1 vccd1 _1890_/A sky130_fd_sc_hd__inv_2
X_3476_ _3501_/CLK _3476_/D vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2427_ _2430_/A _2603_/X vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__and2_1
XFILLER_84_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2358_ _2358_/A vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _3089_/Q _2282_/A _2132_/X _2283_/A vssd1 vssd1 vccd1 vccd1 _3089_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1660_ _1660_/A vssd1 vssd1 vccd1 vccd1 _1660_/X sky130_fd_sc_hd__clkbuf_2
X_1591_ _1591_/A _2855_/X vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__and2_1
X_3330_ _3331_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3261_ _3301_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2212_ _3138_/Q _2206_/X _2130_/X _2207_/X vssd1 vssd1 vccd1 vccd1 _3138_/D sky130_fd_sc_hd__a22o_1
X_3192_ _3504_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_1
X_2143_ _3181_/Q _2136_/X _2142_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__a22o_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2074_ _2088_/A vssd1 vssd1 vccd1 vccd1 _2089_/A sky130_fd_sc_hd__inv_2
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2976_ _3282_/Q _3258_/Q _3234_/Q _3210_/Q input5/X input6/X vssd1 vssd1 vccd1 vccd1
+ _2976_/X sky130_fd_sc_hd__mux4_2
X_1927_ _3310_/Q _1922_/X _1636_/X _1924_/X vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__a22o_1
X_1858_ _1865_/A vssd1 vssd1 vccd1 vccd1 _1858_/X sky130_fd_sc_hd__clkbuf_2
X_1789_ _1815_/A input8/X _1789_/C vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__or3_4
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3459_ _3485_/CLK _3459_/D vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2830_ _3081_/Q _3365_/Q _3033_/Q _3025_/Q _2851_/S0 _2851_/S1 vssd1 vssd1 vccd1
+ vccd1 _2830_/X sky130_fd_sc_hd__mux4_2
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _3103_/Q _3079_/Q _3055_/Q _3359_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2761_/X sky130_fd_sc_hd__mux4_1
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2692_ _2688_/X _2689_/X _2690_/X _2691_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2692_/X sky130_fd_sc_hd__mux4_2
X_1712_ _2326_/A vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1643_ _1658_/A vssd1 vssd1 vccd1 vccd1 _1643_/X sky130_fd_sc_hd__clkbuf_2
X_1574_ _1575_/A _2629_/X vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__nor2b_1
X_3313_ _3433_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
X_3244_ _3297_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3175_ _3506_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
X_2126_ _2561_/A vssd1 vssd1 vccd1 vccd1 _2126_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _3237_/Q _2052_/X _2056_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__a22o_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2959_ input22/X input54/X input70/X input86/X _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2959_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater390 _2905_/S1 vssd1 vssd1 vccd1 vccd1 _2911_/S1 sky130_fd_sc_hd__buf_8
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput160 io_b_dat_o_8[12] vssd1 vssd1 vccd1 vccd1 _2585_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput171 io_b_dat_o_8[8] vssd1 vssd1 vccd1 vccd1 _2594_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput182 io_b_dat_o_9[3] vssd1 vssd1 vccd1 vccd1 _2604_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput193 io_dat_i[12] vssd1 vssd1 vccd1 vccd1 _2570_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2813_ _3060_/Q _3252_/Q _3228_/Q _3204_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2813_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2744_ _3148_/Q _3124_/Q _3196_/Q _3444_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2744_/X sky130_fd_sc_hd__mux4_1
X_2675_ _2971_/X _2674_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__mux2_1
X_1626_ _1626_/A input2/X input3/X _1626_/D vssd1 vssd1 vccd1 vccd1 _2342_/D sky130_fd_sc_hd__or4_4
X_1557_ _3495_/Q vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__buf_2
X_1488_ _1482_/A _3499_/Q _1482_/A _3499_/Q vssd1 vssd1 vccd1 vccd1 _1490_/C sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3227_ _3371_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
X_3158_ _3456_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2109_ _2123_/A vssd1 vssd1 vccd1 vccd1 _2109_/X sky130_fd_sc_hd__clkbuf_2
X_3089_ _3502_/CLK _3089_/D vssd1 vssd1 vccd1 vccd1 _3089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3409_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2460_ _3496_/Q vssd1 vssd1 vccd1 vccd1 _2460_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2391_ _3021_/Q _2387_/X _2332_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _3021_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3012_ _3277_/CLK _3012_/D vssd1 vssd1 vccd1 vccd1 _3012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2727_ _2723_/X _2724_/X _2725_/X _2726_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2727_/X sky130_fd_sc_hd__mux4_2
X_2658_ _2658_/A0 _2658_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__mux2_2
X_2589_ _2588_/X _2486_/X _2595_/S vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__mux2_1
X_1609_ _1609_/A _3000_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__and2_1
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1978_/A sky130_fd_sc_hd__inv_2
X_1891_ _3334_/Q _1889_/X _1659_/X _1890_/X vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__a22o_1
X_2512_ _2523_/A _2580_/X vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__and2_1
X_3492_ _3518_/CLK _3492_/D vssd1 vssd1 vccd1 vccd1 _3492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2443_ _3422_/Q vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__inv_2
X_2374_ _3034_/Q _2367_/A _2338_/X _2368_/A vssd1 vssd1 vccd1 vccd1 _3034_/D sky130_fd_sc_hd__a22o_1
XFILLER_37_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_1 _2624_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2090_ _3214_/Q _2088_/X _2053_/X _2089_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__a22o_1
XFILLER_81_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2992_ _2988_/X _2989_/X _2990_/X _2991_/X _2992_/S0 _2992_/S1 vssd1 vssd1 vccd1
+ vccd1 _2992_/X sky130_fd_sc_hd__mux4_1
X_1943_ _1943_/A vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1874_ _1889_/A vssd1 vssd1 vccd1 vccd1 _1874_/X sky130_fd_sc_hd__clkbuf_2
X_3475_ _3497_/CLK _3475_/D vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfxtp_4
X_2426_ _2429_/A _2426_/B vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__and2_1
XFILLER_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2357_ _3047_/Q _2351_/X _2336_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3047_/D sky130_fd_sc_hd__a22o_1
X_2288_ _3090_/Q _2282_/X _2130_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _3090_/D sky130_fd_sc_hd__a22o_1
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1590_ _1590_/A _2554_/A vssd1 vssd1 vccd1 vccd1 _3473_/D sky130_fd_sc_hd__nor2_1
X_3260_ _3295_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2211_ _3139_/Q _2206_/X _2128_/X _2207_/X vssd1 vssd1 vccd1 vccd1 _3139_/D sky130_fd_sc_hd__a22o_1
X_3191_ _3502_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2142_ _2566_/A vssd1 vssd1 vccd1 vccd1 _2142_/X sky130_fd_sc_hd__buf_2
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _2088_/A vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _3162_/Q _3330_/Q _3314_/Q _3298_/Q _1700_/A input6/X vssd1 vssd1 vccd1 vccd1
+ _2975_/X sky130_fd_sc_hd__mux4_2
X_1926_ _3311_/Q _1922_/X _1634_/X _1924_/X vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__a22o_1
X_1857_ _1864_/A vssd1 vssd1 vccd1 vccd1 _1857_/X sky130_fd_sc_hd__clkbuf_2
X_1788_ _3389_/Q _1782_/X _1778_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3458_ _3485_/CLK _3458_/D vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfxtp_1
X_2409_ _3007_/Q _2407_/X _2041_/A _2408_/X vssd1 vssd1 vccd1 vccd1 _3007_/D sky130_fd_sc_hd__a22o_1
X_3389_ _3392_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_36_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2760_ _3199_/Q _3447_/Q _3151_/Q _3127_/Q _2910_/S0 _2913_/S1 vssd1 vssd1 vccd1
+ vccd1 _2760_/X sky130_fd_sc_hd__mux4_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2691_ _3313_/Q _3297_/Q _3161_/Q _3329_/Q _2716_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2691_/X sky130_fd_sc_hd__mux4_1
X_1711_ _1760_/A _2553_/A vssd1 vssd1 vccd1 vccd1 _2326_/A sky130_fd_sc_hd__or2_4
XFILLER_6_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1642_ _3444_/Q _1629_/X _1641_/X _1632_/X vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__a22o_1
X_1573_ _1575_/A _2628_/X vssd1 vssd1 vccd1 vccd1 _3487_/D sky130_fd_sc_hd__nor2b_1
X_3312_ _3344_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
X_3243_ _3303_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
X_3174_ _3506_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2125_ _3189_/Q _2122_/X _2056_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2562_/A vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__buf_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2958_ _2954_/X _2955_/X _2956_/X _2957_/X _2684_/S _2997_/S1 vssd1 vssd1 vccd1 vccd1
+ _2958_/X sky130_fd_sc_hd__mux4_1
X_1909_ _3322_/Q _1906_/X _1649_/X _1907_/X vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__a22o_1
X_2889_ _3061_/Q _3253_/Q _3229_/Q _3205_/Q _2918_/S0 _2905_/S1 vssd1 vssd1 vccd1
+ vccd1 _2889_/X sky130_fd_sc_hd__mux4_1
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater380 _3476_/Q vssd1 vssd1 vccd1 vccd1 _2851_/S1 sky130_fd_sc_hd__buf_12
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater391 _2944_/S1 vssd1 vssd1 vccd1 vccd1 _2905_/S1 sky130_fd_sc_hd__buf_8
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput150 io_b_dat_o_7[3] vssd1 vssd1 vccd1 vccd1 _2960_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput161 io_b_dat_o_8[13] vssd1 vssd1 vccd1 vccd1 _2582_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput172 io_b_dat_o_8[9] vssd1 vssd1 vccd1 vccd1 _2592_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput183 io_b_dat_o_9[4] vssd1 vssd1 vccd1 vccd1 _2602_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput194 io_dat_i[13] vssd1 vssd1 vccd1 vccd1 _2571_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2812_ _2808_/X _2809_/X _2810_/X _2811_/X _3477_/Q _3478_/Q vssd1 vssd1 vccd1 vccd1
+ _2812_/X sky130_fd_sc_hd__mux4_2
X_2743_ _3052_/Q _3356_/Q _3100_/Q _3076_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2743_/X sky130_fd_sc_hd__mux4_2
X_2674_ _2674_/A0 _2674_/A1 _2682_/S vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__mux2_4
X_1625_ _2224_/A _1847_/A _2300_/C vssd1 vssd1 vccd1 vccd1 _2543_/A sky130_fd_sc_hd__or3_4
X_1556_ _3496_/Q _1539_/A _1941_/A _1541_/A _1592_/A vssd1 vssd1 vccd1 vccd1 _3496_/D
+ sky130_fd_sc_hd__o221a_1
X_1487_ _1482_/B _3498_/Q _1482_/B _3498_/Q vssd1 vssd1 vccd1 vccd1 _1490_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _3372_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3157_ _3180_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2108_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__inv_2
XFILLER_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3088_ _3398_/CLK _3088_/D vssd1 vssd1 vccd1 vccd1 _3088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2039_ _3244_/Q _2031_/X _2038_/X _2033_/X vssd1 vssd1 vccd1 vccd1 _3244_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3336_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2390_ _3022_/Q _2387_/X _2330_/X _2388_/X vssd1 vssd1 vccd1 vccd1 _3022_/D sky130_fd_sc_hd__a22o_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3011_ _3019_/CLK _3011_/D vssd1 vssd1 vccd1 vccd1 _3011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2726_ _3320_/Q _3304_/Q _3168_/Q _3336_/Q _2750_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2726_/X sky130_fd_sc_hd__mux4_1
X_2657_ _3496_/Q _2914_/X _2669_/S vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__mux2_1
X_1608_ _1609_/A _2987_/X vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__and2_1
X_2588_ _2588_/A0 _2588_/A1 _2594_/S vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1539_ _1539_/A vssd1 vssd1 vccd1 vccd1 _1539_/X sky130_fd_sc_hd__buf_2
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3209_ _3297_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1890_ _1890_/A vssd1 vssd1 vccd1 vccd1 _1890_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2511_ _2522_/A _2511_/B vssd1 vssd1 vccd1 vccd1 _2511_/X sky130_fd_sc_hd__and2_1
X_3491_ _3518_/CLK _3491_/D vssd1 vssd1 vccd1 vccd1 _3491_/Q sky130_fd_sc_hd__dfxtp_1
X_2442_ _3378_/Q vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2373_ _3035_/Q _2367_/X _2336_/X _2368_/X vssd1 vssd1 vccd1 vccd1 _3035_/D sky130_fd_sc_hd__a22o_1
XFILLER_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _3141_/Q _3117_/Q _3189_/Q _3437_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2709_/X sky130_fd_sc_hd__mux4_2
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_2 _2674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2991_ _3089_/Q _3065_/Q _3041_/Q _3345_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2991_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1942_ _3303_/Q _1931_/X _1941_/X _1933_/X vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__a22o_1
X_1873_ _1995_/A _2552_/A vssd1 vssd1 vccd1 vccd1 _1889_/A sky130_fd_sc_hd__or2_4
X_3474_ _3474_/CLK _3474_/D vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2425_ _2430_/A _2605_/X vssd1 vssd1 vccd1 vccd1 _2425_/X sky130_fd_sc_hd__and2_1
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2356_ _3048_/Q _2351_/X _2334_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3048_/D sky130_fd_sc_hd__a22o_1
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2287_ _3091_/Q _2282_/X _2128_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _3091_/D sky130_fd_sc_hd__a22o_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _3140_/Q _2206_/X _2126_/X _2207_/X vssd1 vssd1 vccd1 vccd1 _3140_/D sky130_fd_sc_hd__a22o_1
X_3190_ _3438_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2141_ _3182_/Q _2136_/X _2140_/X _2138_/X vssd1 vssd1 vccd1 vccd1 _3182_/D sky130_fd_sc_hd__a22o_1
XFILLER_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2072_ _2190_/A _2545_/A vssd1 vssd1 vccd1 vccd1 _2088_/A sky130_fd_sc_hd__or2_4
XFILLER_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2974_ _2673_/X _2675_/X _2676_/X _2417_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2974_/X sky130_fd_sc_hd__mux4_1
X_1925_ _3312_/Q _1922_/X _1630_/X _1924_/X vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3372_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1856_ _3356_/Q _1849_/X _1641_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__a22o_1
XFILLER_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1787_ _3390_/Q _1782_/X _1776_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__a22o_1
X_3457_ _3485_/CLK _3457_/D vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _2408_/A vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__clkbuf_2
X_3388_ _3420_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2339_ _3058_/Q _2326_/A _2338_/X _2328_/A vssd1 vssd1 vccd1 vccd1 _3058_/D sky130_fd_sc_hd__a22o_1
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ _3233_/Q _3209_/Q _3281_/Q _3257_/Q _2750_/S0 _2847_/X vssd1 vssd1 vccd1 vccd1
+ _2690_/X sky130_fd_sc_hd__mux4_1
X_1710_ _2224_/A _1780_/B _2266_/C vssd1 vssd1 vccd1 vccd1 _2553_/A sky130_fd_sc_hd__or3_4
XFILLER_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1641_ _2038_/A vssd1 vssd1 vccd1 vccd1 _1641_/X sky130_fd_sc_hd__buf_2
X_1572_ _1575_/A _2627_/X vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__nor2b_1
X_3311_ _3344_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3242_ _3514_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
X_3173_ _3506_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2124_ _3190_/Q _2122_/X _2053_/X _2123_/X vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__a22o_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2055_ _3238_/Q _2052_/X _2053_/X _2054_/X vssd1 vssd1 vccd1 vccd1 _3238_/D sky130_fd_sc_hd__a22o_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2957_ _3408_/Q _3404_/Q _3412_/Q _3384_/Q _2610_/S _1700_/B vssd1 vssd1 vccd1 vccd1
+ _2957_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2888_ _2467_/X _2648_/X _2649_/X _2473_/X _3000_/S0 _2575_/S vssd1 vssd1 vccd1 vccd1
+ _2888_/X sky130_fd_sc_hd__mux4_2
X_1908_ _3323_/Q _1906_/X _1645_/X _1907_/X vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__a22o_1
X_1839_ _3367_/Q _1837_/X _1656_/X _1838_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3509_ _3509_/CLK _3509_/D vssd1 vssd1 vccd1 vccd1 _3509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater381 _3475_/Q vssd1 vssd1 vccd1 vccd1 _2851_/S0 sky130_fd_sc_hd__clkbuf_16
XFILLER_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater392 _2609_/S vssd1 vssd1 vccd1 vccd1 _2595_/S sky130_fd_sc_hd__buf_8
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput151 io_b_dat_o_7[4] vssd1 vssd1 vccd1 vccd1 _2947_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput162 io_b_dat_o_8[14] vssd1 vssd1 vccd1 vccd1 _2579_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput140 io_b_dat_o_6[9] vssd1 vssd1 vccd1 vccd1 _2887_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput184 io_b_dat_o_9[5] vssd1 vssd1 vccd1 vccd1 _2600_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput173 io_b_dat_o_9[0] vssd1 vssd1 vccd1 vccd1 _2610_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput195 io_dat_i[14] vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2811_ _3021_/Q _3013_/Q _3005_/Q _3277_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2811_/X sky130_fd_sc_hd__mux4_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ _2738_/X _2739_/X _2740_/X _2741_/X _2752_/S0 _2837_/X vssd1 vssd1 vccd1 vccd1
+ _2742_/X sky130_fd_sc_hd__mux4_2
X_2673_ _3499_/Q _2966_/X _2683_/S vssd1 vssd1 vccd1 vccd1 _2673_/X sky130_fd_sc_hd__mux2_1
X_1624_ _2485_/A _2611_/S vssd1 vssd1 vccd1 vccd1 _2300_/C sky130_fd_sc_hd__or2_2
X_1555_ _1555_/A vssd1 vssd1 vccd1 vccd1 _1592_/A sky130_fd_sc_hd__clkbuf_2
X_1486_ _3518_/Q _3500_/Q _3518_/Q _3500_/Q vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__a2bb2oi_1
X_3225_ _3372_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3156_ _3180_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3087_ _3087_/CLK _3087_/D vssd1 vssd1 vccd1 vccd1 _3087_/Q sky130_fd_sc_hd__dfxtp_1
X_2107_ _2122_/A vssd1 vssd1 vccd1 vccd1 _2107_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _2038_/A vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__buf_2
XFILLER_23_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3010_ _3273_/CLK _3010_/D vssd1 vssd1 vccd1 vccd1 _3010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2725_ _3240_/Q _3216_/Q _3288_/Q _3264_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2725_/X sky130_fd_sc_hd__mux4_2
X_2656_ _2907_/X _2908_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2656_/X sky130_fd_sc_hd__mux2_1
X_1607_ _1609_/A _2974_/X vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__and2_1
X_2587_ _2587_/A0 _2587_/A1 _2644_/S vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__mux2_1
X_1538_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__inv_2
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3208_ _3372_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3139_ _3333_/CLK _3139_/D vssd1 vssd1 vccd1 vccd1 _3139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3490_ _3518_/CLK _3490_/D vssd1 vssd1 vccd1 vccd1 _3490_/Q sky130_fd_sc_hd__dfxtp_1
X_2510_ _3376_/Q vssd1 vssd1 vccd1 vccd1 _2510_/Y sky130_fd_sc_hd__inv_2
X_2441_ _3363_/Q vssd1 vssd1 vccd1 vccd1 _2441_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2372_ _3036_/Q _2367_/X _2334_/X _2368_/X vssd1 vssd1 vccd1 vccd1 _3036_/D sky130_fd_sc_hd__a22o_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2708_ _3045_/Q _3349_/Q _3093_/Q _3069_/Q _2710_/S0 _2716_/S1 vssd1 vssd1 vccd1
+ vccd1 _2708_/X sky130_fd_sc_hd__mux4_2
X_2639_ _2859_/X _2860_/X _2660_/S vssd1 vssd1 vccd1 vccd1 _2639_/X sky130_fd_sc_hd__mux2_1
Xoutput296 _2554_/Y vssd1 vssd1 vccd1 vccd1 io_ack_o sky130_fd_sc_hd__clkbuf_2
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_3 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2990_ _3185_/Q _3433_/Q _3137_/Q _3113_/Q _2991_/S0 _2991_/S1 vssd1 vssd1 vccd1
+ vccd1 _2990_/X sky130_fd_sc_hd__mux4_1
X_1941_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1941_/X sky130_fd_sc_hd__buf_2
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1872_ _2342_/D vssd1 vssd1 vccd1 vccd1 _1995_/A sky130_fd_sc_hd__buf_1
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3473_ _3474_/CLK _3473_/D vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfxtp_1
X_2424_ _2429_/A _2424_/B vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__and2_1
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2355_ _3049_/Q _2351_/X _2332_/X _2352_/X vssd1 vssd1 vccd1 vccd1 _3049_/D sky130_fd_sc_hd__a22o_1
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2286_ _3092_/Q _2282_/X _2126_/X _2283_/X vssd1 vssd1 vccd1 vccd1 _3092_/D sky130_fd_sc_hd__a22o_1
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2140_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2140_/X sky130_fd_sc_hd__buf_2
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _3225_/Q _2063_/A _2056_/X _2064_/A vssd1 vssd1 vccd1 vccd1 _3225_/D sky130_fd_sc_hd__a22o_1
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2973_ _2973_/A0 _2973_/A1 _2973_/A2 _2973_/A3 _2606_/S _2609_/S vssd1 vssd1 vccd1
+ vccd1 _2973_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _1945_/A vssd1 vssd1 vccd1 vccd1 _1924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1855_ _3357_/Q _1849_/X _1638_/X _1851_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__a22o_1
X_1786_ _3391_/Q _1782_/X _1774_/X _1784_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__a22o_1
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3456_ _3456_/CLK _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfxtp_1
X_2407_ _2407_/A vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__buf_2
X_3387_ _3423_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
X_2338_ _2563_/A vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__clkbuf_2
X_2269_ _2283_/A vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _3340_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _2569_/A vssd1 vssd1 vccd1 vccd1 _2038_/A sky130_fd_sc_hd__clkbuf_2
X_1571_ _1575_/A _2626_/X vssd1 vssd1 vccd1 vccd1 _3489_/D sky130_fd_sc_hd__nor2b_1
XFILLER_6_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3310_ _3344_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_1
X_3241_ _3307_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _3445_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
X_2123_ _2123_/A vssd1 vssd1 vccd1 vccd1 _2123_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2054_ _2054_/A vssd1 vssd1 vccd1 vccd1 _2054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _3424_/Q _3364_/Q _3400_/Q _3396_/Q _2996_/S0 _2611_/S vssd1 vssd1 vccd1 vccd1
+ _2956_/X sky130_fd_sc_hd__mux4_1
X_2887_ _2887_/A0 _2887_/A1 _2887_/A2 _2887_/A3 _2594_/S _2595_/S vssd1 vssd1 vccd1
+ vccd1 _2887_/X sky130_fd_sc_hd__mux4_1
X_1907_ _1914_/A vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__clkbuf_2
X_1838_ _1838_/A vssd1 vssd1 vccd1 vccd1 _1838_/X sky130_fd_sc_hd__buf_2
X_1769_ _2377_/A vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__clkbuf_2
X_3508_ _3509_/CLK _3508_/D vssd1 vssd1 vccd1 vccd1 _3508_/Q sky130_fd_sc_hd__dfxtp_1
X_3439_ _3439_/CLK _3439_/D vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater393 _2611_/S vssd1 vssd1 vccd1 vccd1 _2609_/S sky130_fd_sc_hd__buf_8
Xrepeater382 _2575_/X vssd1 vssd1 vccd1 vccd1 _3000_/S0 sky130_fd_sc_hd__buf_12
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput130 io_b_dat_o_6[14] vssd1 vssd1 vccd1 vccd1 _2857_/A2 sky130_fd_sc_hd__clkbuf_1
Xinput152 io_b_dat_o_7[5] vssd1 vssd1 vccd1 vccd1 _2934_/A3 sky130_fd_sc_hd__clkbuf_1
Xinput163 io_b_dat_o_8[15] vssd1 vssd1 vccd1 vccd1 _2576_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput141 io_b_dat_o_7[0] vssd1 vssd1 vccd1 vccd1 _2999_/A3 sky130_fd_sc_hd__clkbuf_1
XFILLER_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput174 io_b_dat_o_9[10] vssd1 vssd1 vccd1 vccd1 _2590_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput185 io_b_dat_o_9[6] vssd1 vssd1 vccd1 vccd1 _2598_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput196 io_dat_i[15] vssd1 vssd1 vccd1 vccd1 _2573_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2810_ _3085_/Q _3369_/Q _3037_/Q _3029_/Q _3475_/Q _3476_/Q vssd1 vssd1 vccd1 vccd1
+ _2810_/X sky130_fd_sc_hd__mux4_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _3323_/Q _3307_/Q _3171_/Q _3339_/Q _2751_/S0 _2751_/S1 vssd1 vssd1 vccd1
+ vccd1 _2741_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2672_ _2959_/X _2960_/X _2684_/S vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1623_ _1689_/A vssd1 vssd1 vccd1 vccd1 _2485_/A sky130_fd_sc_hd__clkbuf_4
X_1554_ _2564_/A vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__clkbuf_2
X_1485_ _3519_/Q vssd1 vssd1 vccd1 vccd1 _1485_/Y sky130_fd_sc_hd__inv_2
X_3224_ _3294_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
.ends

