VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cic_block
  CLASS BLOCK ;
  FOREIGN cic_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 170.000 BY 280.000 ;
  PIN io_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 -4.000 34.870 4.000 ;
    END
  END io_adr_i[0]
  PIN io_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 -4.000 42.690 4.000 ;
    END
  END io_adr_i[1]
  PIN io_cs_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 -4.000 19.230 4.000 ;
    END
  END io_cs_i
  PIN io_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 -4.000 50.050 4.000 ;
    END
  END io_dat_i[0]
  PIN io_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 -4.000 127.790 4.000 ;
    END
  END io_dat_i[10]
  PIN io_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 -4.000 135.150 4.000 ;
    END
  END io_dat_i[11]
  PIN io_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 -4.000 142.970 4.000 ;
    END
  END io_dat_i[12]
  PIN io_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 -4.000 150.790 4.000 ;
    END
  END io_dat_i[13]
  PIN io_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 -4.000 158.610 4.000 ;
    END
  END io_dat_i[14]
  PIN io_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 -4.000 166.430 4.000 ;
    END
  END io_dat_i[15]
  PIN io_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 -4.000 57.870 4.000 ;
    END
  END io_dat_i[1]
  PIN io_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 -4.000 65.690 4.000 ;
    END
  END io_dat_i[2]
  PIN io_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END io_dat_i[3]
  PIN io_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 -4.000 81.330 4.000 ;
    END
  END io_dat_i[4]
  PIN io_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 -4.000 89.150 4.000 ;
    END
  END io_dat_i[5]
  PIN io_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 -4.000 96.510 4.000 ;
    END
  END io_dat_i[6]
  PIN io_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 -4.000 104.330 4.000 ;
    END
  END io_dat_i[7]
  PIN io_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 -4.000 112.150 4.000 ;
    END
  END io_dat_i[8]
  PIN io_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 -4.000 119.970 4.000 ;
    END
  END io_dat_i[9]
  PIN io_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 276.000 5.430 284.000 ;
    END
  END io_dat_o[0]
  PIN io_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 276.000 111.690 284.000 ;
    END
  END io_dat_o[10]
  PIN io_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 276.000 122.270 284.000 ;
    END
  END io_dat_o[11]
  PIN io_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 276.000 132.850 284.000 ;
    END
  END io_dat_o[12]
  PIN io_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 276.000 143.430 284.000 ;
    END
  END io_dat_o[13]
  PIN io_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 276.000 154.010 284.000 ;
    END
  END io_dat_o[14]
  PIN io_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 276.000 164.590 284.000 ;
    END
  END io_dat_o[15]
  PIN io_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 276.000 16.010 284.000 ;
    END
  END io_dat_o[1]
  PIN io_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 276.000 26.590 284.000 ;
    END
  END io_dat_o[2]
  PIN io_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 276.000 37.170 284.000 ;
    END
  END io_dat_o[3]
  PIN io_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 276.000 47.750 284.000 ;
    END
  END io_dat_o[4]
  PIN io_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 276.000 58.330 284.000 ;
    END
  END io_dat_o[5]
  PIN io_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 276.000 68.910 284.000 ;
    END
  END io_dat_o[6]
  PIN io_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 276.000 79.490 284.000 ;
    END
  END io_dat_o[7]
  PIN io_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 276.000 90.530 284.000 ;
    END
  END io_dat_o[8]
  PIN io_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 276.000 101.110 284.000 ;
    END
  END io_dat_o[9]
  PIN io_eo[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 146.240 174.000 146.840 ;
    END
  END io_eo[0]
  PIN io_eo[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 166.640 174.000 167.240 ;
    END
  END io_eo[10]
  PIN io_eo[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 168.680 174.000 169.280 ;
    END
  END io_eo[11]
  PIN io_eo[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 170.720 174.000 171.320 ;
    END
  END io_eo[12]
  PIN io_eo[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 172.760 174.000 173.360 ;
    END
  END io_eo[13]
  PIN io_eo[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 174.800 174.000 175.400 ;
    END
  END io_eo[14]
  PIN io_eo[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 176.840 174.000 177.440 ;
    END
  END io_eo[15]
  PIN io_eo[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 178.880 174.000 179.480 ;
    END
  END io_eo[16]
  PIN io_eo[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 180.920 174.000 181.520 ;
    END
  END io_eo[17]
  PIN io_eo[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 182.960 174.000 183.560 ;
    END
  END io_eo[18]
  PIN io_eo[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 185.000 174.000 185.600 ;
    END
  END io_eo[19]
  PIN io_eo[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 148.280 174.000 148.880 ;
    END
  END io_eo[1]
  PIN io_eo[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 187.040 174.000 187.640 ;
    END
  END io_eo[20]
  PIN io_eo[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 189.080 174.000 189.680 ;
    END
  END io_eo[21]
  PIN io_eo[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 191.120 174.000 191.720 ;
    END
  END io_eo[22]
  PIN io_eo[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 193.160 174.000 193.760 ;
    END
  END io_eo[23]
  PIN io_eo[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 195.200 174.000 195.800 ;
    END
  END io_eo[24]
  PIN io_eo[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 197.240 174.000 197.840 ;
    END
  END io_eo[25]
  PIN io_eo[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 199.280 174.000 199.880 ;
    END
  END io_eo[26]
  PIN io_eo[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 201.320 174.000 201.920 ;
    END
  END io_eo[27]
  PIN io_eo[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 203.360 174.000 203.960 ;
    END
  END io_eo[28]
  PIN io_eo[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 205.400 174.000 206.000 ;
    END
  END io_eo[29]
  PIN io_eo[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 150.320 174.000 150.920 ;
    END
  END io_eo[2]
  PIN io_eo[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 207.440 174.000 208.040 ;
    END
  END io_eo[30]
  PIN io_eo[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 209.480 174.000 210.080 ;
    END
  END io_eo[31]
  PIN io_eo[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 211.520 174.000 212.120 ;
    END
  END io_eo[32]
  PIN io_eo[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 213.560 174.000 214.160 ;
    END
  END io_eo[33]
  PIN io_eo[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 215.600 174.000 216.200 ;
    END
  END io_eo[34]
  PIN io_eo[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 217.640 174.000 218.240 ;
    END
  END io_eo[35]
  PIN io_eo[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 219.680 174.000 220.280 ;
    END
  END io_eo[36]
  PIN io_eo[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 221.720 174.000 222.320 ;
    END
  END io_eo[37]
  PIN io_eo[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 223.760 174.000 224.360 ;
    END
  END io_eo[38]
  PIN io_eo[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 225.800 174.000 226.400 ;
    END
  END io_eo[39]
  PIN io_eo[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 152.360 174.000 152.960 ;
    END
  END io_eo[3]
  PIN io_eo[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 227.840 174.000 228.440 ;
    END
  END io_eo[40]
  PIN io_eo[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 229.880 174.000 230.480 ;
    END
  END io_eo[41]
  PIN io_eo[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 231.920 174.000 232.520 ;
    END
  END io_eo[42]
  PIN io_eo[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 233.960 174.000 234.560 ;
    END
  END io_eo[43]
  PIN io_eo[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 236.000 174.000 236.600 ;
    END
  END io_eo[44]
  PIN io_eo[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 238.040 174.000 238.640 ;
    END
  END io_eo[45]
  PIN io_eo[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 240.080 174.000 240.680 ;
    END
  END io_eo[46]
  PIN io_eo[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 242.120 174.000 242.720 ;
    END
  END io_eo[47]
  PIN io_eo[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 244.160 174.000 244.760 ;
    END
  END io_eo[48]
  PIN io_eo[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 246.200 174.000 246.800 ;
    END
  END io_eo[49]
  PIN io_eo[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 154.400 174.000 155.000 ;
    END
  END io_eo[4]
  PIN io_eo[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 248.240 174.000 248.840 ;
    END
  END io_eo[50]
  PIN io_eo[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 250.280 174.000 250.880 ;
    END
  END io_eo[51]
  PIN io_eo[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 252.320 174.000 252.920 ;
    END
  END io_eo[52]
  PIN io_eo[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 254.360 174.000 254.960 ;
    END
  END io_eo[53]
  PIN io_eo[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 256.400 174.000 257.000 ;
    END
  END io_eo[54]
  PIN io_eo[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 258.440 174.000 259.040 ;
    END
  END io_eo[55]
  PIN io_eo[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 260.480 174.000 261.080 ;
    END
  END io_eo[56]
  PIN io_eo[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 262.520 174.000 263.120 ;
    END
  END io_eo[57]
  PIN io_eo[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 264.560 174.000 265.160 ;
    END
  END io_eo[58]
  PIN io_eo[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 266.600 174.000 267.200 ;
    END
  END io_eo[59]
  PIN io_eo[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 156.440 174.000 157.040 ;
    END
  END io_eo[5]
  PIN io_eo[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 268.640 174.000 269.240 ;
    END
  END io_eo[60]
  PIN io_eo[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 270.680 174.000 271.280 ;
    END
  END io_eo[61]
  PIN io_eo[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 272.720 174.000 273.320 ;
    END
  END io_eo[62]
  PIN io_eo[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 274.760 174.000 275.360 ;
    END
  END io_eo[63]
  PIN io_eo[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 158.480 174.000 159.080 ;
    END
  END io_eo[6]
  PIN io_eo[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 160.520 174.000 161.120 ;
    END
  END io_eo[7]
  PIN io_eo[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 162.560 174.000 163.160 ;
    END
  END io_eo[8]
  PIN io_eo[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 164.600 174.000 165.200 ;
    END
  END io_eo[9]
  PIN io_i_0_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 0.720 4.000 1.320 ;
    END
  END io_i_0_ci
  PIN io_i_0_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 17.040 4.000 17.640 ;
    END
  END io_i_0_in1[0]
  PIN io_i_0_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 33.360 4.000 33.960 ;
    END
  END io_i_0_in1[1]
  PIN io_i_0_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 49.680 4.000 50.280 ;
    END
  END io_i_0_in1[2]
  PIN io_i_0_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 66.000 4.000 66.600 ;
    END
  END io_i_0_in1[3]
  PIN io_i_0_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 82.320 4.000 82.920 ;
    END
  END io_i_0_in1[4]
  PIN io_i_0_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 98.640 4.000 99.240 ;
    END
  END io_i_0_in1[5]
  PIN io_i_0_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 114.960 4.000 115.560 ;
    END
  END io_i_0_in1[6]
  PIN io_i_0_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 131.280 4.000 131.880 ;
    END
  END io_i_0_in1[7]
  PIN io_i_1_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.760 4.000 3.360 ;
    END
  END io_i_1_ci
  PIN io_i_1_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 19.080 4.000 19.680 ;
    END
  END io_i_1_in1[0]
  PIN io_i_1_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 35.400 4.000 36.000 ;
    END
  END io_i_1_in1[1]
  PIN io_i_1_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 51.720 4.000 52.320 ;
    END
  END io_i_1_in1[2]
  PIN io_i_1_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.040 4.000 68.640 ;
    END
  END io_i_1_in1[3]
  PIN io_i_1_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.360 4.000 84.960 ;
    END
  END io_i_1_in1[4]
  PIN io_i_1_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.680 4.000 101.280 ;
    END
  END io_i_1_in1[5]
  PIN io_i_1_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 117.000 4.000 117.600 ;
    END
  END io_i_1_in1[6]
  PIN io_i_1_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 133.320 4.000 133.920 ;
    END
  END io_i_1_in1[7]
  PIN io_i_2_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.800 4.000 5.400 ;
    END
  END io_i_2_ci
  PIN io_i_2_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 21.120 4.000 21.720 ;
    END
  END io_i_2_in1[0]
  PIN io_i_2_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 37.440 4.000 38.040 ;
    END
  END io_i_2_in1[1]
  PIN io_i_2_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 53.760 4.000 54.360 ;
    END
  END io_i_2_in1[2]
  PIN io_i_2_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 70.080 4.000 70.680 ;
    END
  END io_i_2_in1[3]
  PIN io_i_2_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 86.400 4.000 87.000 ;
    END
  END io_i_2_in1[4]
  PIN io_i_2_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 102.720 4.000 103.320 ;
    END
  END io_i_2_in1[5]
  PIN io_i_2_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 119.040 4.000 119.640 ;
    END
  END io_i_2_in1[6]
  PIN io_i_2_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 135.360 4.000 135.960 ;
    END
  END io_i_2_in1[7]
  PIN io_i_3_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.840 4.000 7.440 ;
    END
  END io_i_3_ci
  PIN io_i_3_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 23.160 4.000 23.760 ;
    END
  END io_i_3_in1[0]
  PIN io_i_3_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 39.480 4.000 40.080 ;
    END
  END io_i_3_in1[1]
  PIN io_i_3_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 55.800 4.000 56.400 ;
    END
  END io_i_3_in1[2]
  PIN io_i_3_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.120 4.000 72.720 ;
    END
  END io_i_3_in1[3]
  PIN io_i_3_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.440 4.000 89.040 ;
    END
  END io_i_3_in1[4]
  PIN io_i_3_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.760 4.000 105.360 ;
    END
  END io_i_3_in1[5]
  PIN io_i_3_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 121.080 4.000 121.680 ;
    END
  END io_i_3_in1[6]
  PIN io_i_3_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 137.400 4.000 138.000 ;
    END
  END io_i_3_in1[7]
  PIN io_i_4_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.880 4.000 9.480 ;
    END
  END io_i_4_ci
  PIN io_i_4_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 25.200 4.000 25.800 ;
    END
  END io_i_4_in1[0]
  PIN io_i_4_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 41.520 4.000 42.120 ;
    END
  END io_i_4_in1[1]
  PIN io_i_4_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 57.840 4.000 58.440 ;
    END
  END io_i_4_in1[2]
  PIN io_i_4_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 74.160 4.000 74.760 ;
    END
  END io_i_4_in1[3]
  PIN io_i_4_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 90.480 4.000 91.080 ;
    END
  END io_i_4_in1[4]
  PIN io_i_4_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 106.800 4.000 107.400 ;
    END
  END io_i_4_in1[5]
  PIN io_i_4_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 123.120 4.000 123.720 ;
    END
  END io_i_4_in1[6]
  PIN io_i_4_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 139.440 4.000 140.040 ;
    END
  END io_i_4_in1[7]
  PIN io_i_5_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.920 4.000 11.520 ;
    END
  END io_i_5_ci
  PIN io_i_5_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 27.240 4.000 27.840 ;
    END
  END io_i_5_in1[0]
  PIN io_i_5_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 43.560 4.000 44.160 ;
    END
  END io_i_5_in1[1]
  PIN io_i_5_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 59.880 4.000 60.480 ;
    END
  END io_i_5_in1[2]
  PIN io_i_5_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.200 4.000 76.800 ;
    END
  END io_i_5_in1[3]
  PIN io_i_5_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.520 4.000 93.120 ;
    END
  END io_i_5_in1[4]
  PIN io_i_5_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.840 4.000 109.440 ;
    END
  END io_i_5_in1[5]
  PIN io_i_5_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 125.160 4.000 125.760 ;
    END
  END io_i_5_in1[6]
  PIN io_i_5_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 141.480 4.000 142.080 ;
    END
  END io_i_5_in1[7]
  PIN io_i_6_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.960 4.000 13.560 ;
    END
  END io_i_6_ci
  PIN io_i_6_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 29.280 4.000 29.880 ;
    END
  END io_i_6_in1[0]
  PIN io_i_6_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 45.600 4.000 46.200 ;
    END
  END io_i_6_in1[1]
  PIN io_i_6_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 61.920 4.000 62.520 ;
    END
  END io_i_6_in1[2]
  PIN io_i_6_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 78.240 4.000 78.840 ;
    END
  END io_i_6_in1[3]
  PIN io_i_6_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 94.560 4.000 95.160 ;
    END
  END io_i_6_in1[4]
  PIN io_i_6_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 110.880 4.000 111.480 ;
    END
  END io_i_6_in1[5]
  PIN io_i_6_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 127.200 4.000 127.800 ;
    END
  END io_i_6_in1[6]
  PIN io_i_6_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 143.520 4.000 144.120 ;
    END
  END io_i_6_in1[7]
  PIN io_i_7_ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 15.000 4.000 15.600 ;
    END
  END io_i_7_ci
  PIN io_i_7_in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 31.320 4.000 31.920 ;
    END
  END io_i_7_in1[0]
  PIN io_i_7_in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 47.640 4.000 48.240 ;
    END
  END io_i_7_in1[1]
  PIN io_i_7_in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 63.960 4.000 64.560 ;
    END
  END io_i_7_in1[2]
  PIN io_i_7_in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.280 4.000 80.880 ;
    END
  END io_i_7_in1[3]
  PIN io_i_7_in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.600 4.000 97.200 ;
    END
  END io_i_7_in1[4]
  PIN io_i_7_in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.920 4.000 113.520 ;
    END
  END io_i_7_in1[5]
  PIN io_i_7_in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 129.240 4.000 129.840 ;
    END
  END io_i_7_in1[6]
  PIN io_i_7_in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 145.560 4.000 146.160 ;
    END
  END io_i_7_in1[7]
  PIN io_o_0_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 0.720 174.000 1.320 ;
    END
  END io_o_0_co
  PIN io_o_0_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 16.360 174.000 16.960 ;
    END
  END io_o_0_out[0]
  PIN io_o_0_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 32.680 174.000 33.280 ;
    END
  END io_o_0_out[1]
  PIN io_o_0_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 49.000 174.000 49.600 ;
    END
  END io_o_0_out[2]
  PIN io_o_0_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 65.320 174.000 65.920 ;
    END
  END io_o_0_out[3]
  PIN io_o_0_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 81.640 174.000 82.240 ;
    END
  END io_o_0_out[4]
  PIN io_o_0_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 97.960 174.000 98.560 ;
    END
  END io_o_0_out[5]
  PIN io_o_0_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 114.280 174.000 114.880 ;
    END
  END io_o_0_out[6]
  PIN io_o_0_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 130.600 174.000 131.200 ;
    END
  END io_o_0_out[7]
  PIN io_o_1_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 2.080 174.000 2.680 ;
    END
  END io_o_1_co
  PIN io_o_1_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 18.400 174.000 19.000 ;
    END
  END io_o_1_out[0]
  PIN io_o_1_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 34.720 174.000 35.320 ;
    END
  END io_o_1_out[1]
  PIN io_o_1_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 51.040 174.000 51.640 ;
    END
  END io_o_1_out[2]
  PIN io_o_1_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 67.360 174.000 67.960 ;
    END
  END io_o_1_out[3]
  PIN io_o_1_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 83.680 174.000 84.280 ;
    END
  END io_o_1_out[4]
  PIN io_o_1_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 100.000 174.000 100.600 ;
    END
  END io_o_1_out[5]
  PIN io_o_1_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 116.320 174.000 116.920 ;
    END
  END io_o_1_out[6]
  PIN io_o_1_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 132.640 174.000 133.240 ;
    END
  END io_o_1_out[7]
  PIN io_o_2_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 4.120 174.000 4.720 ;
    END
  END io_o_2_co
  PIN io_o_2_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 20.440 174.000 21.040 ;
    END
  END io_o_2_out[0]
  PIN io_o_2_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 36.760 174.000 37.360 ;
    END
  END io_o_2_out[1]
  PIN io_o_2_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 53.080 174.000 53.680 ;
    END
  END io_o_2_out[2]
  PIN io_o_2_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 69.400 174.000 70.000 ;
    END
  END io_o_2_out[3]
  PIN io_o_2_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 85.720 174.000 86.320 ;
    END
  END io_o_2_out[4]
  PIN io_o_2_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 102.040 174.000 102.640 ;
    END
  END io_o_2_out[5]
  PIN io_o_2_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 118.360 174.000 118.960 ;
    END
  END io_o_2_out[6]
  PIN io_o_2_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 134.680 174.000 135.280 ;
    END
  END io_o_2_out[7]
  PIN io_o_3_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 6.160 174.000 6.760 ;
    END
  END io_o_3_co
  PIN io_o_3_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 22.480 174.000 23.080 ;
    END
  END io_o_3_out[0]
  PIN io_o_3_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 38.800 174.000 39.400 ;
    END
  END io_o_3_out[1]
  PIN io_o_3_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 55.120 174.000 55.720 ;
    END
  END io_o_3_out[2]
  PIN io_o_3_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 71.440 174.000 72.040 ;
    END
  END io_o_3_out[3]
  PIN io_o_3_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 87.760 174.000 88.360 ;
    END
  END io_o_3_out[4]
  PIN io_o_3_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 104.080 174.000 104.680 ;
    END
  END io_o_3_out[5]
  PIN io_o_3_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 120.400 174.000 121.000 ;
    END
  END io_o_3_out[6]
  PIN io_o_3_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 136.720 174.000 137.320 ;
    END
  END io_o_3_out[7]
  PIN io_o_4_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 8.200 174.000 8.800 ;
    END
  END io_o_4_co
  PIN io_o_4_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 24.520 174.000 25.120 ;
    END
  END io_o_4_out[0]
  PIN io_o_4_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 40.840 174.000 41.440 ;
    END
  END io_o_4_out[1]
  PIN io_o_4_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 57.160 174.000 57.760 ;
    END
  END io_o_4_out[2]
  PIN io_o_4_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 73.480 174.000 74.080 ;
    END
  END io_o_4_out[3]
  PIN io_o_4_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 89.800 174.000 90.400 ;
    END
  END io_o_4_out[4]
  PIN io_o_4_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 106.120 174.000 106.720 ;
    END
  END io_o_4_out[5]
  PIN io_o_4_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 122.440 174.000 123.040 ;
    END
  END io_o_4_out[6]
  PIN io_o_4_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 138.760 174.000 139.360 ;
    END
  END io_o_4_out[7]
  PIN io_o_5_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 10.240 174.000 10.840 ;
    END
  END io_o_5_co
  PIN io_o_5_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 26.560 174.000 27.160 ;
    END
  END io_o_5_out[0]
  PIN io_o_5_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 42.880 174.000 43.480 ;
    END
  END io_o_5_out[1]
  PIN io_o_5_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 59.200 174.000 59.800 ;
    END
  END io_o_5_out[2]
  PIN io_o_5_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 75.520 174.000 76.120 ;
    END
  END io_o_5_out[3]
  PIN io_o_5_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 91.840 174.000 92.440 ;
    END
  END io_o_5_out[4]
  PIN io_o_5_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 108.160 174.000 108.760 ;
    END
  END io_o_5_out[5]
  PIN io_o_5_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 124.480 174.000 125.080 ;
    END
  END io_o_5_out[6]
  PIN io_o_5_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 140.800 174.000 141.400 ;
    END
  END io_o_5_out[7]
  PIN io_o_6_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 12.280 174.000 12.880 ;
    END
  END io_o_6_co
  PIN io_o_6_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 28.600 174.000 29.200 ;
    END
  END io_o_6_out[0]
  PIN io_o_6_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 44.920 174.000 45.520 ;
    END
  END io_o_6_out[1]
  PIN io_o_6_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 61.240 174.000 61.840 ;
    END
  END io_o_6_out[2]
  PIN io_o_6_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 77.560 174.000 78.160 ;
    END
  END io_o_6_out[3]
  PIN io_o_6_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 93.880 174.000 94.480 ;
    END
  END io_o_6_out[4]
  PIN io_o_6_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 110.200 174.000 110.800 ;
    END
  END io_o_6_out[5]
  PIN io_o_6_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 126.520 174.000 127.120 ;
    END
  END io_o_6_out[6]
  PIN io_o_6_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 142.160 174.000 142.760 ;
    END
  END io_o_6_out[7]
  PIN io_o_7_co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 14.320 174.000 14.920 ;
    END
  END io_o_7_co
  PIN io_o_7_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 30.640 174.000 31.240 ;
    END
  END io_o_7_out[0]
  PIN io_o_7_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 46.960 174.000 47.560 ;
    END
  END io_o_7_out[1]
  PIN io_o_7_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 63.280 174.000 63.880 ;
    END
  END io_o_7_out[2]
  PIN io_o_7_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 79.600 174.000 80.200 ;
    END
  END io_o_7_out[3]
  PIN io_o_7_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 95.920 174.000 96.520 ;
    END
  END io_o_7_out[4]
  PIN io_o_7_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 112.240 174.000 112.840 ;
    END
  END io_o_7_out[5]
  PIN io_o_7_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 128.560 174.000 129.160 ;
    END
  END io_o_7_out[6]
  PIN io_o_7_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 144.200 174.000 144.800 ;
    END
  END io_o_7_out[7]
  PIN io_vci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 -4.000 4.050 4.000 ;
    END
  END io_vci
  PIN io_vco
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 -4.000 11.410 4.000 ;
    END
  END io_vco
  PIN io_vi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 276.800 174.000 277.400 ;
    END
  END io_vi
  PIN io_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 -4.000 27.050 4.000 ;
    END
  END io_we_i
  PIN io_wo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 147.600 4.000 148.200 ;
    END
  END io_wo[0]
  PIN io_wo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.000 4.000 168.600 ;
    END
  END io_wo[10]
  PIN io_wo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 170.040 4.000 170.640 ;
    END
  END io_wo[11]
  PIN io_wo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.080 4.000 172.680 ;
    END
  END io_wo[12]
  PIN io_wo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 174.120 4.000 174.720 ;
    END
  END io_wo[13]
  PIN io_wo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.160 4.000 176.760 ;
    END
  END io_wo[14]
  PIN io_wo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 178.200 4.000 178.800 ;
    END
  END io_wo[15]
  PIN io_wo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.240 4.000 180.840 ;
    END
  END io_wo[16]
  PIN io_wo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 182.280 4.000 182.880 ;
    END
  END io_wo[17]
  PIN io_wo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 184.320 4.000 184.920 ;
    END
  END io_wo[18]
  PIN io_wo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 186.360 4.000 186.960 ;
    END
  END io_wo[19]
  PIN io_wo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 149.640 4.000 150.240 ;
    END
  END io_wo[1]
  PIN io_wo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 188.400 4.000 189.000 ;
    END
  END io_wo[20]
  PIN io_wo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 190.440 4.000 191.040 ;
    END
  END io_wo[21]
  PIN io_wo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 192.480 4.000 193.080 ;
    END
  END io_wo[22]
  PIN io_wo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 194.520 4.000 195.120 ;
    END
  END io_wo[23]
  PIN io_wo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 196.560 4.000 197.160 ;
    END
  END io_wo[24]
  PIN io_wo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 198.600 4.000 199.200 ;
    END
  END io_wo[25]
  PIN io_wo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.640 4.000 201.240 ;
    END
  END io_wo[26]
  PIN io_wo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 202.680 4.000 203.280 ;
    END
  END io_wo[27]
  PIN io_wo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.720 4.000 205.320 ;
    END
  END io_wo[28]
  PIN io_wo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 206.760 4.000 207.360 ;
    END
  END io_wo[29]
  PIN io_wo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 151.680 4.000 152.280 ;
    END
  END io_wo[2]
  PIN io_wo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.800 4.000 209.400 ;
    END
  END io_wo[30]
  PIN io_wo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 210.840 4.000 211.440 ;
    END
  END io_wo[31]
  PIN io_wo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.880 4.000 213.480 ;
    END
  END io_wo[32]
  PIN io_wo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 214.920 4.000 215.520 ;
    END
  END io_wo[33]
  PIN io_wo[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.960 4.000 217.560 ;
    END
  END io_wo[34]
  PIN io_wo[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 219.000 4.000 219.600 ;
    END
  END io_wo[35]
  PIN io_wo[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 221.040 4.000 221.640 ;
    END
  END io_wo[36]
  PIN io_wo[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 223.080 4.000 223.680 ;
    END
  END io_wo[37]
  PIN io_wo[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 225.120 4.000 225.720 ;
    END
  END io_wo[38]
  PIN io_wo[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 227.160 4.000 227.760 ;
    END
  END io_wo[39]
  PIN io_wo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 153.720 4.000 154.320 ;
    END
  END io_wo[3]
  PIN io_wo[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 229.200 4.000 229.800 ;
    END
  END io_wo[40]
  PIN io_wo[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 231.240 4.000 231.840 ;
    END
  END io_wo[41]
  PIN io_wo[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 233.280 4.000 233.880 ;
    END
  END io_wo[42]
  PIN io_wo[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 235.320 4.000 235.920 ;
    END
  END io_wo[43]
  PIN io_wo[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 237.360 4.000 237.960 ;
    END
  END io_wo[44]
  PIN io_wo[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 239.400 4.000 240.000 ;
    END
  END io_wo[45]
  PIN io_wo[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 241.440 4.000 242.040 ;
    END
  END io_wo[46]
  PIN io_wo[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 243.480 4.000 244.080 ;
    END
  END io_wo[47]
  PIN io_wo[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 245.520 4.000 246.120 ;
    END
  END io_wo[48]
  PIN io_wo[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 247.560 4.000 248.160 ;
    END
  END io_wo[49]
  PIN io_wo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 155.760 4.000 156.360 ;
    END
  END io_wo[4]
  PIN io_wo[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 249.600 4.000 250.200 ;
    END
  END io_wo[50]
  PIN io_wo[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 251.640 4.000 252.240 ;
    END
  END io_wo[51]
  PIN io_wo[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 253.680 4.000 254.280 ;
    END
  END io_wo[52]
  PIN io_wo[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 255.720 4.000 256.320 ;
    END
  END io_wo[53]
  PIN io_wo[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 257.760 4.000 258.360 ;
    END
  END io_wo[54]
  PIN io_wo[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 259.800 4.000 260.400 ;
    END
  END io_wo[55]
  PIN io_wo[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 261.840 4.000 262.440 ;
    END
  END io_wo[56]
  PIN io_wo[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 263.880 4.000 264.480 ;
    END
  END io_wo[57]
  PIN io_wo[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 265.920 4.000 266.520 ;
    END
  END io_wo[58]
  PIN io_wo[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 267.960 4.000 268.560 ;
    END
  END io_wo[59]
  PIN io_wo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 157.800 4.000 158.400 ;
    END
  END io_wo[5]
  PIN io_wo[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 270.000 4.000 270.600 ;
    END
  END io_wo[60]
  PIN io_wo[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.040 4.000 272.640 ;
    END
  END io_wo[61]
  PIN io_wo[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 274.080 4.000 274.680 ;
    END
  END io_wo[62]
  PIN io_wo[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.120 4.000 276.720 ;
    END
  END io_wo[63]
  PIN io_wo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 159.840 4.000 160.440 ;
    END
  END io_wo[6]
  PIN io_wo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 161.880 4.000 162.480 ;
    END
  END io_wo[7]
  PIN io_wo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 163.920 4.000 164.520 ;
    END
  END io_wo[8]
  PIN io_wo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 165.960 4.000 166.560 ;
    END
  END io_wo[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 278.160 4.000 278.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 166.000 278.840 174.000 279.440 ;
    END
  END wb_rst_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 137.185 10.640 138.785 266.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 84.200 10.640 85.800 266.800 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 31.215 10.640 32.815 266.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 110.695 10.640 112.295 266.800 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 57.705 10.640 59.305 266.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 8.245 164.995 266.645 ;
      LAYER met1 ;
        RECT 3.750 6.500 166.450 273.660 ;
      LAYER met2 ;
        RECT 3.780 275.720 4.870 279.325 ;
        RECT 5.710 275.720 15.450 279.325 ;
        RECT 16.290 275.720 26.030 279.325 ;
        RECT 26.870 275.720 36.610 279.325 ;
        RECT 37.450 275.720 47.190 279.325 ;
        RECT 48.030 275.720 57.770 279.325 ;
        RECT 58.610 275.720 68.350 279.325 ;
        RECT 69.190 275.720 78.930 279.325 ;
        RECT 79.770 275.720 89.970 279.325 ;
        RECT 90.810 275.720 100.550 279.325 ;
        RECT 101.390 275.720 111.130 279.325 ;
        RECT 111.970 275.720 121.710 279.325 ;
        RECT 122.550 275.720 132.290 279.325 ;
        RECT 133.130 275.720 142.870 279.325 ;
        RECT 143.710 275.720 153.450 279.325 ;
        RECT 154.290 275.720 164.030 279.325 ;
        RECT 164.870 275.720 166.420 279.325 ;
        RECT 3.780 4.280 166.420 275.720 ;
        RECT 4.330 0.835 10.850 4.280 ;
        RECT 11.690 0.835 18.670 4.280 ;
        RECT 19.510 0.835 26.490 4.280 ;
        RECT 27.330 0.835 34.310 4.280 ;
        RECT 35.150 0.835 42.130 4.280 ;
        RECT 42.970 0.835 49.490 4.280 ;
        RECT 50.330 0.835 57.310 4.280 ;
        RECT 58.150 0.835 65.130 4.280 ;
        RECT 65.970 0.835 72.950 4.280 ;
        RECT 73.790 0.835 80.770 4.280 ;
        RECT 81.610 0.835 88.590 4.280 ;
        RECT 89.430 0.835 95.950 4.280 ;
        RECT 96.790 0.835 103.770 4.280 ;
        RECT 104.610 0.835 111.590 4.280 ;
        RECT 112.430 0.835 119.410 4.280 ;
        RECT 120.250 0.835 127.230 4.280 ;
        RECT 128.070 0.835 134.590 4.280 ;
        RECT 135.430 0.835 142.410 4.280 ;
        RECT 143.250 0.835 150.230 4.280 ;
        RECT 151.070 0.835 158.050 4.280 ;
        RECT 158.890 0.835 165.870 4.280 ;
      LAYER met3 ;
        RECT 4.000 279.160 165.600 279.305 ;
        RECT 4.400 278.440 165.600 279.160 ;
        RECT 4.400 277.800 166.000 278.440 ;
        RECT 4.400 277.760 165.600 277.800 ;
        RECT 4.000 277.120 165.600 277.760 ;
        RECT 4.400 276.400 165.600 277.120 ;
        RECT 4.400 275.760 166.000 276.400 ;
        RECT 4.400 275.720 165.600 275.760 ;
        RECT 4.000 275.080 165.600 275.720 ;
        RECT 4.400 274.360 165.600 275.080 ;
        RECT 4.400 273.720 166.000 274.360 ;
        RECT 4.400 273.680 165.600 273.720 ;
        RECT 4.000 273.040 165.600 273.680 ;
        RECT 4.400 272.320 165.600 273.040 ;
        RECT 4.400 271.680 166.000 272.320 ;
        RECT 4.400 271.640 165.600 271.680 ;
        RECT 4.000 271.000 165.600 271.640 ;
        RECT 4.400 270.280 165.600 271.000 ;
        RECT 4.400 269.640 166.000 270.280 ;
        RECT 4.400 269.600 165.600 269.640 ;
        RECT 4.000 268.960 165.600 269.600 ;
        RECT 4.400 268.240 165.600 268.960 ;
        RECT 4.400 267.600 166.000 268.240 ;
        RECT 4.400 267.560 165.600 267.600 ;
        RECT 4.000 266.920 165.600 267.560 ;
        RECT 4.400 266.200 165.600 266.920 ;
        RECT 4.400 265.560 166.000 266.200 ;
        RECT 4.400 265.520 165.600 265.560 ;
        RECT 4.000 264.880 165.600 265.520 ;
        RECT 4.400 264.160 165.600 264.880 ;
        RECT 4.400 263.520 166.000 264.160 ;
        RECT 4.400 263.480 165.600 263.520 ;
        RECT 4.000 262.840 165.600 263.480 ;
        RECT 4.400 262.120 165.600 262.840 ;
        RECT 4.400 261.480 166.000 262.120 ;
        RECT 4.400 261.440 165.600 261.480 ;
        RECT 4.000 260.800 165.600 261.440 ;
        RECT 4.400 260.080 165.600 260.800 ;
        RECT 4.400 259.440 166.000 260.080 ;
        RECT 4.400 259.400 165.600 259.440 ;
        RECT 4.000 258.760 165.600 259.400 ;
        RECT 4.400 258.040 165.600 258.760 ;
        RECT 4.400 257.400 166.000 258.040 ;
        RECT 4.400 257.360 165.600 257.400 ;
        RECT 4.000 256.720 165.600 257.360 ;
        RECT 4.400 256.000 165.600 256.720 ;
        RECT 4.400 255.360 166.000 256.000 ;
        RECT 4.400 255.320 165.600 255.360 ;
        RECT 4.000 254.680 165.600 255.320 ;
        RECT 4.400 253.960 165.600 254.680 ;
        RECT 4.400 253.320 166.000 253.960 ;
        RECT 4.400 253.280 165.600 253.320 ;
        RECT 4.000 252.640 165.600 253.280 ;
        RECT 4.400 251.920 165.600 252.640 ;
        RECT 4.400 251.280 166.000 251.920 ;
        RECT 4.400 251.240 165.600 251.280 ;
        RECT 4.000 250.600 165.600 251.240 ;
        RECT 4.400 249.880 165.600 250.600 ;
        RECT 4.400 249.240 166.000 249.880 ;
        RECT 4.400 249.200 165.600 249.240 ;
        RECT 4.000 248.560 165.600 249.200 ;
        RECT 4.400 247.840 165.600 248.560 ;
        RECT 4.400 247.200 166.000 247.840 ;
        RECT 4.400 247.160 165.600 247.200 ;
        RECT 4.000 246.520 165.600 247.160 ;
        RECT 4.400 245.800 165.600 246.520 ;
        RECT 4.400 245.160 166.000 245.800 ;
        RECT 4.400 245.120 165.600 245.160 ;
        RECT 4.000 244.480 165.600 245.120 ;
        RECT 4.400 243.760 165.600 244.480 ;
        RECT 4.400 243.120 166.000 243.760 ;
        RECT 4.400 243.080 165.600 243.120 ;
        RECT 4.000 242.440 165.600 243.080 ;
        RECT 4.400 241.720 165.600 242.440 ;
        RECT 4.400 241.080 166.000 241.720 ;
        RECT 4.400 241.040 165.600 241.080 ;
        RECT 4.000 240.400 165.600 241.040 ;
        RECT 4.400 239.680 165.600 240.400 ;
        RECT 4.400 239.040 166.000 239.680 ;
        RECT 4.400 239.000 165.600 239.040 ;
        RECT 4.000 238.360 165.600 239.000 ;
        RECT 4.400 237.640 165.600 238.360 ;
        RECT 4.400 237.000 166.000 237.640 ;
        RECT 4.400 236.960 165.600 237.000 ;
        RECT 4.000 236.320 165.600 236.960 ;
        RECT 4.400 235.600 165.600 236.320 ;
        RECT 4.400 234.960 166.000 235.600 ;
        RECT 4.400 234.920 165.600 234.960 ;
        RECT 4.000 234.280 165.600 234.920 ;
        RECT 4.400 233.560 165.600 234.280 ;
        RECT 4.400 232.920 166.000 233.560 ;
        RECT 4.400 232.880 165.600 232.920 ;
        RECT 4.000 232.240 165.600 232.880 ;
        RECT 4.400 231.520 165.600 232.240 ;
        RECT 4.400 230.880 166.000 231.520 ;
        RECT 4.400 230.840 165.600 230.880 ;
        RECT 4.000 230.200 165.600 230.840 ;
        RECT 4.400 229.480 165.600 230.200 ;
        RECT 4.400 228.840 166.000 229.480 ;
        RECT 4.400 228.800 165.600 228.840 ;
        RECT 4.000 228.160 165.600 228.800 ;
        RECT 4.400 227.440 165.600 228.160 ;
        RECT 4.400 226.800 166.000 227.440 ;
        RECT 4.400 226.760 165.600 226.800 ;
        RECT 4.000 226.120 165.600 226.760 ;
        RECT 4.400 225.400 165.600 226.120 ;
        RECT 4.400 224.760 166.000 225.400 ;
        RECT 4.400 224.720 165.600 224.760 ;
        RECT 4.000 224.080 165.600 224.720 ;
        RECT 4.400 223.360 165.600 224.080 ;
        RECT 4.400 222.720 166.000 223.360 ;
        RECT 4.400 222.680 165.600 222.720 ;
        RECT 4.000 222.040 165.600 222.680 ;
        RECT 4.400 221.320 165.600 222.040 ;
        RECT 4.400 220.680 166.000 221.320 ;
        RECT 4.400 220.640 165.600 220.680 ;
        RECT 4.000 220.000 165.600 220.640 ;
        RECT 4.400 219.280 165.600 220.000 ;
        RECT 4.400 218.640 166.000 219.280 ;
        RECT 4.400 218.600 165.600 218.640 ;
        RECT 4.000 217.960 165.600 218.600 ;
        RECT 4.400 217.240 165.600 217.960 ;
        RECT 4.400 216.600 166.000 217.240 ;
        RECT 4.400 216.560 165.600 216.600 ;
        RECT 4.000 215.920 165.600 216.560 ;
        RECT 4.400 215.200 165.600 215.920 ;
        RECT 4.400 214.560 166.000 215.200 ;
        RECT 4.400 214.520 165.600 214.560 ;
        RECT 4.000 213.880 165.600 214.520 ;
        RECT 4.400 213.160 165.600 213.880 ;
        RECT 4.400 212.520 166.000 213.160 ;
        RECT 4.400 212.480 165.600 212.520 ;
        RECT 4.000 211.840 165.600 212.480 ;
        RECT 4.400 211.120 165.600 211.840 ;
        RECT 4.400 210.480 166.000 211.120 ;
        RECT 4.400 210.440 165.600 210.480 ;
        RECT 4.000 209.800 165.600 210.440 ;
        RECT 4.400 209.080 165.600 209.800 ;
        RECT 4.400 208.440 166.000 209.080 ;
        RECT 4.400 208.400 165.600 208.440 ;
        RECT 4.000 207.760 165.600 208.400 ;
        RECT 4.400 207.040 165.600 207.760 ;
        RECT 4.400 206.400 166.000 207.040 ;
        RECT 4.400 206.360 165.600 206.400 ;
        RECT 4.000 205.720 165.600 206.360 ;
        RECT 4.400 205.000 165.600 205.720 ;
        RECT 4.400 204.360 166.000 205.000 ;
        RECT 4.400 204.320 165.600 204.360 ;
        RECT 4.000 203.680 165.600 204.320 ;
        RECT 4.400 202.960 165.600 203.680 ;
        RECT 4.400 202.320 166.000 202.960 ;
        RECT 4.400 202.280 165.600 202.320 ;
        RECT 4.000 201.640 165.600 202.280 ;
        RECT 4.400 200.920 165.600 201.640 ;
        RECT 4.400 200.280 166.000 200.920 ;
        RECT 4.400 200.240 165.600 200.280 ;
        RECT 4.000 199.600 165.600 200.240 ;
        RECT 4.400 198.880 165.600 199.600 ;
        RECT 4.400 198.240 166.000 198.880 ;
        RECT 4.400 198.200 165.600 198.240 ;
        RECT 4.000 197.560 165.600 198.200 ;
        RECT 4.400 196.840 165.600 197.560 ;
        RECT 4.400 196.200 166.000 196.840 ;
        RECT 4.400 196.160 165.600 196.200 ;
        RECT 4.000 195.520 165.600 196.160 ;
        RECT 4.400 194.800 165.600 195.520 ;
        RECT 4.400 194.160 166.000 194.800 ;
        RECT 4.400 194.120 165.600 194.160 ;
        RECT 4.000 193.480 165.600 194.120 ;
        RECT 4.400 192.760 165.600 193.480 ;
        RECT 4.400 192.120 166.000 192.760 ;
        RECT 4.400 192.080 165.600 192.120 ;
        RECT 4.000 191.440 165.600 192.080 ;
        RECT 4.400 190.720 165.600 191.440 ;
        RECT 4.400 190.080 166.000 190.720 ;
        RECT 4.400 190.040 165.600 190.080 ;
        RECT 4.000 189.400 165.600 190.040 ;
        RECT 4.400 188.680 165.600 189.400 ;
        RECT 4.400 188.040 166.000 188.680 ;
        RECT 4.400 188.000 165.600 188.040 ;
        RECT 4.000 187.360 165.600 188.000 ;
        RECT 4.400 186.640 165.600 187.360 ;
        RECT 4.400 186.000 166.000 186.640 ;
        RECT 4.400 185.960 165.600 186.000 ;
        RECT 4.000 185.320 165.600 185.960 ;
        RECT 4.400 184.600 165.600 185.320 ;
        RECT 4.400 183.960 166.000 184.600 ;
        RECT 4.400 183.920 165.600 183.960 ;
        RECT 4.000 183.280 165.600 183.920 ;
        RECT 4.400 182.560 165.600 183.280 ;
        RECT 4.400 181.920 166.000 182.560 ;
        RECT 4.400 181.880 165.600 181.920 ;
        RECT 4.000 181.240 165.600 181.880 ;
        RECT 4.400 180.520 165.600 181.240 ;
        RECT 4.400 179.880 166.000 180.520 ;
        RECT 4.400 179.840 165.600 179.880 ;
        RECT 4.000 179.200 165.600 179.840 ;
        RECT 4.400 178.480 165.600 179.200 ;
        RECT 4.400 177.840 166.000 178.480 ;
        RECT 4.400 177.800 165.600 177.840 ;
        RECT 4.000 177.160 165.600 177.800 ;
        RECT 4.400 176.440 165.600 177.160 ;
        RECT 4.400 175.800 166.000 176.440 ;
        RECT 4.400 175.760 165.600 175.800 ;
        RECT 4.000 175.120 165.600 175.760 ;
        RECT 4.400 174.400 165.600 175.120 ;
        RECT 4.400 173.760 166.000 174.400 ;
        RECT 4.400 173.720 165.600 173.760 ;
        RECT 4.000 173.080 165.600 173.720 ;
        RECT 4.400 172.360 165.600 173.080 ;
        RECT 4.400 171.720 166.000 172.360 ;
        RECT 4.400 171.680 165.600 171.720 ;
        RECT 4.000 171.040 165.600 171.680 ;
        RECT 4.400 170.320 165.600 171.040 ;
        RECT 4.400 169.680 166.000 170.320 ;
        RECT 4.400 169.640 165.600 169.680 ;
        RECT 4.000 169.000 165.600 169.640 ;
        RECT 4.400 168.280 165.600 169.000 ;
        RECT 4.400 167.640 166.000 168.280 ;
        RECT 4.400 167.600 165.600 167.640 ;
        RECT 4.000 166.960 165.600 167.600 ;
        RECT 4.400 166.240 165.600 166.960 ;
        RECT 4.400 165.600 166.000 166.240 ;
        RECT 4.400 165.560 165.600 165.600 ;
        RECT 4.000 164.920 165.600 165.560 ;
        RECT 4.400 164.200 165.600 164.920 ;
        RECT 4.400 163.560 166.000 164.200 ;
        RECT 4.400 163.520 165.600 163.560 ;
        RECT 4.000 162.880 165.600 163.520 ;
        RECT 4.400 162.160 165.600 162.880 ;
        RECT 4.400 161.520 166.000 162.160 ;
        RECT 4.400 161.480 165.600 161.520 ;
        RECT 4.000 160.840 165.600 161.480 ;
        RECT 4.400 160.120 165.600 160.840 ;
        RECT 4.400 159.480 166.000 160.120 ;
        RECT 4.400 159.440 165.600 159.480 ;
        RECT 4.000 158.800 165.600 159.440 ;
        RECT 4.400 158.080 165.600 158.800 ;
        RECT 4.400 157.440 166.000 158.080 ;
        RECT 4.400 157.400 165.600 157.440 ;
        RECT 4.000 156.760 165.600 157.400 ;
        RECT 4.400 156.040 165.600 156.760 ;
        RECT 4.400 155.400 166.000 156.040 ;
        RECT 4.400 155.360 165.600 155.400 ;
        RECT 4.000 154.720 165.600 155.360 ;
        RECT 4.400 154.000 165.600 154.720 ;
        RECT 4.400 153.360 166.000 154.000 ;
        RECT 4.400 153.320 165.600 153.360 ;
        RECT 4.000 152.680 165.600 153.320 ;
        RECT 4.400 151.960 165.600 152.680 ;
        RECT 4.400 151.320 166.000 151.960 ;
        RECT 4.400 151.280 165.600 151.320 ;
        RECT 4.000 150.640 165.600 151.280 ;
        RECT 4.400 149.920 165.600 150.640 ;
        RECT 4.400 149.280 166.000 149.920 ;
        RECT 4.400 149.240 165.600 149.280 ;
        RECT 4.000 148.600 165.600 149.240 ;
        RECT 4.400 147.880 165.600 148.600 ;
        RECT 4.400 147.240 166.000 147.880 ;
        RECT 4.400 147.200 165.600 147.240 ;
        RECT 4.000 146.560 165.600 147.200 ;
        RECT 4.400 145.840 165.600 146.560 ;
        RECT 4.400 145.200 166.000 145.840 ;
        RECT 4.400 145.160 165.600 145.200 ;
        RECT 4.000 144.520 165.600 145.160 ;
        RECT 4.400 143.800 165.600 144.520 ;
        RECT 4.400 143.160 166.000 143.800 ;
        RECT 4.400 143.120 165.600 143.160 ;
        RECT 4.000 142.480 165.600 143.120 ;
        RECT 4.400 141.080 165.600 142.480 ;
        RECT 4.000 140.440 165.600 141.080 ;
        RECT 4.400 140.400 165.600 140.440 ;
        RECT 4.400 139.760 166.000 140.400 ;
        RECT 4.400 139.040 165.600 139.760 ;
        RECT 4.000 138.400 165.600 139.040 ;
        RECT 4.400 138.360 165.600 138.400 ;
        RECT 4.400 137.720 166.000 138.360 ;
        RECT 4.400 137.000 165.600 137.720 ;
        RECT 4.000 136.360 165.600 137.000 ;
        RECT 4.400 136.320 165.600 136.360 ;
        RECT 4.400 135.680 166.000 136.320 ;
        RECT 4.400 134.960 165.600 135.680 ;
        RECT 4.000 134.320 165.600 134.960 ;
        RECT 4.400 134.280 165.600 134.320 ;
        RECT 4.400 133.640 166.000 134.280 ;
        RECT 4.400 132.920 165.600 133.640 ;
        RECT 4.000 132.280 165.600 132.920 ;
        RECT 4.400 132.240 165.600 132.280 ;
        RECT 4.400 131.600 166.000 132.240 ;
        RECT 4.400 130.880 165.600 131.600 ;
        RECT 4.000 130.240 165.600 130.880 ;
        RECT 4.400 130.200 165.600 130.240 ;
        RECT 4.400 129.560 166.000 130.200 ;
        RECT 4.400 128.840 165.600 129.560 ;
        RECT 4.000 128.200 165.600 128.840 ;
        RECT 4.400 128.160 165.600 128.200 ;
        RECT 4.400 127.520 166.000 128.160 ;
        RECT 4.400 126.800 165.600 127.520 ;
        RECT 4.000 126.160 165.600 126.800 ;
        RECT 4.400 126.120 165.600 126.160 ;
        RECT 4.400 125.480 166.000 126.120 ;
        RECT 4.400 124.760 165.600 125.480 ;
        RECT 4.000 124.120 165.600 124.760 ;
        RECT 4.400 124.080 165.600 124.120 ;
        RECT 4.400 123.440 166.000 124.080 ;
        RECT 4.400 122.720 165.600 123.440 ;
        RECT 4.000 122.080 165.600 122.720 ;
        RECT 4.400 122.040 165.600 122.080 ;
        RECT 4.400 121.400 166.000 122.040 ;
        RECT 4.400 120.680 165.600 121.400 ;
        RECT 4.000 120.040 165.600 120.680 ;
        RECT 4.400 120.000 165.600 120.040 ;
        RECT 4.400 119.360 166.000 120.000 ;
        RECT 4.400 118.640 165.600 119.360 ;
        RECT 4.000 118.000 165.600 118.640 ;
        RECT 4.400 117.960 165.600 118.000 ;
        RECT 4.400 117.320 166.000 117.960 ;
        RECT 4.400 116.600 165.600 117.320 ;
        RECT 4.000 115.960 165.600 116.600 ;
        RECT 4.400 115.920 165.600 115.960 ;
        RECT 4.400 115.280 166.000 115.920 ;
        RECT 4.400 114.560 165.600 115.280 ;
        RECT 4.000 113.920 165.600 114.560 ;
        RECT 4.400 113.880 165.600 113.920 ;
        RECT 4.400 113.240 166.000 113.880 ;
        RECT 4.400 112.520 165.600 113.240 ;
        RECT 4.000 111.880 165.600 112.520 ;
        RECT 4.400 111.840 165.600 111.880 ;
        RECT 4.400 111.200 166.000 111.840 ;
        RECT 4.400 110.480 165.600 111.200 ;
        RECT 4.000 109.840 165.600 110.480 ;
        RECT 4.400 109.800 165.600 109.840 ;
        RECT 4.400 109.160 166.000 109.800 ;
        RECT 4.400 108.440 165.600 109.160 ;
        RECT 4.000 107.800 165.600 108.440 ;
        RECT 4.400 107.760 165.600 107.800 ;
        RECT 4.400 107.120 166.000 107.760 ;
        RECT 4.400 106.400 165.600 107.120 ;
        RECT 4.000 105.760 165.600 106.400 ;
        RECT 4.400 105.720 165.600 105.760 ;
        RECT 4.400 105.080 166.000 105.720 ;
        RECT 4.400 104.360 165.600 105.080 ;
        RECT 4.000 103.720 165.600 104.360 ;
        RECT 4.400 103.680 165.600 103.720 ;
        RECT 4.400 103.040 166.000 103.680 ;
        RECT 4.400 102.320 165.600 103.040 ;
        RECT 4.000 101.680 165.600 102.320 ;
        RECT 4.400 101.640 165.600 101.680 ;
        RECT 4.400 101.000 166.000 101.640 ;
        RECT 4.400 100.280 165.600 101.000 ;
        RECT 4.000 99.640 165.600 100.280 ;
        RECT 4.400 99.600 165.600 99.640 ;
        RECT 4.400 98.960 166.000 99.600 ;
        RECT 4.400 98.240 165.600 98.960 ;
        RECT 4.000 97.600 165.600 98.240 ;
        RECT 4.400 97.560 165.600 97.600 ;
        RECT 4.400 96.920 166.000 97.560 ;
        RECT 4.400 96.200 165.600 96.920 ;
        RECT 4.000 95.560 165.600 96.200 ;
        RECT 4.400 95.520 165.600 95.560 ;
        RECT 4.400 94.880 166.000 95.520 ;
        RECT 4.400 94.160 165.600 94.880 ;
        RECT 4.000 93.520 165.600 94.160 ;
        RECT 4.400 93.480 165.600 93.520 ;
        RECT 4.400 92.840 166.000 93.480 ;
        RECT 4.400 92.120 165.600 92.840 ;
        RECT 4.000 91.480 165.600 92.120 ;
        RECT 4.400 91.440 165.600 91.480 ;
        RECT 4.400 90.800 166.000 91.440 ;
        RECT 4.400 90.080 165.600 90.800 ;
        RECT 4.000 89.440 165.600 90.080 ;
        RECT 4.400 89.400 165.600 89.440 ;
        RECT 4.400 88.760 166.000 89.400 ;
        RECT 4.400 88.040 165.600 88.760 ;
        RECT 4.000 87.400 165.600 88.040 ;
        RECT 4.400 87.360 165.600 87.400 ;
        RECT 4.400 86.720 166.000 87.360 ;
        RECT 4.400 86.000 165.600 86.720 ;
        RECT 4.000 85.360 165.600 86.000 ;
        RECT 4.400 85.320 165.600 85.360 ;
        RECT 4.400 84.680 166.000 85.320 ;
        RECT 4.400 83.960 165.600 84.680 ;
        RECT 4.000 83.320 165.600 83.960 ;
        RECT 4.400 83.280 165.600 83.320 ;
        RECT 4.400 82.640 166.000 83.280 ;
        RECT 4.400 81.920 165.600 82.640 ;
        RECT 4.000 81.280 165.600 81.920 ;
        RECT 4.400 81.240 165.600 81.280 ;
        RECT 4.400 80.600 166.000 81.240 ;
        RECT 4.400 79.880 165.600 80.600 ;
        RECT 4.000 79.240 165.600 79.880 ;
        RECT 4.400 79.200 165.600 79.240 ;
        RECT 4.400 78.560 166.000 79.200 ;
        RECT 4.400 77.840 165.600 78.560 ;
        RECT 4.000 77.200 165.600 77.840 ;
        RECT 4.400 77.160 165.600 77.200 ;
        RECT 4.400 76.520 166.000 77.160 ;
        RECT 4.400 75.800 165.600 76.520 ;
        RECT 4.000 75.160 165.600 75.800 ;
        RECT 4.400 75.120 165.600 75.160 ;
        RECT 4.400 74.480 166.000 75.120 ;
        RECT 4.400 73.760 165.600 74.480 ;
        RECT 4.000 73.120 165.600 73.760 ;
        RECT 4.400 73.080 165.600 73.120 ;
        RECT 4.400 72.440 166.000 73.080 ;
        RECT 4.400 71.720 165.600 72.440 ;
        RECT 4.000 71.080 165.600 71.720 ;
        RECT 4.400 71.040 165.600 71.080 ;
        RECT 4.400 70.400 166.000 71.040 ;
        RECT 4.400 69.680 165.600 70.400 ;
        RECT 4.000 69.040 165.600 69.680 ;
        RECT 4.400 69.000 165.600 69.040 ;
        RECT 4.400 68.360 166.000 69.000 ;
        RECT 4.400 67.640 165.600 68.360 ;
        RECT 4.000 67.000 165.600 67.640 ;
        RECT 4.400 66.960 165.600 67.000 ;
        RECT 4.400 66.320 166.000 66.960 ;
        RECT 4.400 65.600 165.600 66.320 ;
        RECT 4.000 64.960 165.600 65.600 ;
        RECT 4.400 64.920 165.600 64.960 ;
        RECT 4.400 64.280 166.000 64.920 ;
        RECT 4.400 63.560 165.600 64.280 ;
        RECT 4.000 62.920 165.600 63.560 ;
        RECT 4.400 62.880 165.600 62.920 ;
        RECT 4.400 62.240 166.000 62.880 ;
        RECT 4.400 61.520 165.600 62.240 ;
        RECT 4.000 60.880 165.600 61.520 ;
        RECT 4.400 60.840 165.600 60.880 ;
        RECT 4.400 60.200 166.000 60.840 ;
        RECT 4.400 59.480 165.600 60.200 ;
        RECT 4.000 58.840 165.600 59.480 ;
        RECT 4.400 58.800 165.600 58.840 ;
        RECT 4.400 58.160 166.000 58.800 ;
        RECT 4.400 57.440 165.600 58.160 ;
        RECT 4.000 56.800 165.600 57.440 ;
        RECT 4.400 56.760 165.600 56.800 ;
        RECT 4.400 56.120 166.000 56.760 ;
        RECT 4.400 55.400 165.600 56.120 ;
        RECT 4.000 54.760 165.600 55.400 ;
        RECT 4.400 54.720 165.600 54.760 ;
        RECT 4.400 54.080 166.000 54.720 ;
        RECT 4.400 53.360 165.600 54.080 ;
        RECT 4.000 52.720 165.600 53.360 ;
        RECT 4.400 52.680 165.600 52.720 ;
        RECT 4.400 52.040 166.000 52.680 ;
        RECT 4.400 51.320 165.600 52.040 ;
        RECT 4.000 50.680 165.600 51.320 ;
        RECT 4.400 50.640 165.600 50.680 ;
        RECT 4.400 50.000 166.000 50.640 ;
        RECT 4.400 49.280 165.600 50.000 ;
        RECT 4.000 48.640 165.600 49.280 ;
        RECT 4.400 48.600 165.600 48.640 ;
        RECT 4.400 47.960 166.000 48.600 ;
        RECT 4.400 47.240 165.600 47.960 ;
        RECT 4.000 46.600 165.600 47.240 ;
        RECT 4.400 46.560 165.600 46.600 ;
        RECT 4.400 45.920 166.000 46.560 ;
        RECT 4.400 45.200 165.600 45.920 ;
        RECT 4.000 44.560 165.600 45.200 ;
        RECT 4.400 44.520 165.600 44.560 ;
        RECT 4.400 43.880 166.000 44.520 ;
        RECT 4.400 43.160 165.600 43.880 ;
        RECT 4.000 42.520 165.600 43.160 ;
        RECT 4.400 42.480 165.600 42.520 ;
        RECT 4.400 41.840 166.000 42.480 ;
        RECT 4.400 41.120 165.600 41.840 ;
        RECT 4.000 40.480 165.600 41.120 ;
        RECT 4.400 40.440 165.600 40.480 ;
        RECT 4.400 39.800 166.000 40.440 ;
        RECT 4.400 39.080 165.600 39.800 ;
        RECT 4.000 38.440 165.600 39.080 ;
        RECT 4.400 38.400 165.600 38.440 ;
        RECT 4.400 37.760 166.000 38.400 ;
        RECT 4.400 37.040 165.600 37.760 ;
        RECT 4.000 36.400 165.600 37.040 ;
        RECT 4.400 36.360 165.600 36.400 ;
        RECT 4.400 35.720 166.000 36.360 ;
        RECT 4.400 35.000 165.600 35.720 ;
        RECT 4.000 34.360 165.600 35.000 ;
        RECT 4.400 34.320 165.600 34.360 ;
        RECT 4.400 33.680 166.000 34.320 ;
        RECT 4.400 32.960 165.600 33.680 ;
        RECT 4.000 32.320 165.600 32.960 ;
        RECT 4.400 32.280 165.600 32.320 ;
        RECT 4.400 31.640 166.000 32.280 ;
        RECT 4.400 30.920 165.600 31.640 ;
        RECT 4.000 30.280 165.600 30.920 ;
        RECT 4.400 30.240 165.600 30.280 ;
        RECT 4.400 29.600 166.000 30.240 ;
        RECT 4.400 28.880 165.600 29.600 ;
        RECT 4.000 28.240 165.600 28.880 ;
        RECT 4.400 28.200 165.600 28.240 ;
        RECT 4.400 27.560 166.000 28.200 ;
        RECT 4.400 26.840 165.600 27.560 ;
        RECT 4.000 26.200 165.600 26.840 ;
        RECT 4.400 26.160 165.600 26.200 ;
        RECT 4.400 25.520 166.000 26.160 ;
        RECT 4.400 24.800 165.600 25.520 ;
        RECT 4.000 24.160 165.600 24.800 ;
        RECT 4.400 24.120 165.600 24.160 ;
        RECT 4.400 23.480 166.000 24.120 ;
        RECT 4.400 22.760 165.600 23.480 ;
        RECT 4.000 22.120 165.600 22.760 ;
        RECT 4.400 22.080 165.600 22.120 ;
        RECT 4.400 21.440 166.000 22.080 ;
        RECT 4.400 20.720 165.600 21.440 ;
        RECT 4.000 20.080 165.600 20.720 ;
        RECT 4.400 20.040 165.600 20.080 ;
        RECT 4.400 19.400 166.000 20.040 ;
        RECT 4.400 18.680 165.600 19.400 ;
        RECT 4.000 18.040 165.600 18.680 ;
        RECT 4.400 18.000 165.600 18.040 ;
        RECT 4.400 17.360 166.000 18.000 ;
        RECT 4.400 16.640 165.600 17.360 ;
        RECT 4.000 16.000 165.600 16.640 ;
        RECT 4.400 15.960 165.600 16.000 ;
        RECT 4.400 15.320 166.000 15.960 ;
        RECT 4.400 14.600 165.600 15.320 ;
        RECT 4.000 13.960 165.600 14.600 ;
        RECT 4.400 13.920 165.600 13.960 ;
        RECT 4.400 13.280 166.000 13.920 ;
        RECT 4.400 12.560 165.600 13.280 ;
        RECT 4.000 11.920 165.600 12.560 ;
        RECT 4.400 11.880 165.600 11.920 ;
        RECT 4.400 11.240 166.000 11.880 ;
        RECT 4.400 10.520 165.600 11.240 ;
        RECT 4.000 9.880 165.600 10.520 ;
        RECT 4.400 9.840 165.600 9.880 ;
        RECT 4.400 9.200 166.000 9.840 ;
        RECT 4.400 8.480 165.600 9.200 ;
        RECT 4.000 7.840 165.600 8.480 ;
        RECT 4.400 7.800 165.600 7.840 ;
        RECT 4.400 7.160 166.000 7.800 ;
        RECT 4.400 6.440 165.600 7.160 ;
        RECT 4.000 5.800 165.600 6.440 ;
        RECT 4.400 5.760 165.600 5.800 ;
        RECT 4.400 5.120 166.000 5.760 ;
        RECT 4.400 4.400 165.600 5.120 ;
        RECT 4.000 3.760 165.600 4.400 ;
        RECT 4.400 3.720 165.600 3.760 ;
        RECT 4.400 3.080 166.000 3.720 ;
        RECT 4.400 2.360 165.600 3.080 ;
        RECT 4.000 1.720 165.600 2.360 ;
        RECT 4.400 0.855 165.600 1.720 ;
      LAYER met4 ;
        RECT 33.215 10.640 57.305 266.800 ;
        RECT 59.705 10.640 83.800 266.800 ;
        RECT 86.200 10.640 110.295 266.800 ;
  END
END cic_block
END LIBRARY

