magic
tech sky130A
magscale 1 2
timestamp 1624040213
<< obsli1 >>
rect 1104 1649 32999 53329
<< obsm1 >>
rect 750 1300 33290 54732
<< metal2 >>
rect 1030 55200 1086 56800
rect 3146 55200 3202 56800
rect 5262 55200 5318 56800
rect 7378 55200 7434 56800
rect 9494 55200 9550 56800
rect 11610 55200 11666 56800
rect 13726 55200 13782 56800
rect 15842 55200 15898 56800
rect 18050 55200 18106 56800
rect 20166 55200 20222 56800
rect 22282 55200 22338 56800
rect 24398 55200 24454 56800
rect 26514 55200 26570 56800
rect 28630 55200 28686 56800
rect 30746 55200 30802 56800
rect 32862 55200 32918 56800
rect 754 -800 810 800
rect 2226 -800 2282 800
rect 3790 -800 3846 800
rect 5354 -800 5410 800
rect 6918 -800 6974 800
rect 8482 -800 8538 800
rect 9954 -800 10010 800
rect 11518 -800 11574 800
rect 13082 -800 13138 800
rect 14646 -800 14702 800
rect 16210 -800 16266 800
rect 17774 -800 17830 800
rect 19246 -800 19302 800
rect 20810 -800 20866 800
rect 22374 -800 22430 800
rect 23938 -800 23994 800
rect 25502 -800 25558 800
rect 26974 -800 27030 800
rect 28538 -800 28594 800
rect 30102 -800 30158 800
rect 31666 -800 31722 800
rect 33230 -800 33286 800
<< obsm2 >>
rect 756 55144 974 55865
rect 1142 55144 3090 55865
rect 3258 55144 5206 55865
rect 5374 55144 7322 55865
rect 7490 55144 9438 55865
rect 9606 55144 11554 55865
rect 11722 55144 13670 55865
rect 13838 55144 15786 55865
rect 15954 55144 17994 55865
rect 18162 55144 20110 55865
rect 20278 55144 22226 55865
rect 22394 55144 24342 55865
rect 24510 55144 26458 55865
rect 26626 55144 28574 55865
rect 28742 55144 30690 55865
rect 30858 55144 32806 55865
rect 32974 55144 33284 55865
rect 756 856 33284 55144
rect 866 167 2170 856
rect 2338 167 3734 856
rect 3902 167 5298 856
rect 5466 167 6862 856
rect 7030 167 8426 856
rect 8594 167 9898 856
rect 10066 167 11462 856
rect 11630 167 13026 856
rect 13194 167 14590 856
rect 14758 167 16154 856
rect 16322 167 17718 856
rect 17886 167 19190 856
rect 19358 167 20754 856
rect 20922 167 22318 856
rect 22486 167 23882 856
rect 24050 167 25446 856
rect 25614 167 26918 856
rect 27086 167 28482 856
rect 28650 167 30046 856
rect 30214 167 31610 856
rect 31778 167 33174 856
<< metal3 >>
rect -800 55632 800 55752
rect 33200 55768 34800 55888
rect -800 55224 800 55344
rect 33200 55360 34800 55480
rect -800 54816 800 54936
rect 33200 54952 34800 55072
rect -800 54408 800 54528
rect 33200 54544 34800 54664
rect -800 54000 800 54120
rect 33200 54136 34800 54256
rect -800 53592 800 53712
rect 33200 53728 34800 53848
rect -800 53184 800 53304
rect 33200 53320 34800 53440
rect -800 52776 800 52896
rect 33200 52912 34800 53032
rect -800 52368 800 52488
rect 33200 52504 34800 52624
rect -800 51960 800 52080
rect 33200 52096 34800 52216
rect -800 51552 800 51672
rect 33200 51688 34800 51808
rect -800 51144 800 51264
rect 33200 51280 34800 51400
rect -800 50736 800 50856
rect 33200 50872 34800 50992
rect -800 50328 800 50448
rect 33200 50464 34800 50584
rect -800 49920 800 50040
rect 33200 50056 34800 50176
rect -800 49512 800 49632
rect 33200 49648 34800 49768
rect -800 49104 800 49224
rect 33200 49240 34800 49360
rect -800 48696 800 48816
rect 33200 48832 34800 48952
rect -800 48288 800 48408
rect 33200 48424 34800 48544
rect -800 47880 800 48000
rect 33200 48016 34800 48136
rect -800 47472 800 47592
rect 33200 47608 34800 47728
rect -800 47064 800 47184
rect 33200 47200 34800 47320
rect -800 46656 800 46776
rect 33200 46792 34800 46912
rect -800 46248 800 46368
rect 33200 46384 34800 46504
rect -800 45840 800 45960
rect 33200 45976 34800 46096
rect -800 45432 800 45552
rect 33200 45568 34800 45688
rect -800 45024 800 45144
rect 33200 45160 34800 45280
rect -800 44616 800 44736
rect 33200 44752 34800 44872
rect -800 44208 800 44328
rect 33200 44344 34800 44464
rect -800 43800 800 43920
rect 33200 43936 34800 44056
rect -800 43392 800 43512
rect 33200 43528 34800 43648
rect -800 42984 800 43104
rect 33200 43120 34800 43240
rect -800 42576 800 42696
rect 33200 42712 34800 42832
rect -800 42168 800 42288
rect 33200 42304 34800 42424
rect -800 41760 800 41880
rect 33200 41896 34800 42016
rect -800 41352 800 41472
rect 33200 41488 34800 41608
rect -800 40944 800 41064
rect 33200 41080 34800 41200
rect -800 40536 800 40656
rect 33200 40672 34800 40792
rect -800 40128 800 40248
rect 33200 40264 34800 40384
rect -800 39720 800 39840
rect 33200 39856 34800 39976
rect -800 39312 800 39432
rect 33200 39448 34800 39568
rect -800 38904 800 39024
rect 33200 39040 34800 39160
rect -800 38496 800 38616
rect 33200 38632 34800 38752
rect -800 38088 800 38208
rect 33200 38224 34800 38344
rect -800 37680 800 37800
rect 33200 37816 34800 37936
rect -800 37272 800 37392
rect 33200 37408 34800 37528
rect -800 36864 800 36984
rect 33200 37000 34800 37120
rect -800 36456 800 36576
rect 33200 36592 34800 36712
rect -800 36048 800 36168
rect 33200 36184 34800 36304
rect -800 35640 800 35760
rect 33200 35776 34800 35896
rect -800 35232 800 35352
rect 33200 35368 34800 35488
rect -800 34824 800 34944
rect 33200 34960 34800 35080
rect -800 34416 800 34536
rect 33200 34552 34800 34672
rect -800 34008 800 34128
rect 33200 34144 34800 34264
rect -800 33600 800 33720
rect 33200 33736 34800 33856
rect -800 33192 800 33312
rect 33200 33328 34800 33448
rect -800 32784 800 32904
rect 33200 32920 34800 33040
rect -800 32376 800 32496
rect 33200 32512 34800 32632
rect -800 31968 800 32088
rect 33200 32104 34800 32224
rect -800 31560 800 31680
rect 33200 31696 34800 31816
rect -800 31152 800 31272
rect 33200 31288 34800 31408
rect -800 30744 800 30864
rect 33200 30880 34800 31000
rect -800 30336 800 30456
rect 33200 30472 34800 30592
rect -800 29928 800 30048
rect 33200 30064 34800 30184
rect -800 29520 800 29640
rect 33200 29656 34800 29776
rect -800 29112 800 29232
rect 33200 29248 34800 29368
rect -800 28704 800 28824
rect 33200 28840 34800 28960
rect -800 28296 800 28416
rect 33200 28432 34800 28552
rect 33200 28160 34800 28280
rect -800 27888 800 28008
rect 33200 27752 34800 27872
rect -800 27480 800 27600
rect 33200 27344 34800 27464
rect -800 27072 800 27192
rect 33200 26936 34800 27056
rect -800 26664 800 26784
rect 33200 26528 34800 26648
rect -800 26256 800 26376
rect 33200 26120 34800 26240
rect -800 25848 800 25968
rect 33200 25712 34800 25832
rect -800 25440 800 25560
rect 33200 25304 34800 25424
rect -800 25032 800 25152
rect 33200 24896 34800 25016
rect -800 24624 800 24744
rect 33200 24488 34800 24608
rect -800 24216 800 24336
rect 33200 24080 34800 24200
rect -800 23808 800 23928
rect 33200 23672 34800 23792
rect -800 23400 800 23520
rect 33200 23264 34800 23384
rect -800 22992 800 23112
rect 33200 22856 34800 22976
rect -800 22584 800 22704
rect 33200 22448 34800 22568
rect -800 22176 800 22296
rect 33200 22040 34800 22160
rect -800 21768 800 21888
rect 33200 21632 34800 21752
rect -800 21360 800 21480
rect 33200 21224 34800 21344
rect -800 20952 800 21072
rect 33200 20816 34800 20936
rect -800 20544 800 20664
rect 33200 20408 34800 20528
rect -800 20136 800 20256
rect 33200 20000 34800 20120
rect -800 19728 800 19848
rect 33200 19592 34800 19712
rect -800 19320 800 19440
rect 33200 19184 34800 19304
rect -800 18912 800 19032
rect 33200 18776 34800 18896
rect -800 18504 800 18624
rect 33200 18368 34800 18488
rect -800 18096 800 18216
rect 33200 17960 34800 18080
rect -800 17688 800 17808
rect 33200 17552 34800 17672
rect -800 17280 800 17400
rect 33200 17144 34800 17264
rect -800 16872 800 16992
rect 33200 16736 34800 16856
rect -800 16464 800 16584
rect 33200 16328 34800 16448
rect -800 16056 800 16176
rect 33200 15920 34800 16040
rect -800 15648 800 15768
rect 33200 15512 34800 15632
rect -800 15240 800 15360
rect 33200 15104 34800 15224
rect -800 14832 800 14952
rect 33200 14696 34800 14816
rect -800 14424 800 14544
rect 33200 14288 34800 14408
rect -800 14016 800 14136
rect 33200 13880 34800 14000
rect -800 13608 800 13728
rect 33200 13472 34800 13592
rect -800 13200 800 13320
rect 33200 13064 34800 13184
rect -800 12792 800 12912
rect 33200 12656 34800 12776
rect -800 12384 800 12504
rect 33200 12248 34800 12368
rect -800 11976 800 12096
rect 33200 11840 34800 11960
rect -800 11568 800 11688
rect 33200 11432 34800 11552
rect -800 11160 800 11280
rect 33200 11024 34800 11144
rect -800 10752 800 10872
rect 33200 10616 34800 10736
rect -800 10344 800 10464
rect 33200 10208 34800 10328
rect -800 9936 800 10056
rect 33200 9800 34800 9920
rect -800 9528 800 9648
rect 33200 9392 34800 9512
rect -800 9120 800 9240
rect 33200 8984 34800 9104
rect -800 8712 800 8832
rect 33200 8576 34800 8696
rect -800 8304 800 8424
rect 33200 8168 34800 8288
rect -800 7896 800 8016
rect 33200 7760 34800 7880
rect -800 7488 800 7608
rect 33200 7352 34800 7472
rect -800 7080 800 7200
rect 33200 6944 34800 7064
rect -800 6672 800 6792
rect 33200 6536 34800 6656
rect -800 6264 800 6384
rect 33200 6128 34800 6248
rect -800 5856 800 5976
rect 33200 5720 34800 5840
rect -800 5448 800 5568
rect 33200 5312 34800 5432
rect -800 5040 800 5160
rect 33200 4904 34800 5024
rect -800 4632 800 4752
rect 33200 4496 34800 4616
rect -800 4224 800 4344
rect 33200 4088 34800 4208
rect -800 3816 800 3936
rect 33200 3680 34800 3800
rect -800 3408 800 3528
rect 33200 3272 34800 3392
rect -800 3000 800 3120
rect 33200 2864 34800 2984
rect -800 2592 800 2712
rect 33200 2456 34800 2576
rect -800 2184 800 2304
rect 33200 2048 34800 2168
rect -800 1776 800 1896
rect 33200 1640 34800 1760
rect -800 1368 800 1488
rect 33200 1232 34800 1352
rect -800 960 800 1080
rect 33200 824 34800 944
rect -800 552 800 672
rect 33200 416 34800 536
rect -800 144 800 264
rect 33200 144 34800 264
<< obsm3 >>
rect 800 55832 33120 55861
rect 880 55688 33120 55832
rect 880 55560 33200 55688
rect 880 55552 33120 55560
rect 800 55424 33120 55552
rect 880 55280 33120 55424
rect 880 55152 33200 55280
rect 880 55144 33120 55152
rect 800 55016 33120 55144
rect 880 54872 33120 55016
rect 880 54744 33200 54872
rect 880 54736 33120 54744
rect 800 54608 33120 54736
rect 880 54464 33120 54608
rect 880 54336 33200 54464
rect 880 54328 33120 54336
rect 800 54200 33120 54328
rect 880 54056 33120 54200
rect 880 53928 33200 54056
rect 880 53920 33120 53928
rect 800 53792 33120 53920
rect 880 53648 33120 53792
rect 880 53520 33200 53648
rect 880 53512 33120 53520
rect 800 53384 33120 53512
rect 880 53240 33120 53384
rect 880 53112 33200 53240
rect 880 53104 33120 53112
rect 800 52976 33120 53104
rect 880 52832 33120 52976
rect 880 52704 33200 52832
rect 880 52696 33120 52704
rect 800 52568 33120 52696
rect 880 52424 33120 52568
rect 880 52296 33200 52424
rect 880 52288 33120 52296
rect 800 52160 33120 52288
rect 880 52016 33120 52160
rect 880 51888 33200 52016
rect 880 51880 33120 51888
rect 800 51752 33120 51880
rect 880 51608 33120 51752
rect 880 51480 33200 51608
rect 880 51472 33120 51480
rect 800 51344 33120 51472
rect 880 51200 33120 51344
rect 880 51072 33200 51200
rect 880 51064 33120 51072
rect 800 50936 33120 51064
rect 880 50792 33120 50936
rect 880 50664 33200 50792
rect 880 50656 33120 50664
rect 800 50528 33120 50656
rect 880 50384 33120 50528
rect 880 50256 33200 50384
rect 880 50248 33120 50256
rect 800 50120 33120 50248
rect 880 49976 33120 50120
rect 880 49848 33200 49976
rect 880 49840 33120 49848
rect 800 49712 33120 49840
rect 880 49568 33120 49712
rect 880 49440 33200 49568
rect 880 49432 33120 49440
rect 800 49304 33120 49432
rect 880 49160 33120 49304
rect 880 49032 33200 49160
rect 880 49024 33120 49032
rect 800 48896 33120 49024
rect 880 48752 33120 48896
rect 880 48624 33200 48752
rect 880 48616 33120 48624
rect 800 48488 33120 48616
rect 880 48344 33120 48488
rect 880 48216 33200 48344
rect 880 48208 33120 48216
rect 800 48080 33120 48208
rect 880 47936 33120 48080
rect 880 47808 33200 47936
rect 880 47800 33120 47808
rect 800 47672 33120 47800
rect 880 47528 33120 47672
rect 880 47400 33200 47528
rect 880 47392 33120 47400
rect 800 47264 33120 47392
rect 880 47120 33120 47264
rect 880 46992 33200 47120
rect 880 46984 33120 46992
rect 800 46856 33120 46984
rect 880 46712 33120 46856
rect 880 46584 33200 46712
rect 880 46576 33120 46584
rect 800 46448 33120 46576
rect 880 46304 33120 46448
rect 880 46176 33200 46304
rect 880 46168 33120 46176
rect 800 46040 33120 46168
rect 880 45896 33120 46040
rect 880 45768 33200 45896
rect 880 45760 33120 45768
rect 800 45632 33120 45760
rect 880 45488 33120 45632
rect 880 45360 33200 45488
rect 880 45352 33120 45360
rect 800 45224 33120 45352
rect 880 45080 33120 45224
rect 880 44952 33200 45080
rect 880 44944 33120 44952
rect 800 44816 33120 44944
rect 880 44672 33120 44816
rect 880 44544 33200 44672
rect 880 44536 33120 44544
rect 800 44408 33120 44536
rect 880 44264 33120 44408
rect 880 44136 33200 44264
rect 880 44128 33120 44136
rect 800 44000 33120 44128
rect 880 43856 33120 44000
rect 880 43728 33200 43856
rect 880 43720 33120 43728
rect 800 43592 33120 43720
rect 880 43448 33120 43592
rect 880 43320 33200 43448
rect 880 43312 33120 43320
rect 800 43184 33120 43312
rect 880 43040 33120 43184
rect 880 42912 33200 43040
rect 880 42904 33120 42912
rect 800 42776 33120 42904
rect 880 42632 33120 42776
rect 880 42504 33200 42632
rect 880 42496 33120 42504
rect 800 42368 33120 42496
rect 880 42224 33120 42368
rect 880 42096 33200 42224
rect 880 42088 33120 42096
rect 800 41960 33120 42088
rect 880 41816 33120 41960
rect 880 41688 33200 41816
rect 880 41680 33120 41688
rect 800 41552 33120 41680
rect 880 41408 33120 41552
rect 880 41280 33200 41408
rect 880 41272 33120 41280
rect 800 41144 33120 41272
rect 880 41000 33120 41144
rect 880 40872 33200 41000
rect 880 40864 33120 40872
rect 800 40736 33120 40864
rect 880 40592 33120 40736
rect 880 40464 33200 40592
rect 880 40456 33120 40464
rect 800 40328 33120 40456
rect 880 40184 33120 40328
rect 880 40056 33200 40184
rect 880 40048 33120 40056
rect 800 39920 33120 40048
rect 880 39776 33120 39920
rect 880 39648 33200 39776
rect 880 39640 33120 39648
rect 800 39512 33120 39640
rect 880 39368 33120 39512
rect 880 39240 33200 39368
rect 880 39232 33120 39240
rect 800 39104 33120 39232
rect 880 38960 33120 39104
rect 880 38832 33200 38960
rect 880 38824 33120 38832
rect 800 38696 33120 38824
rect 880 38552 33120 38696
rect 880 38424 33200 38552
rect 880 38416 33120 38424
rect 800 38288 33120 38416
rect 880 38144 33120 38288
rect 880 38016 33200 38144
rect 880 38008 33120 38016
rect 800 37880 33120 38008
rect 880 37736 33120 37880
rect 880 37608 33200 37736
rect 880 37600 33120 37608
rect 800 37472 33120 37600
rect 880 37328 33120 37472
rect 880 37200 33200 37328
rect 880 37192 33120 37200
rect 800 37064 33120 37192
rect 880 36920 33120 37064
rect 880 36792 33200 36920
rect 880 36784 33120 36792
rect 800 36656 33120 36784
rect 880 36512 33120 36656
rect 880 36384 33200 36512
rect 880 36376 33120 36384
rect 800 36248 33120 36376
rect 880 36104 33120 36248
rect 880 35976 33200 36104
rect 880 35968 33120 35976
rect 800 35840 33120 35968
rect 880 35696 33120 35840
rect 880 35568 33200 35696
rect 880 35560 33120 35568
rect 800 35432 33120 35560
rect 880 35288 33120 35432
rect 880 35160 33200 35288
rect 880 35152 33120 35160
rect 800 35024 33120 35152
rect 880 34880 33120 35024
rect 880 34752 33200 34880
rect 880 34744 33120 34752
rect 800 34616 33120 34744
rect 880 34472 33120 34616
rect 880 34344 33200 34472
rect 880 34336 33120 34344
rect 800 34208 33120 34336
rect 880 34064 33120 34208
rect 880 33936 33200 34064
rect 880 33928 33120 33936
rect 800 33800 33120 33928
rect 880 33656 33120 33800
rect 880 33528 33200 33656
rect 880 33520 33120 33528
rect 800 33392 33120 33520
rect 880 33248 33120 33392
rect 880 33120 33200 33248
rect 880 33112 33120 33120
rect 800 32984 33120 33112
rect 880 32840 33120 32984
rect 880 32712 33200 32840
rect 880 32704 33120 32712
rect 800 32576 33120 32704
rect 880 32432 33120 32576
rect 880 32304 33200 32432
rect 880 32296 33120 32304
rect 800 32168 33120 32296
rect 880 32024 33120 32168
rect 880 31896 33200 32024
rect 880 31888 33120 31896
rect 800 31760 33120 31888
rect 880 31616 33120 31760
rect 880 31488 33200 31616
rect 880 31480 33120 31488
rect 800 31352 33120 31480
rect 880 31208 33120 31352
rect 880 31080 33200 31208
rect 880 31072 33120 31080
rect 800 30944 33120 31072
rect 880 30800 33120 30944
rect 880 30672 33200 30800
rect 880 30664 33120 30672
rect 800 30536 33120 30664
rect 880 30392 33120 30536
rect 880 30264 33200 30392
rect 880 30256 33120 30264
rect 800 30128 33120 30256
rect 880 29984 33120 30128
rect 880 29856 33200 29984
rect 880 29848 33120 29856
rect 800 29720 33120 29848
rect 880 29576 33120 29720
rect 880 29448 33200 29576
rect 880 29440 33120 29448
rect 800 29312 33120 29440
rect 880 29168 33120 29312
rect 880 29040 33200 29168
rect 880 29032 33120 29040
rect 800 28904 33120 29032
rect 880 28760 33120 28904
rect 880 28632 33200 28760
rect 880 28624 33120 28632
rect 800 28496 33120 28624
rect 880 28216 33120 28496
rect 800 28088 33120 28216
rect 880 28080 33120 28088
rect 880 27952 33200 28080
rect 880 27808 33120 27952
rect 800 27680 33120 27808
rect 880 27672 33120 27680
rect 880 27544 33200 27672
rect 880 27400 33120 27544
rect 800 27272 33120 27400
rect 880 27264 33120 27272
rect 880 27136 33200 27264
rect 880 26992 33120 27136
rect 800 26864 33120 26992
rect 880 26856 33120 26864
rect 880 26728 33200 26856
rect 880 26584 33120 26728
rect 800 26456 33120 26584
rect 880 26448 33120 26456
rect 880 26320 33200 26448
rect 880 26176 33120 26320
rect 800 26048 33120 26176
rect 880 26040 33120 26048
rect 880 25912 33200 26040
rect 880 25768 33120 25912
rect 800 25640 33120 25768
rect 880 25632 33120 25640
rect 880 25504 33200 25632
rect 880 25360 33120 25504
rect 800 25232 33120 25360
rect 880 25224 33120 25232
rect 880 25096 33200 25224
rect 880 24952 33120 25096
rect 800 24824 33120 24952
rect 880 24816 33120 24824
rect 880 24688 33200 24816
rect 880 24544 33120 24688
rect 800 24416 33120 24544
rect 880 24408 33120 24416
rect 880 24280 33200 24408
rect 880 24136 33120 24280
rect 800 24008 33120 24136
rect 880 24000 33120 24008
rect 880 23872 33200 24000
rect 880 23728 33120 23872
rect 800 23600 33120 23728
rect 880 23592 33120 23600
rect 880 23464 33200 23592
rect 880 23320 33120 23464
rect 800 23192 33120 23320
rect 880 23184 33120 23192
rect 880 23056 33200 23184
rect 880 22912 33120 23056
rect 800 22784 33120 22912
rect 880 22776 33120 22784
rect 880 22648 33200 22776
rect 880 22504 33120 22648
rect 800 22376 33120 22504
rect 880 22368 33120 22376
rect 880 22240 33200 22368
rect 880 22096 33120 22240
rect 800 21968 33120 22096
rect 880 21960 33120 21968
rect 880 21832 33200 21960
rect 880 21688 33120 21832
rect 800 21560 33120 21688
rect 880 21552 33120 21560
rect 880 21424 33200 21552
rect 880 21280 33120 21424
rect 800 21152 33120 21280
rect 880 21144 33120 21152
rect 880 21016 33200 21144
rect 880 20872 33120 21016
rect 800 20744 33120 20872
rect 880 20736 33120 20744
rect 880 20608 33200 20736
rect 880 20464 33120 20608
rect 800 20336 33120 20464
rect 880 20328 33120 20336
rect 880 20200 33200 20328
rect 880 20056 33120 20200
rect 800 19928 33120 20056
rect 880 19920 33120 19928
rect 880 19792 33200 19920
rect 880 19648 33120 19792
rect 800 19520 33120 19648
rect 880 19512 33120 19520
rect 880 19384 33200 19512
rect 880 19240 33120 19384
rect 800 19112 33120 19240
rect 880 19104 33120 19112
rect 880 18976 33200 19104
rect 880 18832 33120 18976
rect 800 18704 33120 18832
rect 880 18696 33120 18704
rect 880 18568 33200 18696
rect 880 18424 33120 18568
rect 800 18296 33120 18424
rect 880 18288 33120 18296
rect 880 18160 33200 18288
rect 880 18016 33120 18160
rect 800 17888 33120 18016
rect 880 17880 33120 17888
rect 880 17752 33200 17880
rect 880 17608 33120 17752
rect 800 17480 33120 17608
rect 880 17472 33120 17480
rect 880 17344 33200 17472
rect 880 17200 33120 17344
rect 800 17072 33120 17200
rect 880 17064 33120 17072
rect 880 16936 33200 17064
rect 880 16792 33120 16936
rect 800 16664 33120 16792
rect 880 16656 33120 16664
rect 880 16528 33200 16656
rect 880 16384 33120 16528
rect 800 16256 33120 16384
rect 880 16248 33120 16256
rect 880 16120 33200 16248
rect 880 15976 33120 16120
rect 800 15848 33120 15976
rect 880 15840 33120 15848
rect 880 15712 33200 15840
rect 880 15568 33120 15712
rect 800 15440 33120 15568
rect 880 15432 33120 15440
rect 880 15304 33200 15432
rect 880 15160 33120 15304
rect 800 15032 33120 15160
rect 880 15024 33120 15032
rect 880 14896 33200 15024
rect 880 14752 33120 14896
rect 800 14624 33120 14752
rect 880 14616 33120 14624
rect 880 14488 33200 14616
rect 880 14344 33120 14488
rect 800 14216 33120 14344
rect 880 14208 33120 14216
rect 880 14080 33200 14208
rect 880 13936 33120 14080
rect 800 13808 33120 13936
rect 880 13800 33120 13808
rect 880 13672 33200 13800
rect 880 13528 33120 13672
rect 800 13400 33120 13528
rect 880 13392 33120 13400
rect 880 13264 33200 13392
rect 880 13120 33120 13264
rect 800 12992 33120 13120
rect 880 12984 33120 12992
rect 880 12856 33200 12984
rect 880 12712 33120 12856
rect 800 12584 33120 12712
rect 880 12576 33120 12584
rect 880 12448 33200 12576
rect 880 12304 33120 12448
rect 800 12176 33120 12304
rect 880 12168 33120 12176
rect 880 12040 33200 12168
rect 880 11896 33120 12040
rect 800 11768 33120 11896
rect 880 11760 33120 11768
rect 880 11632 33200 11760
rect 880 11488 33120 11632
rect 800 11360 33120 11488
rect 880 11352 33120 11360
rect 880 11224 33200 11352
rect 880 11080 33120 11224
rect 800 10952 33120 11080
rect 880 10944 33120 10952
rect 880 10816 33200 10944
rect 880 10672 33120 10816
rect 800 10544 33120 10672
rect 880 10536 33120 10544
rect 880 10408 33200 10536
rect 880 10264 33120 10408
rect 800 10136 33120 10264
rect 880 10128 33120 10136
rect 880 10000 33200 10128
rect 880 9856 33120 10000
rect 800 9728 33120 9856
rect 880 9720 33120 9728
rect 880 9592 33200 9720
rect 880 9448 33120 9592
rect 800 9320 33120 9448
rect 880 9312 33120 9320
rect 880 9184 33200 9312
rect 880 9040 33120 9184
rect 800 8912 33120 9040
rect 880 8904 33120 8912
rect 880 8776 33200 8904
rect 880 8632 33120 8776
rect 800 8504 33120 8632
rect 880 8496 33120 8504
rect 880 8368 33200 8496
rect 880 8224 33120 8368
rect 800 8096 33120 8224
rect 880 8088 33120 8096
rect 880 7960 33200 8088
rect 880 7816 33120 7960
rect 800 7688 33120 7816
rect 880 7680 33120 7688
rect 880 7552 33200 7680
rect 880 7408 33120 7552
rect 800 7280 33120 7408
rect 880 7272 33120 7280
rect 880 7144 33200 7272
rect 880 7000 33120 7144
rect 800 6872 33120 7000
rect 880 6864 33120 6872
rect 880 6736 33200 6864
rect 880 6592 33120 6736
rect 800 6464 33120 6592
rect 880 6456 33120 6464
rect 880 6328 33200 6456
rect 880 6184 33120 6328
rect 800 6056 33120 6184
rect 880 6048 33120 6056
rect 880 5920 33200 6048
rect 880 5776 33120 5920
rect 800 5648 33120 5776
rect 880 5640 33120 5648
rect 880 5512 33200 5640
rect 880 5368 33120 5512
rect 800 5240 33120 5368
rect 880 5232 33120 5240
rect 880 5104 33200 5232
rect 880 4960 33120 5104
rect 800 4832 33120 4960
rect 880 4824 33120 4832
rect 880 4696 33200 4824
rect 880 4552 33120 4696
rect 800 4424 33120 4552
rect 880 4416 33120 4424
rect 880 4288 33200 4416
rect 880 4144 33120 4288
rect 800 4016 33120 4144
rect 880 4008 33120 4016
rect 880 3880 33200 4008
rect 880 3736 33120 3880
rect 800 3608 33120 3736
rect 880 3600 33120 3608
rect 880 3472 33200 3600
rect 880 3328 33120 3472
rect 800 3200 33120 3328
rect 880 3192 33120 3200
rect 880 3064 33200 3192
rect 880 2920 33120 3064
rect 800 2792 33120 2920
rect 880 2784 33120 2792
rect 880 2656 33200 2784
rect 880 2512 33120 2656
rect 800 2384 33120 2512
rect 880 2376 33120 2384
rect 880 2248 33200 2376
rect 880 2104 33120 2248
rect 800 1976 33120 2104
rect 880 1968 33120 1976
rect 880 1840 33200 1968
rect 880 1696 33120 1840
rect 800 1568 33120 1696
rect 880 1560 33120 1568
rect 880 1432 33200 1560
rect 880 1288 33120 1432
rect 800 1160 33120 1288
rect 880 1152 33120 1160
rect 880 1024 33200 1152
rect 880 880 33120 1024
rect 800 752 33120 880
rect 880 744 33120 752
rect 880 616 33200 744
rect 880 472 33120 616
rect 800 344 33120 472
rect 880 171 33120 344
<< metal4 >>
rect 6243 2128 6563 53360
rect 11541 2128 11861 53360
rect 16840 2128 17160 53360
rect 22139 2128 22459 53360
rect 27437 2128 27757 53360
<< obsm4 >>
rect 6643 2128 11461 53360
rect 11941 2128 16760 53360
rect 17240 2128 22059 53360
<< labels >>
rlabel metal2 s 6918 -800 6974 800 8 io_adr_i[0]
port 1 nsew signal input
rlabel metal2 s 8482 -800 8538 800 8 io_adr_i[1]
port 2 nsew signal input
rlabel metal2 s 3790 -800 3846 800 8 io_cs_i
port 3 nsew signal input
rlabel metal2 s 9954 -800 10010 800 8 io_dat_i[0]
port 4 nsew signal input
rlabel metal2 s 25502 -800 25558 800 8 io_dat_i[10]
port 5 nsew signal input
rlabel metal2 s 26974 -800 27030 800 8 io_dat_i[11]
port 6 nsew signal input
rlabel metal2 s 28538 -800 28594 800 8 io_dat_i[12]
port 7 nsew signal input
rlabel metal2 s 30102 -800 30158 800 8 io_dat_i[13]
port 8 nsew signal input
rlabel metal2 s 31666 -800 31722 800 8 io_dat_i[14]
port 9 nsew signal input
rlabel metal2 s 33230 -800 33286 800 8 io_dat_i[15]
port 10 nsew signal input
rlabel metal2 s 11518 -800 11574 800 8 io_dat_i[1]
port 11 nsew signal input
rlabel metal2 s 13082 -800 13138 800 8 io_dat_i[2]
port 12 nsew signal input
rlabel metal2 s 14646 -800 14702 800 8 io_dat_i[3]
port 13 nsew signal input
rlabel metal2 s 16210 -800 16266 800 8 io_dat_i[4]
port 14 nsew signal input
rlabel metal2 s 17774 -800 17830 800 8 io_dat_i[5]
port 15 nsew signal input
rlabel metal2 s 19246 -800 19302 800 8 io_dat_i[6]
port 16 nsew signal input
rlabel metal2 s 20810 -800 20866 800 8 io_dat_i[7]
port 17 nsew signal input
rlabel metal2 s 22374 -800 22430 800 8 io_dat_i[8]
port 18 nsew signal input
rlabel metal2 s 23938 -800 23994 800 8 io_dat_i[9]
port 19 nsew signal input
rlabel metal2 s 1030 55200 1086 56800 6 io_dat_o[0]
port 20 nsew signal output
rlabel metal2 s 22282 55200 22338 56800 6 io_dat_o[10]
port 21 nsew signal output
rlabel metal2 s 24398 55200 24454 56800 6 io_dat_o[11]
port 22 nsew signal output
rlabel metal2 s 26514 55200 26570 56800 6 io_dat_o[12]
port 23 nsew signal output
rlabel metal2 s 28630 55200 28686 56800 6 io_dat_o[13]
port 24 nsew signal output
rlabel metal2 s 30746 55200 30802 56800 6 io_dat_o[14]
port 25 nsew signal output
rlabel metal2 s 32862 55200 32918 56800 6 io_dat_o[15]
port 26 nsew signal output
rlabel metal2 s 3146 55200 3202 56800 6 io_dat_o[1]
port 27 nsew signal output
rlabel metal2 s 5262 55200 5318 56800 6 io_dat_o[2]
port 28 nsew signal output
rlabel metal2 s 7378 55200 7434 56800 6 io_dat_o[3]
port 29 nsew signal output
rlabel metal2 s 9494 55200 9550 56800 6 io_dat_o[4]
port 30 nsew signal output
rlabel metal2 s 11610 55200 11666 56800 6 io_dat_o[5]
port 31 nsew signal output
rlabel metal2 s 13726 55200 13782 56800 6 io_dat_o[6]
port 32 nsew signal output
rlabel metal2 s 15842 55200 15898 56800 6 io_dat_o[7]
port 33 nsew signal output
rlabel metal2 s 18050 55200 18106 56800 6 io_dat_o[8]
port 34 nsew signal output
rlabel metal2 s 20166 55200 20222 56800 6 io_dat_o[9]
port 35 nsew signal output
rlabel metal3 s 33200 29248 34800 29368 6 io_eo[0]
port 36 nsew signal input
rlabel metal3 s 33200 33328 34800 33448 6 io_eo[10]
port 37 nsew signal input
rlabel metal3 s 33200 33736 34800 33856 6 io_eo[11]
port 38 nsew signal input
rlabel metal3 s 33200 34144 34800 34264 6 io_eo[12]
port 39 nsew signal input
rlabel metal3 s 33200 34552 34800 34672 6 io_eo[13]
port 40 nsew signal input
rlabel metal3 s 33200 34960 34800 35080 6 io_eo[14]
port 41 nsew signal input
rlabel metal3 s 33200 35368 34800 35488 6 io_eo[15]
port 42 nsew signal input
rlabel metal3 s 33200 35776 34800 35896 6 io_eo[16]
port 43 nsew signal input
rlabel metal3 s 33200 36184 34800 36304 6 io_eo[17]
port 44 nsew signal input
rlabel metal3 s 33200 36592 34800 36712 6 io_eo[18]
port 45 nsew signal input
rlabel metal3 s 33200 37000 34800 37120 6 io_eo[19]
port 46 nsew signal input
rlabel metal3 s 33200 29656 34800 29776 6 io_eo[1]
port 47 nsew signal input
rlabel metal3 s 33200 37408 34800 37528 6 io_eo[20]
port 48 nsew signal input
rlabel metal3 s 33200 37816 34800 37936 6 io_eo[21]
port 49 nsew signal input
rlabel metal3 s 33200 38224 34800 38344 6 io_eo[22]
port 50 nsew signal input
rlabel metal3 s 33200 38632 34800 38752 6 io_eo[23]
port 51 nsew signal input
rlabel metal3 s 33200 39040 34800 39160 6 io_eo[24]
port 52 nsew signal input
rlabel metal3 s 33200 39448 34800 39568 6 io_eo[25]
port 53 nsew signal input
rlabel metal3 s 33200 39856 34800 39976 6 io_eo[26]
port 54 nsew signal input
rlabel metal3 s 33200 40264 34800 40384 6 io_eo[27]
port 55 nsew signal input
rlabel metal3 s 33200 40672 34800 40792 6 io_eo[28]
port 56 nsew signal input
rlabel metal3 s 33200 41080 34800 41200 6 io_eo[29]
port 57 nsew signal input
rlabel metal3 s 33200 30064 34800 30184 6 io_eo[2]
port 58 nsew signal input
rlabel metal3 s 33200 41488 34800 41608 6 io_eo[30]
port 59 nsew signal input
rlabel metal3 s 33200 41896 34800 42016 6 io_eo[31]
port 60 nsew signal input
rlabel metal3 s 33200 42304 34800 42424 6 io_eo[32]
port 61 nsew signal input
rlabel metal3 s 33200 42712 34800 42832 6 io_eo[33]
port 62 nsew signal input
rlabel metal3 s 33200 43120 34800 43240 6 io_eo[34]
port 63 nsew signal input
rlabel metal3 s 33200 43528 34800 43648 6 io_eo[35]
port 64 nsew signal input
rlabel metal3 s 33200 43936 34800 44056 6 io_eo[36]
port 65 nsew signal input
rlabel metal3 s 33200 44344 34800 44464 6 io_eo[37]
port 66 nsew signal input
rlabel metal3 s 33200 44752 34800 44872 6 io_eo[38]
port 67 nsew signal input
rlabel metal3 s 33200 45160 34800 45280 6 io_eo[39]
port 68 nsew signal input
rlabel metal3 s 33200 30472 34800 30592 6 io_eo[3]
port 69 nsew signal input
rlabel metal3 s 33200 45568 34800 45688 6 io_eo[40]
port 70 nsew signal input
rlabel metal3 s 33200 45976 34800 46096 6 io_eo[41]
port 71 nsew signal input
rlabel metal3 s 33200 46384 34800 46504 6 io_eo[42]
port 72 nsew signal input
rlabel metal3 s 33200 46792 34800 46912 6 io_eo[43]
port 73 nsew signal input
rlabel metal3 s 33200 47200 34800 47320 6 io_eo[44]
port 74 nsew signal input
rlabel metal3 s 33200 47608 34800 47728 6 io_eo[45]
port 75 nsew signal input
rlabel metal3 s 33200 48016 34800 48136 6 io_eo[46]
port 76 nsew signal input
rlabel metal3 s 33200 48424 34800 48544 6 io_eo[47]
port 77 nsew signal input
rlabel metal3 s 33200 48832 34800 48952 6 io_eo[48]
port 78 nsew signal input
rlabel metal3 s 33200 49240 34800 49360 6 io_eo[49]
port 79 nsew signal input
rlabel metal3 s 33200 30880 34800 31000 6 io_eo[4]
port 80 nsew signal input
rlabel metal3 s 33200 49648 34800 49768 6 io_eo[50]
port 81 nsew signal input
rlabel metal3 s 33200 50056 34800 50176 6 io_eo[51]
port 82 nsew signal input
rlabel metal3 s 33200 50464 34800 50584 6 io_eo[52]
port 83 nsew signal input
rlabel metal3 s 33200 50872 34800 50992 6 io_eo[53]
port 84 nsew signal input
rlabel metal3 s 33200 51280 34800 51400 6 io_eo[54]
port 85 nsew signal input
rlabel metal3 s 33200 51688 34800 51808 6 io_eo[55]
port 86 nsew signal input
rlabel metal3 s 33200 52096 34800 52216 6 io_eo[56]
port 87 nsew signal input
rlabel metal3 s 33200 52504 34800 52624 6 io_eo[57]
port 88 nsew signal input
rlabel metal3 s 33200 52912 34800 53032 6 io_eo[58]
port 89 nsew signal input
rlabel metal3 s 33200 53320 34800 53440 6 io_eo[59]
port 90 nsew signal input
rlabel metal3 s 33200 31288 34800 31408 6 io_eo[5]
port 91 nsew signal input
rlabel metal3 s 33200 53728 34800 53848 6 io_eo[60]
port 92 nsew signal input
rlabel metal3 s 33200 54136 34800 54256 6 io_eo[61]
port 93 nsew signal input
rlabel metal3 s 33200 54544 34800 54664 6 io_eo[62]
port 94 nsew signal input
rlabel metal3 s 33200 54952 34800 55072 6 io_eo[63]
port 95 nsew signal input
rlabel metal3 s 33200 31696 34800 31816 6 io_eo[6]
port 96 nsew signal input
rlabel metal3 s 33200 32104 34800 32224 6 io_eo[7]
port 97 nsew signal input
rlabel metal3 s 33200 32512 34800 32632 6 io_eo[8]
port 98 nsew signal input
rlabel metal3 s 33200 32920 34800 33040 6 io_eo[9]
port 99 nsew signal input
rlabel metal3 s -800 144 800 264 4 io_i_0_ci
port 100 nsew signal input
rlabel metal3 s -800 3408 800 3528 4 io_i_0_in1[0]
port 101 nsew signal input
rlabel metal3 s -800 6672 800 6792 4 io_i_0_in1[1]
port 102 nsew signal input
rlabel metal3 s -800 9936 800 10056 4 io_i_0_in1[2]
port 103 nsew signal input
rlabel metal3 s -800 13200 800 13320 4 io_i_0_in1[3]
port 104 nsew signal input
rlabel metal3 s -800 16464 800 16584 4 io_i_0_in1[4]
port 105 nsew signal input
rlabel metal3 s -800 19728 800 19848 4 io_i_0_in1[5]
port 106 nsew signal input
rlabel metal3 s -800 22992 800 23112 4 io_i_0_in1[6]
port 107 nsew signal input
rlabel metal3 s -800 26256 800 26376 4 io_i_0_in1[7]
port 108 nsew signal input
rlabel metal3 s -800 552 800 672 4 io_i_1_ci
port 109 nsew signal input
rlabel metal3 s -800 3816 800 3936 4 io_i_1_in1[0]
port 110 nsew signal input
rlabel metal3 s -800 7080 800 7200 4 io_i_1_in1[1]
port 111 nsew signal input
rlabel metal3 s -800 10344 800 10464 4 io_i_1_in1[2]
port 112 nsew signal input
rlabel metal3 s -800 13608 800 13728 4 io_i_1_in1[3]
port 113 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 io_i_1_in1[4]
port 114 nsew signal input
rlabel metal3 s -800 20136 800 20256 4 io_i_1_in1[5]
port 115 nsew signal input
rlabel metal3 s -800 23400 800 23520 4 io_i_1_in1[6]
port 116 nsew signal input
rlabel metal3 s -800 26664 800 26784 4 io_i_1_in1[7]
port 117 nsew signal input
rlabel metal3 s -800 960 800 1080 4 io_i_2_ci
port 118 nsew signal input
rlabel metal3 s -800 4224 800 4344 4 io_i_2_in1[0]
port 119 nsew signal input
rlabel metal3 s -800 7488 800 7608 4 io_i_2_in1[1]
port 120 nsew signal input
rlabel metal3 s -800 10752 800 10872 4 io_i_2_in1[2]
port 121 nsew signal input
rlabel metal3 s -800 14016 800 14136 4 io_i_2_in1[3]
port 122 nsew signal input
rlabel metal3 s -800 17280 800 17400 4 io_i_2_in1[4]
port 123 nsew signal input
rlabel metal3 s -800 20544 800 20664 4 io_i_2_in1[5]
port 124 nsew signal input
rlabel metal3 s -800 23808 800 23928 4 io_i_2_in1[6]
port 125 nsew signal input
rlabel metal3 s -800 27072 800 27192 4 io_i_2_in1[7]
port 126 nsew signal input
rlabel metal3 s -800 1368 800 1488 4 io_i_3_ci
port 127 nsew signal input
rlabel metal3 s -800 4632 800 4752 4 io_i_3_in1[0]
port 128 nsew signal input
rlabel metal3 s -800 7896 800 8016 4 io_i_3_in1[1]
port 129 nsew signal input
rlabel metal3 s -800 11160 800 11280 4 io_i_3_in1[2]
port 130 nsew signal input
rlabel metal3 s -800 14424 800 14544 4 io_i_3_in1[3]
port 131 nsew signal input
rlabel metal3 s -800 17688 800 17808 4 io_i_3_in1[4]
port 132 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 io_i_3_in1[5]
port 133 nsew signal input
rlabel metal3 s -800 24216 800 24336 4 io_i_3_in1[6]
port 134 nsew signal input
rlabel metal3 s -800 27480 800 27600 4 io_i_3_in1[7]
port 135 nsew signal input
rlabel metal3 s -800 1776 800 1896 4 io_i_4_ci
port 136 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 io_i_4_in1[0]
port 137 nsew signal input
rlabel metal3 s -800 8304 800 8424 4 io_i_4_in1[1]
port 138 nsew signal input
rlabel metal3 s -800 11568 800 11688 4 io_i_4_in1[2]
port 139 nsew signal input
rlabel metal3 s -800 14832 800 14952 4 io_i_4_in1[3]
port 140 nsew signal input
rlabel metal3 s -800 18096 800 18216 4 io_i_4_in1[4]
port 141 nsew signal input
rlabel metal3 s -800 21360 800 21480 4 io_i_4_in1[5]
port 142 nsew signal input
rlabel metal3 s -800 24624 800 24744 4 io_i_4_in1[6]
port 143 nsew signal input
rlabel metal3 s -800 27888 800 28008 4 io_i_4_in1[7]
port 144 nsew signal input
rlabel metal3 s -800 2184 800 2304 4 io_i_5_ci
port 145 nsew signal input
rlabel metal3 s -800 5448 800 5568 4 io_i_5_in1[0]
port 146 nsew signal input
rlabel metal3 s -800 8712 800 8832 4 io_i_5_in1[1]
port 147 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 io_i_5_in1[2]
port 148 nsew signal input
rlabel metal3 s -800 15240 800 15360 4 io_i_5_in1[3]
port 149 nsew signal input
rlabel metal3 s -800 18504 800 18624 4 io_i_5_in1[4]
port 150 nsew signal input
rlabel metal3 s -800 21768 800 21888 4 io_i_5_in1[5]
port 151 nsew signal input
rlabel metal3 s -800 25032 800 25152 4 io_i_5_in1[6]
port 152 nsew signal input
rlabel metal3 s -800 28296 800 28416 4 io_i_5_in1[7]
port 153 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 io_i_6_ci
port 154 nsew signal input
rlabel metal3 s -800 5856 800 5976 4 io_i_6_in1[0]
port 155 nsew signal input
rlabel metal3 s -800 9120 800 9240 4 io_i_6_in1[1]
port 156 nsew signal input
rlabel metal3 s -800 12384 800 12504 4 io_i_6_in1[2]
port 157 nsew signal input
rlabel metal3 s -800 15648 800 15768 4 io_i_6_in1[3]
port 158 nsew signal input
rlabel metal3 s -800 18912 800 19032 4 io_i_6_in1[4]
port 159 nsew signal input
rlabel metal3 s -800 22176 800 22296 4 io_i_6_in1[5]
port 160 nsew signal input
rlabel metal3 s -800 25440 800 25560 4 io_i_6_in1[6]
port 161 nsew signal input
rlabel metal3 s -800 28704 800 28824 4 io_i_6_in1[7]
port 162 nsew signal input
rlabel metal3 s -800 3000 800 3120 4 io_i_7_ci
port 163 nsew signal input
rlabel metal3 s -800 6264 800 6384 4 io_i_7_in1[0]
port 164 nsew signal input
rlabel metal3 s -800 9528 800 9648 4 io_i_7_in1[1]
port 165 nsew signal input
rlabel metal3 s -800 12792 800 12912 4 io_i_7_in1[2]
port 166 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 io_i_7_in1[3]
port 167 nsew signal input
rlabel metal3 s -800 19320 800 19440 4 io_i_7_in1[4]
port 168 nsew signal input
rlabel metal3 s -800 22584 800 22704 4 io_i_7_in1[5]
port 169 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 io_i_7_in1[6]
port 170 nsew signal input
rlabel metal3 s -800 29112 800 29232 4 io_i_7_in1[7]
port 171 nsew signal input
rlabel metal3 s 33200 144 34800 264 6 io_o_0_co
port 172 nsew signal output
rlabel metal3 s 33200 3272 34800 3392 6 io_o_0_out[0]
port 173 nsew signal output
rlabel metal3 s 33200 6536 34800 6656 6 io_o_0_out[1]
port 174 nsew signal output
rlabel metal3 s 33200 9800 34800 9920 6 io_o_0_out[2]
port 175 nsew signal output
rlabel metal3 s 33200 13064 34800 13184 6 io_o_0_out[3]
port 176 nsew signal output
rlabel metal3 s 33200 16328 34800 16448 6 io_o_0_out[4]
port 177 nsew signal output
rlabel metal3 s 33200 19592 34800 19712 6 io_o_0_out[5]
port 178 nsew signal output
rlabel metal3 s 33200 22856 34800 22976 6 io_o_0_out[6]
port 179 nsew signal output
rlabel metal3 s 33200 26120 34800 26240 6 io_o_0_out[7]
port 180 nsew signal output
rlabel metal3 s 33200 416 34800 536 6 io_o_1_co
port 181 nsew signal output
rlabel metal3 s 33200 3680 34800 3800 6 io_o_1_out[0]
port 182 nsew signal output
rlabel metal3 s 33200 6944 34800 7064 6 io_o_1_out[1]
port 183 nsew signal output
rlabel metal3 s 33200 10208 34800 10328 6 io_o_1_out[2]
port 184 nsew signal output
rlabel metal3 s 33200 13472 34800 13592 6 io_o_1_out[3]
port 185 nsew signal output
rlabel metal3 s 33200 16736 34800 16856 6 io_o_1_out[4]
port 186 nsew signal output
rlabel metal3 s 33200 20000 34800 20120 6 io_o_1_out[5]
port 187 nsew signal output
rlabel metal3 s 33200 23264 34800 23384 6 io_o_1_out[6]
port 188 nsew signal output
rlabel metal3 s 33200 26528 34800 26648 6 io_o_1_out[7]
port 189 nsew signal output
rlabel metal3 s 33200 824 34800 944 6 io_o_2_co
port 190 nsew signal output
rlabel metal3 s 33200 4088 34800 4208 6 io_o_2_out[0]
port 191 nsew signal output
rlabel metal3 s 33200 7352 34800 7472 6 io_o_2_out[1]
port 192 nsew signal output
rlabel metal3 s 33200 10616 34800 10736 6 io_o_2_out[2]
port 193 nsew signal output
rlabel metal3 s 33200 13880 34800 14000 6 io_o_2_out[3]
port 194 nsew signal output
rlabel metal3 s 33200 17144 34800 17264 6 io_o_2_out[4]
port 195 nsew signal output
rlabel metal3 s 33200 20408 34800 20528 6 io_o_2_out[5]
port 196 nsew signal output
rlabel metal3 s 33200 23672 34800 23792 6 io_o_2_out[6]
port 197 nsew signal output
rlabel metal3 s 33200 26936 34800 27056 6 io_o_2_out[7]
port 198 nsew signal output
rlabel metal3 s 33200 1232 34800 1352 6 io_o_3_co
port 199 nsew signal output
rlabel metal3 s 33200 4496 34800 4616 6 io_o_3_out[0]
port 200 nsew signal output
rlabel metal3 s 33200 7760 34800 7880 6 io_o_3_out[1]
port 201 nsew signal output
rlabel metal3 s 33200 11024 34800 11144 6 io_o_3_out[2]
port 202 nsew signal output
rlabel metal3 s 33200 14288 34800 14408 6 io_o_3_out[3]
port 203 nsew signal output
rlabel metal3 s 33200 17552 34800 17672 6 io_o_3_out[4]
port 204 nsew signal output
rlabel metal3 s 33200 20816 34800 20936 6 io_o_3_out[5]
port 205 nsew signal output
rlabel metal3 s 33200 24080 34800 24200 6 io_o_3_out[6]
port 206 nsew signal output
rlabel metal3 s 33200 27344 34800 27464 6 io_o_3_out[7]
port 207 nsew signal output
rlabel metal3 s 33200 1640 34800 1760 6 io_o_4_co
port 208 nsew signal output
rlabel metal3 s 33200 4904 34800 5024 6 io_o_4_out[0]
port 209 nsew signal output
rlabel metal3 s 33200 8168 34800 8288 6 io_o_4_out[1]
port 210 nsew signal output
rlabel metal3 s 33200 11432 34800 11552 6 io_o_4_out[2]
port 211 nsew signal output
rlabel metal3 s 33200 14696 34800 14816 6 io_o_4_out[3]
port 212 nsew signal output
rlabel metal3 s 33200 17960 34800 18080 6 io_o_4_out[4]
port 213 nsew signal output
rlabel metal3 s 33200 21224 34800 21344 6 io_o_4_out[5]
port 214 nsew signal output
rlabel metal3 s 33200 24488 34800 24608 6 io_o_4_out[6]
port 215 nsew signal output
rlabel metal3 s 33200 27752 34800 27872 6 io_o_4_out[7]
port 216 nsew signal output
rlabel metal3 s 33200 2048 34800 2168 6 io_o_5_co
port 217 nsew signal output
rlabel metal3 s 33200 5312 34800 5432 6 io_o_5_out[0]
port 218 nsew signal output
rlabel metal3 s 33200 8576 34800 8696 6 io_o_5_out[1]
port 219 nsew signal output
rlabel metal3 s 33200 11840 34800 11960 6 io_o_5_out[2]
port 220 nsew signal output
rlabel metal3 s 33200 15104 34800 15224 6 io_o_5_out[3]
port 221 nsew signal output
rlabel metal3 s 33200 18368 34800 18488 6 io_o_5_out[4]
port 222 nsew signal output
rlabel metal3 s 33200 21632 34800 21752 6 io_o_5_out[5]
port 223 nsew signal output
rlabel metal3 s 33200 24896 34800 25016 6 io_o_5_out[6]
port 224 nsew signal output
rlabel metal3 s 33200 28160 34800 28280 6 io_o_5_out[7]
port 225 nsew signal output
rlabel metal3 s 33200 2456 34800 2576 6 io_o_6_co
port 226 nsew signal output
rlabel metal3 s 33200 5720 34800 5840 6 io_o_6_out[0]
port 227 nsew signal output
rlabel metal3 s 33200 8984 34800 9104 6 io_o_6_out[1]
port 228 nsew signal output
rlabel metal3 s 33200 12248 34800 12368 6 io_o_6_out[2]
port 229 nsew signal output
rlabel metal3 s 33200 15512 34800 15632 6 io_o_6_out[3]
port 230 nsew signal output
rlabel metal3 s 33200 18776 34800 18896 6 io_o_6_out[4]
port 231 nsew signal output
rlabel metal3 s 33200 22040 34800 22160 6 io_o_6_out[5]
port 232 nsew signal output
rlabel metal3 s 33200 25304 34800 25424 6 io_o_6_out[6]
port 233 nsew signal output
rlabel metal3 s 33200 28432 34800 28552 6 io_o_6_out[7]
port 234 nsew signal output
rlabel metal3 s 33200 2864 34800 2984 6 io_o_7_co
port 235 nsew signal output
rlabel metal3 s 33200 6128 34800 6248 6 io_o_7_out[0]
port 236 nsew signal output
rlabel metal3 s 33200 9392 34800 9512 6 io_o_7_out[1]
port 237 nsew signal output
rlabel metal3 s 33200 12656 34800 12776 6 io_o_7_out[2]
port 238 nsew signal output
rlabel metal3 s 33200 15920 34800 16040 6 io_o_7_out[3]
port 239 nsew signal output
rlabel metal3 s 33200 19184 34800 19304 6 io_o_7_out[4]
port 240 nsew signal output
rlabel metal3 s 33200 22448 34800 22568 6 io_o_7_out[5]
port 241 nsew signal output
rlabel metal3 s 33200 25712 34800 25832 6 io_o_7_out[6]
port 242 nsew signal output
rlabel metal3 s 33200 28840 34800 28960 6 io_o_7_out[7]
port 243 nsew signal output
rlabel metal2 s 754 -800 810 800 8 io_vci
port 244 nsew signal input
rlabel metal2 s 2226 -800 2282 800 8 io_vco
port 245 nsew signal output
rlabel metal3 s 33200 55360 34800 55480 6 io_vi
port 246 nsew signal input
rlabel metal2 s 5354 -800 5410 800 8 io_we_i
port 247 nsew signal input
rlabel metal3 s -800 29520 800 29640 4 io_wo[0]
port 248 nsew signal output
rlabel metal3 s -800 33600 800 33720 4 io_wo[10]
port 249 nsew signal output
rlabel metal3 s -800 34008 800 34128 4 io_wo[11]
port 250 nsew signal output
rlabel metal3 s -800 34416 800 34536 4 io_wo[12]
port 251 nsew signal output
rlabel metal3 s -800 34824 800 34944 4 io_wo[13]
port 252 nsew signal output
rlabel metal3 s -800 35232 800 35352 4 io_wo[14]
port 253 nsew signal output
rlabel metal3 s -800 35640 800 35760 4 io_wo[15]
port 254 nsew signal output
rlabel metal3 s -800 36048 800 36168 4 io_wo[16]
port 255 nsew signal output
rlabel metal3 s -800 36456 800 36576 4 io_wo[17]
port 256 nsew signal output
rlabel metal3 s -800 36864 800 36984 4 io_wo[18]
port 257 nsew signal output
rlabel metal3 s -800 37272 800 37392 4 io_wo[19]
port 258 nsew signal output
rlabel metal3 s -800 29928 800 30048 4 io_wo[1]
port 259 nsew signal output
rlabel metal3 s -800 37680 800 37800 4 io_wo[20]
port 260 nsew signal output
rlabel metal3 s -800 38088 800 38208 4 io_wo[21]
port 261 nsew signal output
rlabel metal3 s -800 38496 800 38616 4 io_wo[22]
port 262 nsew signal output
rlabel metal3 s -800 38904 800 39024 4 io_wo[23]
port 263 nsew signal output
rlabel metal3 s -800 39312 800 39432 4 io_wo[24]
port 264 nsew signal output
rlabel metal3 s -800 39720 800 39840 4 io_wo[25]
port 265 nsew signal output
rlabel metal3 s -800 40128 800 40248 4 io_wo[26]
port 266 nsew signal output
rlabel metal3 s -800 40536 800 40656 4 io_wo[27]
port 267 nsew signal output
rlabel metal3 s -800 40944 800 41064 4 io_wo[28]
port 268 nsew signal output
rlabel metal3 s -800 41352 800 41472 4 io_wo[29]
port 269 nsew signal output
rlabel metal3 s -800 30336 800 30456 4 io_wo[2]
port 270 nsew signal output
rlabel metal3 s -800 41760 800 41880 4 io_wo[30]
port 271 nsew signal output
rlabel metal3 s -800 42168 800 42288 4 io_wo[31]
port 272 nsew signal output
rlabel metal3 s -800 42576 800 42696 4 io_wo[32]
port 273 nsew signal output
rlabel metal3 s -800 42984 800 43104 4 io_wo[33]
port 274 nsew signal output
rlabel metal3 s -800 43392 800 43512 4 io_wo[34]
port 275 nsew signal output
rlabel metal3 s -800 43800 800 43920 4 io_wo[35]
port 276 nsew signal output
rlabel metal3 s -800 44208 800 44328 4 io_wo[36]
port 277 nsew signal output
rlabel metal3 s -800 44616 800 44736 4 io_wo[37]
port 278 nsew signal output
rlabel metal3 s -800 45024 800 45144 4 io_wo[38]
port 279 nsew signal output
rlabel metal3 s -800 45432 800 45552 4 io_wo[39]
port 280 nsew signal output
rlabel metal3 s -800 30744 800 30864 4 io_wo[3]
port 281 nsew signal output
rlabel metal3 s -800 45840 800 45960 4 io_wo[40]
port 282 nsew signal output
rlabel metal3 s -800 46248 800 46368 4 io_wo[41]
port 283 nsew signal output
rlabel metal3 s -800 46656 800 46776 4 io_wo[42]
port 284 nsew signal output
rlabel metal3 s -800 47064 800 47184 4 io_wo[43]
port 285 nsew signal output
rlabel metal3 s -800 47472 800 47592 4 io_wo[44]
port 286 nsew signal output
rlabel metal3 s -800 47880 800 48000 4 io_wo[45]
port 287 nsew signal output
rlabel metal3 s -800 48288 800 48408 4 io_wo[46]
port 288 nsew signal output
rlabel metal3 s -800 48696 800 48816 4 io_wo[47]
port 289 nsew signal output
rlabel metal3 s -800 49104 800 49224 4 io_wo[48]
port 290 nsew signal output
rlabel metal3 s -800 49512 800 49632 4 io_wo[49]
port 291 nsew signal output
rlabel metal3 s -800 31152 800 31272 4 io_wo[4]
port 292 nsew signal output
rlabel metal3 s -800 49920 800 50040 4 io_wo[50]
port 293 nsew signal output
rlabel metal3 s -800 50328 800 50448 4 io_wo[51]
port 294 nsew signal output
rlabel metal3 s -800 50736 800 50856 4 io_wo[52]
port 295 nsew signal output
rlabel metal3 s -800 51144 800 51264 4 io_wo[53]
port 296 nsew signal output
rlabel metal3 s -800 51552 800 51672 4 io_wo[54]
port 297 nsew signal output
rlabel metal3 s -800 51960 800 52080 4 io_wo[55]
port 298 nsew signal output
rlabel metal3 s -800 52368 800 52488 4 io_wo[56]
port 299 nsew signal output
rlabel metal3 s -800 52776 800 52896 4 io_wo[57]
port 300 nsew signal output
rlabel metal3 s -800 53184 800 53304 4 io_wo[58]
port 301 nsew signal output
rlabel metal3 s -800 53592 800 53712 4 io_wo[59]
port 302 nsew signal output
rlabel metal3 s -800 31560 800 31680 4 io_wo[5]
port 303 nsew signal output
rlabel metal3 s -800 54000 800 54120 4 io_wo[60]
port 304 nsew signal output
rlabel metal3 s -800 54408 800 54528 4 io_wo[61]
port 305 nsew signal output
rlabel metal3 s -800 54816 800 54936 4 io_wo[62]
port 306 nsew signal output
rlabel metal3 s -800 55224 800 55344 4 io_wo[63]
port 307 nsew signal output
rlabel metal3 s -800 31968 800 32088 4 io_wo[6]
port 308 nsew signal output
rlabel metal3 s -800 32376 800 32496 4 io_wo[7]
port 309 nsew signal output
rlabel metal3 s -800 32784 800 32904 4 io_wo[8]
port 310 nsew signal output
rlabel metal3 s -800 33192 800 33312 4 io_wo[9]
port 311 nsew signal output
rlabel metal3 s -800 55632 800 55752 4 wb_clk_i
port 312 nsew signal input
rlabel metal3 s 33200 55768 34800 55888 6 wb_rst_i
port 313 nsew signal input
rlabel metal4 s 27437 2128 27757 53360 6 vccd1
port 314 nsew power bidirectional
rlabel metal4 s 16840 2128 17160 53360 6 vccd1
port 315 nsew power bidirectional
rlabel metal4 s 6243 2128 6563 53360 6 vccd1
port 316 nsew power bidirectional
rlabel metal4 s 22139 2128 22459 53360 6 vssd1
port 317 nsew ground bidirectional
rlabel metal4 s 11541 2128 11861 53360 6 vssd1
port 318 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 34000 56000
string LEFview TRUE
string GDS_FILE /project/openlane/cic_block/runs/cic_block/results/magic/cic_block.gds
string GDS_END 6385102
string GDS_START 660770
<< end >>

