VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_local
  CLASS BLOCK ;
  FOREIGN wb_local ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 600.000 ;
  PIN dsi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 596.000 0.830 604.000 ;
    END
  END dsi[0]
  PIN dsi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 596.000 1.750 604.000 ;
    END
  END dsi[1]
  PIN dsi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 596.000 2.670 604.000 ;
    END
  END dsi[2]
  PIN dsi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 596.000 3.590 604.000 ;
    END
  END dsi[3]
  PIN dsi[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 596.000 4.970 604.000 ;
    END
  END dsi[4]
  PIN dsi[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 596.000 5.890 604.000 ;
    END
  END dsi[5]
  PIN dsi[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 596.000 6.810 604.000 ;
    END
  END dsi[6]
  PIN dsi[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 596.000 8.190 604.000 ;
    END
  END dsi[7]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 596.000 9.110 604.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 596.000 40.850 604.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 596.000 44.070 604.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 596.000 47.290 604.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 596.000 50.510 604.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 596.000 53.730 604.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 596.000 56.490 604.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 596.000 59.710 604.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 596.000 62.930 604.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 596.000 66.150 604.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 596.000 69.370 604.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 596.000 12.330 604.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 596.000 72.590 604.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 596.000 75.810 604.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 596.000 79.030 604.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 596.000 82.250 604.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 596.000 85.470 604.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 596.000 88.690 604.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 596.000 91.450 604.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 596.000 94.670 604.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 596.000 97.890 604.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 596.000 101.110 604.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 596.000 15.550 604.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 596.000 104.330 604.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 596.000 107.550 604.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 596.000 110.770 604.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 596.000 113.990 604.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 596.000 117.210 604.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 596.000 120.430 604.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 596.000 123.190 604.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 596.000 126.410 604.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 596.000 18.770 604.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 596.000 21.990 604.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 596.000 24.750 604.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 596.000 27.970 604.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 596.000 31.190 604.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 596.000 34.410 604.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 596.000 37.630 604.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 596.000 10.030 604.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 596.000 41.770 604.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 596.000 44.990 604.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 596.000 48.210 604.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 596.000 51.430 604.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 596.000 54.650 604.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 596.000 57.870 604.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 596.000 61.090 604.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 596.000 64.310 604.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 596.000 67.530 604.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 596.000 70.290 604.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 596.000 13.250 604.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 596.000 73.510 604.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 596.000 76.730 604.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 596.000 79.950 604.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 596.000 83.170 604.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 596.000 86.390 604.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 596.000 89.610 604.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 596.000 92.830 604.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 596.000 96.050 604.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 596.000 99.270 604.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 596.000 102.030 604.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 596.000 16.470 604.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 596.000 105.250 604.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 596.000 108.470 604.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 596.000 111.690 604.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 596.000 114.910 604.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 596.000 118.130 604.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 596.000 121.350 604.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 596.000 124.570 604.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 596.000 127.790 604.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 596.000 19.690 604.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 596.000 22.910 604.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 596.000 26.130 604.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 596.000 29.350 604.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 596.000 32.570 604.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 596.000 35.330 604.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 596.000 38.550 604.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 596.000 11.410 604.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 596.000 43.150 604.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 596.000 45.910 604.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 596.000 49.130 604.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 596.000 52.350 604.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 596.000 55.570 604.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 596.000 58.790 604.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 596.000 62.010 604.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 596.000 65.230 604.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 596.000 68.450 604.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 596.000 71.670 604.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 596.000 14.170 604.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 596.000 74.890 604.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 596.000 78.110 604.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 596.000 80.870 604.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 596.000 84.090 604.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 596.000 87.310 604.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 596.000 90.530 604.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 596.000 93.750 604.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 596.000 96.970 604.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 596.000 100.190 604.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 596.000 103.410 604.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 596.000 17.390 604.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 596.000 106.630 604.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 596.000 109.850 604.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 596.000 112.610 604.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 596.000 115.830 604.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 596.000 119.050 604.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 596.000 122.270 604.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 596.000 125.490 604.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 596.000 128.710 604.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 596.000 20.610 604.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 596.000 23.830 604.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 596.000 27.050 604.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 596.000 30.270 604.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 596.000 33.490 604.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 596.000 36.710 604.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 596.000 39.930 604.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 -4.000 3.590 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 -4.000 4.970 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 -4.000 6.350 4.000 ;
    END
  END irq[2]
  PIN la_reset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 -4.000 159.990 4.000 ;
    END
  END la_reset[0]
  PIN la_reset[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 -4.000 174.250 4.000 ;
    END
  END la_reset[10]
  PIN la_reset[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 -4.000 176.090 4.000 ;
    END
  END la_reset[11]
  PIN la_reset[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 -4.000 161.370 4.000 ;
    END
  END la_reset[1]
  PIN la_reset[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 -4.000 162.750 4.000 ;
    END
  END la_reset[2]
  PIN la_reset[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 -4.000 164.130 4.000 ;
    END
  END la_reset[3]
  PIN la_reset[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 -4.000 165.510 4.000 ;
    END
  END la_reset[4]
  PIN la_reset[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 -4.000 166.890 4.000 ;
    END
  END la_reset[5]
  PIN la_reset[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 -4.000 168.730 4.000 ;
    END
  END la_reset[6]
  PIN la_reset[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 -4.000 170.110 4.000 ;
    END
  END la_reset[7]
  PIN la_reset[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 -4.000 171.490 4.000 ;
    END
  END la_reset[8]
  PIN la_reset[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 -4.000 172.870 4.000 ;
    END
  END la_reset[9]
  PIN m_irqs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 596.000 158.150 604.000 ;
    END
  END m_irqs[0]
  PIN m_irqs[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 596.000 168.730 604.000 ;
    END
  END m_irqs[10]
  PIN m_irqs[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 596.000 170.110 604.000 ;
    END
  END m_irqs[11]
  PIN m_irqs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 596.000 159.530 604.000 ;
    END
  END m_irqs[1]
  PIN m_irqs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 596.000 160.450 604.000 ;
    END
  END m_irqs[2]
  PIN m_irqs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 596.000 161.370 604.000 ;
    END
  END m_irqs[3]
  PIN m_irqs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 596.000 162.750 604.000 ;
    END
  END m_irqs[4]
  PIN m_irqs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 596.000 163.670 604.000 ;
    END
  END m_irqs[5]
  PIN m_irqs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 596.000 164.590 604.000 ;
    END
  END m_irqs[6]
  PIN m_irqs[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 596.000 165.970 604.000 ;
    END
  END m_irqs[7]
  PIN m_irqs[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 596.000 166.890 604.000 ;
    END
  END m_irqs[8]
  PIN m_irqs[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 596.000 167.810 604.000 ;
    END
  END m_irqs[9]
  PIN m_la_reset[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 596.000 171.030 604.000 ;
    END
  END m_la_reset[0]
  PIN m_la_reset[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 596.000 181.610 604.000 ;
    END
  END m_la_reset[10]
  PIN m_la_reset[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 596.000 182.530 604.000 ;
    END
  END m_la_reset[11]
  PIN m_la_reset[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 596.000 171.950 604.000 ;
    END
  END m_la_reset[1]
  PIN m_la_reset[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 596.000 173.330 604.000 ;
    END
  END m_la_reset[2]
  PIN m_la_reset[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 596.000 174.250 604.000 ;
    END
  END m_la_reset[3]
  PIN m_la_reset[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 596.000 175.170 604.000 ;
    END
  END m_la_reset[4]
  PIN m_la_reset[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 596.000 176.550 604.000 ;
    END
  END m_la_reset[5]
  PIN m_la_reset[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 596.000 177.470 604.000 ;
    END
  END m_la_reset[6]
  PIN m_la_reset[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 596.000 178.390 604.000 ;
    END
  END m_la_reset[7]
  PIN m_la_reset[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 596.000 179.310 604.000 ;
    END
  END m_la_reset[8]
  PIN m_la_reset[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 596.000 180.690 604.000 ;
    END
  END m_la_reset[9]
  PIN m_wb_clk_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 -4.000 177.470 4.000 ;
    END
  END m_wb_clk_i
  PIN m_wb_rst_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 531.120 4.000 531.720 ;
    END
  END m_wb_rst_i
  PIN m_wbs_ack_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 552.880 204.000 553.480 ;
    END
  END m_wbs_ack_o[0]
  PIN m_wbs_ack_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 -4.000 191.730 4.000 ;
    END
  END m_wbs_ack_o[10]
  PIN m_wbs_ack_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 582.800 204.000 583.400 ;
    END
  END m_wbs_ack_o[11]
  PIN m_wbs_ack_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 559.000 204.000 559.600 ;
    END
  END m_wbs_ack_o[1]
  PIN m_wbs_ack_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 -4.000 178.850 4.000 ;
    END
  END m_wbs_ack_o[2]
  PIN m_wbs_ack_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 596.000 185.750 604.000 ;
    END
  END m_wbs_ack_o[3]
  PIN m_wbs_ack_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 -4.000 182.990 4.000 ;
    END
  END m_wbs_ack_o[4]
  PIN m_wbs_ack_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 571.920 204.000 572.520 ;
    END
  END m_wbs_ack_o[5]
  PIN m_wbs_ack_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 596.000 188.970 604.000 ;
    END
  END m_wbs_ack_o[6]
  PIN m_wbs_ack_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 576.680 204.000 577.280 ;
    END
  END m_wbs_ack_o[7]
  PIN m_wbs_ack_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.280 4.000 556.880 ;
    END
  END m_wbs_ack_o[8]
  PIN m_wbs_ack_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 564.440 4.000 565.040 ;
    END
  END m_wbs_ack_o[9]
  PIN m_wbs_adr_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 554.920 204.000 555.520 ;
    END
  END m_wbs_adr_i[0]
  PIN m_wbs_adr_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 572.600 4.000 573.200 ;
    END
  END m_wbs_adr_i[10]
  PIN m_wbs_adr_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 584.840 204.000 585.440 ;
    END
  END m_wbs_adr_i[11]
  PIN m_wbs_adr_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 561.040 204.000 561.640 ;
    END
  END m_wbs_adr_i[1]
  PIN m_wbs_adr_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 -4.000 180.230 4.000 ;
    END
  END m_wbs_adr_i[2]
  PIN m_wbs_adr_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 563.760 204.000 564.360 ;
    END
  END m_wbs_adr_i[3]
  PIN m_wbs_adr_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 -4.000 184.830 4.000 ;
    END
  END m_wbs_adr_i[4]
  PIN m_wbs_adr_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 -4.000 186.210 4.000 ;
    END
  END m_wbs_adr_i[5]
  PIN m_wbs_adr_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 596.000 189.890 604.000 ;
    END
  END m_wbs_adr_i[6]
  PIN m_wbs_adr_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 578.720 204.000 579.320 ;
    END
  END m_wbs_adr_i[7]
  PIN m_wbs_adr_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 596.000 191.270 604.000 ;
    END
  END m_wbs_adr_i[8]
  PIN m_wbs_adr_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 568.520 4.000 569.120 ;
    END
  END m_wbs_adr_i[9]
  PIN m_wbs_cs_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 535.200 4.000 535.800 ;
    END
  END m_wbs_cs_i[0]
  PIN m_wbs_cs_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 576.680 4.000 577.280 ;
    END
  END m_wbs_cs_i[10]
  PIN m_wbs_cs_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 -4.000 193.570 4.000 ;
    END
  END m_wbs_cs_i[11]
  PIN m_wbs_cs_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 539.280 4.000 539.880 ;
    END
  END m_wbs_cs_i[1]
  PIN m_wbs_cs_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 543.360 4.000 543.960 ;
    END
  END m_wbs_cs_i[2]
  PIN m_wbs_cs_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 565.800 204.000 566.400 ;
    END
  END m_wbs_cs_i[3]
  PIN m_wbs_cs_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 569.880 204.000 570.480 ;
    END
  END m_wbs_cs_i[4]
  PIN m_wbs_cs_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 547.440 4.000 548.040 ;
    END
  END m_wbs_cs_i[5]
  PIN m_wbs_cs_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 573.960 204.000 574.560 ;
    END
  END m_wbs_cs_i[6]
  PIN m_wbs_cs_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 -4.000 188.970 4.000 ;
    END
  END m_wbs_cs_i[7]
  PIN m_wbs_cs_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 560.360 4.000 560.960 ;
    END
  END m_wbs_cs_i[8]
  PIN m_wbs_cs_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 -4.000 190.350 4.000 ;
    END
  END m_wbs_cs_i[9]
  PIN m_wbs_dat_i[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 556.960 204.000 557.560 ;
    END
  END m_wbs_dat_i[0]
  PIN m_wbs_dat_i[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 580.760 204.000 581.360 ;
    END
  END m_wbs_dat_i[10]
  PIN m_wbs_dat_i[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 580.760 4.000 581.360 ;
    END
  END m_wbs_dat_i[11]
  PIN m_wbs_dat_i[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 -4.000 194.950 4.000 ;
    END
  END m_wbs_dat_i[12]
  PIN m_wbs_dat_i[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.840 4.000 585.440 ;
    END
  END m_wbs_dat_i[13]
  PIN m_wbs_dat_i[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 596.000 194.490 604.000 ;
    END
  END m_wbs_dat_i[14]
  PIN m_wbs_dat_i[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 588.920 4.000 589.520 ;
    END
  END m_wbs_dat_i[15]
  PIN m_wbs_dat_i[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 596.000 195.410 604.000 ;
    END
  END m_wbs_dat_i[16]
  PIN m_wbs_dat_i[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 586.880 204.000 587.480 ;
    END
  END m_wbs_dat_i[17]
  PIN m_wbs_dat_i[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 596.000 196.330 604.000 ;
    END
  END m_wbs_dat_i[18]
  PIN m_wbs_dat_i[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 596.000 197.710 604.000 ;
    END
  END m_wbs_dat_i[19]
  PIN m_wbs_dat_i[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 596.000 184.830 604.000 ;
    END
  END m_wbs_dat_i[1]
  PIN m_wbs_dat_i[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 593.000 4.000 593.600 ;
    END
  END m_wbs_dat_i[20]
  PIN m_wbs_dat_i[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 -4.000 196.330 4.000 ;
    END
  END m_wbs_dat_i[21]
  PIN m_wbs_dat_i[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 589.600 204.000 590.200 ;
    END
  END m_wbs_dat_i[22]
  PIN m_wbs_dat_i[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 591.640 204.000 592.240 ;
    END
  END m_wbs_dat_i[23]
  PIN m_wbs_dat_i[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 -4.000 197.710 4.000 ;
    END
  END m_wbs_dat_i[24]
  PIN m_wbs_dat_i[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 596.000 198.630 604.000 ;
    END
  END m_wbs_dat_i[25]
  PIN m_wbs_dat_i[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 593.680 204.000 594.280 ;
    END
  END m_wbs_dat_i[26]
  PIN m_wbs_dat_i[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 595.720 204.000 596.320 ;
    END
  END m_wbs_dat_i[27]
  PIN m_wbs_dat_i[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 597.760 204.000 598.360 ;
    END
  END m_wbs_dat_i[28]
  PIN m_wbs_dat_i[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 596.000 199.550 604.000 ;
    END
  END m_wbs_dat_i[29]
  PIN m_wbs_dat_i[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 -4.000 181.610 4.000 ;
    END
  END m_wbs_dat_i[2]
  PIN m_wbs_dat_i[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 597.080 4.000 597.680 ;
    END
  END m_wbs_dat_i[30]
  PIN m_wbs_dat_i[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 -4.000 199.090 4.000 ;
    END
  END m_wbs_dat_i[31]
  PIN m_wbs_dat_i[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 567.840 204.000 568.440 ;
    END
  END m_wbs_dat_i[3]
  PIN m_wbs_dat_i[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 596.000 187.130 604.000 ;
    END
  END m_wbs_dat_i[4]
  PIN m_wbs_dat_i[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 596.000 188.050 604.000 ;
    END
  END m_wbs_dat_i[5]
  PIN m_wbs_dat_i[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 -4.000 187.590 4.000 ;
    END
  END m_wbs_dat_i[6]
  PIN m_wbs_dat_i[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 552.200 4.000 552.800 ;
    END
  END m_wbs_dat_i[7]
  PIN m_wbs_dat_i[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 596.000 192.190 604.000 ;
    END
  END m_wbs_dat_i[8]
  PIN m_wbs_dat_i[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 596.000 193.110 604.000 ;
    END
  END m_wbs_dat_i[9]
  PIN m_wbs_dat_o_0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 0.720 204.000 1.320 ;
    END
  END m_wbs_dat_o_0[0]
  PIN m_wbs_dat_o_0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 21.800 204.000 22.400 ;
    END
  END m_wbs_dat_o_0[10]
  PIN m_wbs_dat_o_0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 204.000 24.440 ;
    END
  END m_wbs_dat_o_0[11]
  PIN m_wbs_dat_o_0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 26.560 204.000 27.160 ;
    END
  END m_wbs_dat_o_0[12]
  PIN m_wbs_dat_o_0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 28.600 204.000 29.200 ;
    END
  END m_wbs_dat_o_0[13]
  PIN m_wbs_dat_o_0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 30.640 204.000 31.240 ;
    END
  END m_wbs_dat_o_0[14]
  PIN m_wbs_dat_o_0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.680 204.000 33.280 ;
    END
  END m_wbs_dat_o_0[15]
  PIN m_wbs_dat_o_0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.720 204.000 35.320 ;
    END
  END m_wbs_dat_o_0[16]
  PIN m_wbs_dat_o_0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 36.760 204.000 37.360 ;
    END
  END m_wbs_dat_o_0[17]
  PIN m_wbs_dat_o_0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 39.480 204.000 40.080 ;
    END
  END m_wbs_dat_o_0[18]
  PIN m_wbs_dat_o_0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 41.520 204.000 42.120 ;
    END
  END m_wbs_dat_o_0[19]
  PIN m_wbs_dat_o_0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2.760 204.000 3.360 ;
    END
  END m_wbs_dat_o_0[1]
  PIN m_wbs_dat_o_0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 43.560 204.000 44.160 ;
    END
  END m_wbs_dat_o_0[20]
  PIN m_wbs_dat_o_0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 45.600 204.000 46.200 ;
    END
  END m_wbs_dat_o_0[21]
  PIN m_wbs_dat_o_0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 47.640 204.000 48.240 ;
    END
  END m_wbs_dat_o_0[22]
  PIN m_wbs_dat_o_0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 49.680 204.000 50.280 ;
    END
  END m_wbs_dat_o_0[23]
  PIN m_wbs_dat_o_0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 52.400 204.000 53.000 ;
    END
  END m_wbs_dat_o_0[24]
  PIN m_wbs_dat_o_0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 54.440 204.000 55.040 ;
    END
  END m_wbs_dat_o_0[25]
  PIN m_wbs_dat_o_0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 56.480 204.000 57.080 ;
    END
  END m_wbs_dat_o_0[26]
  PIN m_wbs_dat_o_0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 58.520 204.000 59.120 ;
    END
  END m_wbs_dat_o_0[27]
  PIN m_wbs_dat_o_0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 60.560 204.000 61.160 ;
    END
  END m_wbs_dat_o_0[28]
  PIN m_wbs_dat_o_0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 63.280 204.000 63.880 ;
    END
  END m_wbs_dat_o_0[29]
  PIN m_wbs_dat_o_0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 4.800 204.000 5.400 ;
    END
  END m_wbs_dat_o_0[2]
  PIN m_wbs_dat_o_0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 65.320 204.000 65.920 ;
    END
  END m_wbs_dat_o_0[30]
  PIN m_wbs_dat_o_0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 67.360 204.000 67.960 ;
    END
  END m_wbs_dat_o_0[31]
  PIN m_wbs_dat_o_0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 6.840 204.000 7.440 ;
    END
  END m_wbs_dat_o_0[3]
  PIN m_wbs_dat_o_0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 8.880 204.000 9.480 ;
    END
  END m_wbs_dat_o_0[4]
  PIN m_wbs_dat_o_0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 10.920 204.000 11.520 ;
    END
  END m_wbs_dat_o_0[5]
  PIN m_wbs_dat_o_0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 13.640 204.000 14.240 ;
    END
  END m_wbs_dat_o_0[6]
  PIN m_wbs_dat_o_0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 15.680 204.000 16.280 ;
    END
  END m_wbs_dat_o_0[7]
  PIN m_wbs_dat_o_0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 17.720 204.000 18.320 ;
    END
  END m_wbs_dat_o_0[8]
  PIN m_wbs_dat_o_0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 19.760 204.000 20.360 ;
    END
  END m_wbs_dat_o_0[9]
  PIN m_wbs_dat_o_10[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 204.000 72.040 ;
    END
  END m_wbs_dat_o_10[0]
  PIN m_wbs_dat_o_10[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 136.040 204.000 136.640 ;
    END
  END m_wbs_dat_o_10[10]
  PIN m_wbs_dat_o_10[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 142.840 204.000 143.440 ;
    END
  END m_wbs_dat_o_10[11]
  PIN m_wbs_dat_o_10[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.960 204.000 149.560 ;
    END
  END m_wbs_dat_o_10[12]
  PIN m_wbs_dat_o_10[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.760 204.000 156.360 ;
    END
  END m_wbs_dat_o_10[13]
  PIN m_wbs_dat_o_10[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 161.880 204.000 162.480 ;
    END
  END m_wbs_dat_o_10[14]
  PIN m_wbs_dat_o_10[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 204.000 169.280 ;
    END
  END m_wbs_dat_o_10[15]
  PIN m_wbs_dat_o_10[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.800 204.000 175.400 ;
    END
  END m_wbs_dat_o_10[16]
  PIN m_wbs_dat_o_10[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 181.600 204.000 182.200 ;
    END
  END m_wbs_dat_o_10[17]
  PIN m_wbs_dat_o_10[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 188.400 204.000 189.000 ;
    END
  END m_wbs_dat_o_10[18]
  PIN m_wbs_dat_o_10[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 194.520 204.000 195.120 ;
    END
  END m_wbs_dat_o_10[19]
  PIN m_wbs_dat_o_10[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 204.000 78.840 ;
    END
  END m_wbs_dat_o_10[1]
  PIN m_wbs_dat_o_10[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 201.320 204.000 201.920 ;
    END
  END m_wbs_dat_o_10[20]
  PIN m_wbs_dat_o_10[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 207.440 204.000 208.040 ;
    END
  END m_wbs_dat_o_10[21]
  PIN m_wbs_dat_o_10[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 214.240 204.000 214.840 ;
    END
  END m_wbs_dat_o_10[22]
  PIN m_wbs_dat_o_10[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 220.360 204.000 220.960 ;
    END
  END m_wbs_dat_o_10[23]
  PIN m_wbs_dat_o_10[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 227.160 204.000 227.760 ;
    END
  END m_wbs_dat_o_10[24]
  PIN m_wbs_dat_o_10[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 233.280 204.000 233.880 ;
    END
  END m_wbs_dat_o_10[25]
  PIN m_wbs_dat_o_10[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 240.080 204.000 240.680 ;
    END
  END m_wbs_dat_o_10[26]
  PIN m_wbs_dat_o_10[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 246.200 204.000 246.800 ;
    END
  END m_wbs_dat_o_10[27]
  PIN m_wbs_dat_o_10[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 253.000 204.000 253.600 ;
    END
  END m_wbs_dat_o_10[28]
  PIN m_wbs_dat_o_10[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 259.120 204.000 259.720 ;
    END
  END m_wbs_dat_o_10[29]
  PIN m_wbs_dat_o_10[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 84.360 204.000 84.960 ;
    END
  END m_wbs_dat_o_10[2]
  PIN m_wbs_dat_o_10[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 265.920 204.000 266.520 ;
    END
  END m_wbs_dat_o_10[30]
  PIN m_wbs_dat_o_10[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 272.040 204.000 272.640 ;
    END
  END m_wbs_dat_o_10[31]
  PIN m_wbs_dat_o_10[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.160 204.000 91.760 ;
    END
  END m_wbs_dat_o_10[3]
  PIN m_wbs_dat_o_10[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 97.280 204.000 97.880 ;
    END
  END m_wbs_dat_o_10[4]
  PIN m_wbs_dat_o_10[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 104.080 204.000 104.680 ;
    END
  END m_wbs_dat_o_10[5]
  PIN m_wbs_dat_o_10[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 110.200 204.000 110.800 ;
    END
  END m_wbs_dat_o_10[6]
  PIN m_wbs_dat_o_10[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 117.000 204.000 117.600 ;
    END
  END m_wbs_dat_o_10[7]
  PIN m_wbs_dat_o_10[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 123.120 204.000 123.720 ;
    END
  END m_wbs_dat_o_10[8]
  PIN m_wbs_dat_o_10[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.920 204.000 130.520 ;
    END
  END m_wbs_dat_o_10[9]
  PIN m_wbs_dat_o_11[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 73.480 204.000 74.080 ;
    END
  END m_wbs_dat_o_11[0]
  PIN m_wbs_dat_o_11[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 138.760 204.000 139.360 ;
    END
  END m_wbs_dat_o_11[10]
  PIN m_wbs_dat_o_11[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 144.880 204.000 145.480 ;
    END
  END m_wbs_dat_o_11[11]
  PIN m_wbs_dat_o_11[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 151.680 204.000 152.280 ;
    END
  END m_wbs_dat_o_11[12]
  PIN m_wbs_dat_o_11[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.800 204.000 158.400 ;
    END
  END m_wbs_dat_o_11[13]
  PIN m_wbs_dat_o_11[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 164.600 204.000 165.200 ;
    END
  END m_wbs_dat_o_11[14]
  PIN m_wbs_dat_o_11[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 170.720 204.000 171.320 ;
    END
  END m_wbs_dat_o_11[15]
  PIN m_wbs_dat_o_11[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 177.520 204.000 178.120 ;
    END
  END m_wbs_dat_o_11[16]
  PIN m_wbs_dat_o_11[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 204.000 184.240 ;
    END
  END m_wbs_dat_o_11[17]
  PIN m_wbs_dat_o_11[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 204.000 191.040 ;
    END
  END m_wbs_dat_o_11[18]
  PIN m_wbs_dat_o_11[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 196.560 204.000 197.160 ;
    END
  END m_wbs_dat_o_11[19]
  PIN m_wbs_dat_o_11[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 80.280 204.000 80.880 ;
    END
  END m_wbs_dat_o_11[1]
  PIN m_wbs_dat_o_11[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 203.360 204.000 203.960 ;
    END
  END m_wbs_dat_o_11[20]
  PIN m_wbs_dat_o_11[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 209.480 204.000 210.080 ;
    END
  END m_wbs_dat_o_11[21]
  PIN m_wbs_dat_o_11[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 216.280 204.000 216.880 ;
    END
  END m_wbs_dat_o_11[22]
  PIN m_wbs_dat_o_11[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 222.400 204.000 223.000 ;
    END
  END m_wbs_dat_o_11[23]
  PIN m_wbs_dat_o_11[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 229.200 204.000 229.800 ;
    END
  END m_wbs_dat_o_11[24]
  PIN m_wbs_dat_o_11[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 235.320 204.000 235.920 ;
    END
  END m_wbs_dat_o_11[25]
  PIN m_wbs_dat_o_11[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 242.120 204.000 242.720 ;
    END
  END m_wbs_dat_o_11[26]
  PIN m_wbs_dat_o_11[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 248.240 204.000 248.840 ;
    END
  END m_wbs_dat_o_11[27]
  PIN m_wbs_dat_o_11[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.040 204.000 255.640 ;
    END
  END m_wbs_dat_o_11[28]
  PIN m_wbs_dat_o_11[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 261.160 204.000 261.760 ;
    END
  END m_wbs_dat_o_11[29]
  PIN m_wbs_dat_o_11[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 86.400 204.000 87.000 ;
    END
  END m_wbs_dat_o_11[2]
  PIN m_wbs_dat_o_11[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 267.960 204.000 268.560 ;
    END
  END m_wbs_dat_o_11[30]
  PIN m_wbs_dat_o_11[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 274.080 204.000 274.680 ;
    END
  END m_wbs_dat_o_11[31]
  PIN m_wbs_dat_o_11[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 93.200 204.000 93.800 ;
    END
  END m_wbs_dat_o_11[3]
  PIN m_wbs_dat_o_11[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 99.320 204.000 99.920 ;
    END
  END m_wbs_dat_o_11[4]
  PIN m_wbs_dat_o_11[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 106.120 204.000 106.720 ;
    END
  END m_wbs_dat_o_11[5]
  PIN m_wbs_dat_o_11[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 112.240 204.000 112.840 ;
    END
  END m_wbs_dat_o_11[6]
  PIN m_wbs_dat_o_11[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 119.040 204.000 119.640 ;
    END
  END m_wbs_dat_o_11[7]
  PIN m_wbs_dat_o_11[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 204.000 126.440 ;
    END
  END m_wbs_dat_o_11[8]
  PIN m_wbs_dat_o_11[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 131.960 204.000 132.560 ;
    END
  END m_wbs_dat_o_11[9]
  PIN m_wbs_dat_o_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 69.400 204.000 70.000 ;
    END
  END m_wbs_dat_o_1[0]
  PIN m_wbs_dat_o_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 134.000 204.000 134.600 ;
    END
  END m_wbs_dat_o_1[10]
  PIN m_wbs_dat_o_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 140.800 204.000 141.400 ;
    END
  END m_wbs_dat_o_1[11]
  PIN m_wbs_dat_o_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 146.920 204.000 147.520 ;
    END
  END m_wbs_dat_o_1[12]
  PIN m_wbs_dat_o_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 153.720 204.000 154.320 ;
    END
  END m_wbs_dat_o_1[13]
  PIN m_wbs_dat_o_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 159.840 204.000 160.440 ;
    END
  END m_wbs_dat_o_1[14]
  PIN m_wbs_dat_o_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 166.640 204.000 167.240 ;
    END
  END m_wbs_dat_o_1[15]
  PIN m_wbs_dat_o_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 172.760 204.000 173.360 ;
    END
  END m_wbs_dat_o_1[16]
  PIN m_wbs_dat_o_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 204.000 180.160 ;
    END
  END m_wbs_dat_o_1[17]
  PIN m_wbs_dat_o_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.680 204.000 186.280 ;
    END
  END m_wbs_dat_o_1[18]
  PIN m_wbs_dat_o_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 192.480 204.000 193.080 ;
    END
  END m_wbs_dat_o_1[19]
  PIN m_wbs_dat_o_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 76.200 204.000 76.800 ;
    END
  END m_wbs_dat_o_1[1]
  PIN m_wbs_dat_o_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 198.600 204.000 199.200 ;
    END
  END m_wbs_dat_o_1[20]
  PIN m_wbs_dat_o_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 205.400 204.000 206.000 ;
    END
  END m_wbs_dat_o_1[21]
  PIN m_wbs_dat_o_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 211.520 204.000 212.120 ;
    END
  END m_wbs_dat_o_1[22]
  PIN m_wbs_dat_o_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 218.320 204.000 218.920 ;
    END
  END m_wbs_dat_o_1[23]
  PIN m_wbs_dat_o_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 224.440 204.000 225.040 ;
    END
  END m_wbs_dat_o_1[24]
  PIN m_wbs_dat_o_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 231.240 204.000 231.840 ;
    END
  END m_wbs_dat_o_1[25]
  PIN m_wbs_dat_o_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 237.360 204.000 237.960 ;
    END
  END m_wbs_dat_o_1[26]
  PIN m_wbs_dat_o_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.160 204.000 244.760 ;
    END
  END m_wbs_dat_o_1[27]
  PIN m_wbs_dat_o_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.960 204.000 251.560 ;
    END
  END m_wbs_dat_o_1[28]
  PIN m_wbs_dat_o_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 257.080 204.000 257.680 ;
    END
  END m_wbs_dat_o_1[29]
  PIN m_wbs_dat_o_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 82.320 204.000 82.920 ;
    END
  END m_wbs_dat_o_1[2]
  PIN m_wbs_dat_o_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 263.880 204.000 264.480 ;
    END
  END m_wbs_dat_o_1[30]
  PIN m_wbs_dat_o_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 270.000 204.000 270.600 ;
    END
  END m_wbs_dat_o_1[31]
  PIN m_wbs_dat_o_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.120 204.000 89.720 ;
    END
  END m_wbs_dat_o_1[3]
  PIN m_wbs_dat_o_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 204.000 95.840 ;
    END
  END m_wbs_dat_o_1[4]
  PIN m_wbs_dat_o_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 102.040 204.000 102.640 ;
    END
  END m_wbs_dat_o_1[5]
  PIN m_wbs_dat_o_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 108.160 204.000 108.760 ;
    END
  END m_wbs_dat_o_1[6]
  PIN m_wbs_dat_o_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.960 204.000 115.560 ;
    END
  END m_wbs_dat_o_1[7]
  PIN m_wbs_dat_o_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 121.080 204.000 121.680 ;
    END
  END m_wbs_dat_o_1[8]
  PIN m_wbs_dat_o_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 204.000 128.480 ;
    END
  END m_wbs_dat_o_1[9]
  PIN m_wbs_dat_o_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 276.800 204.000 277.400 ;
    END
  END m_wbs_dat_o_2[0]
  PIN m_wbs_dat_o_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 297.880 204.000 298.480 ;
    END
  END m_wbs_dat_o_2[10]
  PIN m_wbs_dat_o_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 300.600 204.000 301.200 ;
    END
  END m_wbs_dat_o_2[11]
  PIN m_wbs_dat_o_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 302.640 204.000 303.240 ;
    END
  END m_wbs_dat_o_2[12]
  PIN m_wbs_dat_o_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 304.680 204.000 305.280 ;
    END
  END m_wbs_dat_o_2[13]
  PIN m_wbs_dat_o_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 306.720 204.000 307.320 ;
    END
  END m_wbs_dat_o_2[14]
  PIN m_wbs_dat_o_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 308.760 204.000 309.360 ;
    END
  END m_wbs_dat_o_2[15]
  PIN m_wbs_dat_o_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 310.800 204.000 311.400 ;
    END
  END m_wbs_dat_o_2[16]
  PIN m_wbs_dat_o_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 313.520 204.000 314.120 ;
    END
  END m_wbs_dat_o_2[17]
  PIN m_wbs_dat_o_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 315.560 204.000 316.160 ;
    END
  END m_wbs_dat_o_2[18]
  PIN m_wbs_dat_o_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 317.600 204.000 318.200 ;
    END
  END m_wbs_dat_o_2[19]
  PIN m_wbs_dat_o_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 278.840 204.000 279.440 ;
    END
  END m_wbs_dat_o_2[1]
  PIN m_wbs_dat_o_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 319.640 204.000 320.240 ;
    END
  END m_wbs_dat_o_2[20]
  PIN m_wbs_dat_o_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 321.680 204.000 322.280 ;
    END
  END m_wbs_dat_o_2[21]
  PIN m_wbs_dat_o_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 323.720 204.000 324.320 ;
    END
  END m_wbs_dat_o_2[22]
  PIN m_wbs_dat_o_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 326.440 204.000 327.040 ;
    END
  END m_wbs_dat_o_2[23]
  PIN m_wbs_dat_o_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 328.480 204.000 329.080 ;
    END
  END m_wbs_dat_o_2[24]
  PIN m_wbs_dat_o_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 330.520 204.000 331.120 ;
    END
  END m_wbs_dat_o_2[25]
  PIN m_wbs_dat_o_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 332.560 204.000 333.160 ;
    END
  END m_wbs_dat_o_2[26]
  PIN m_wbs_dat_o_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 334.600 204.000 335.200 ;
    END
  END m_wbs_dat_o_2[27]
  PIN m_wbs_dat_o_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 336.640 204.000 337.240 ;
    END
  END m_wbs_dat_o_2[28]
  PIN m_wbs_dat_o_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 339.360 204.000 339.960 ;
    END
  END m_wbs_dat_o_2[29]
  PIN m_wbs_dat_o_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 280.880 204.000 281.480 ;
    END
  END m_wbs_dat_o_2[2]
  PIN m_wbs_dat_o_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 341.400 204.000 342.000 ;
    END
  END m_wbs_dat_o_2[30]
  PIN m_wbs_dat_o_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 343.440 204.000 344.040 ;
    END
  END m_wbs_dat_o_2[31]
  PIN m_wbs_dat_o_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.920 204.000 283.520 ;
    END
  END m_wbs_dat_o_2[3]
  PIN m_wbs_dat_o_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 284.960 204.000 285.560 ;
    END
  END m_wbs_dat_o_2[4]
  PIN m_wbs_dat_o_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 287.000 204.000 287.600 ;
    END
  END m_wbs_dat_o_2[5]
  PIN m_wbs_dat_o_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 289.720 204.000 290.320 ;
    END
  END m_wbs_dat_o_2[6]
  PIN m_wbs_dat_o_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.760 204.000 292.360 ;
    END
  END m_wbs_dat_o_2[7]
  PIN m_wbs_dat_o_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 293.800 204.000 294.400 ;
    END
  END m_wbs_dat_o_2[8]
  PIN m_wbs_dat_o_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 295.840 204.000 296.440 ;
    END
  END m_wbs_dat_o_2[9]
  PIN m_wbs_dat_o_3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 345.480 204.000 346.080 ;
    END
  END m_wbs_dat_o_3[0]
  PIN m_wbs_dat_o_3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 367.240 204.000 367.840 ;
    END
  END m_wbs_dat_o_3[10]
  PIN m_wbs_dat_o_3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 369.280 204.000 369.880 ;
    END
  END m_wbs_dat_o_3[11]
  PIN m_wbs_dat_o_3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 371.320 204.000 371.920 ;
    END
  END m_wbs_dat_o_3[12]
  PIN m_wbs_dat_o_3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 373.360 204.000 373.960 ;
    END
  END m_wbs_dat_o_3[13]
  PIN m_wbs_dat_o_3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 376.080 204.000 376.680 ;
    END
  END m_wbs_dat_o_3[14]
  PIN m_wbs_dat_o_3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 378.120 204.000 378.720 ;
    END
  END m_wbs_dat_o_3[15]
  PIN m_wbs_dat_o_3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 380.160 204.000 380.760 ;
    END
  END m_wbs_dat_o_3[16]
  PIN m_wbs_dat_o_3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 382.200 204.000 382.800 ;
    END
  END m_wbs_dat_o_3[17]
  PIN m_wbs_dat_o_3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 384.240 204.000 384.840 ;
    END
  END m_wbs_dat_o_3[18]
  PIN m_wbs_dat_o_3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 386.280 204.000 386.880 ;
    END
  END m_wbs_dat_o_3[19]
  PIN m_wbs_dat_o_3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 347.520 204.000 348.120 ;
    END
  END m_wbs_dat_o_3[1]
  PIN m_wbs_dat_o_3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 389.000 204.000 389.600 ;
    END
  END m_wbs_dat_o_3[20]
  PIN m_wbs_dat_o_3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 391.040 204.000 391.640 ;
    END
  END m_wbs_dat_o_3[21]
  PIN m_wbs_dat_o_3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 393.080 204.000 393.680 ;
    END
  END m_wbs_dat_o_3[22]
  PIN m_wbs_dat_o_3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 395.120 204.000 395.720 ;
    END
  END m_wbs_dat_o_3[23]
  PIN m_wbs_dat_o_3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 397.160 204.000 397.760 ;
    END
  END m_wbs_dat_o_3[24]
  PIN m_wbs_dat_o_3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 399.200 204.000 399.800 ;
    END
  END m_wbs_dat_o_3[25]
  PIN m_wbs_dat_o_3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 401.920 204.000 402.520 ;
    END
  END m_wbs_dat_o_3[26]
  PIN m_wbs_dat_o_3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 403.960 204.000 404.560 ;
    END
  END m_wbs_dat_o_3[27]
  PIN m_wbs_dat_o_3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 406.000 204.000 406.600 ;
    END
  END m_wbs_dat_o_3[28]
  PIN m_wbs_dat_o_3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 408.040 204.000 408.640 ;
    END
  END m_wbs_dat_o_3[29]
  PIN m_wbs_dat_o_3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 349.560 204.000 350.160 ;
    END
  END m_wbs_dat_o_3[2]
  PIN m_wbs_dat_o_3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 410.080 204.000 410.680 ;
    END
  END m_wbs_dat_o_3[30]
  PIN m_wbs_dat_o_3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 412.120 204.000 412.720 ;
    END
  END m_wbs_dat_o_3[31]
  PIN m_wbs_dat_o_3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 352.280 204.000 352.880 ;
    END
  END m_wbs_dat_o_3[3]
  PIN m_wbs_dat_o_3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 354.320 204.000 354.920 ;
    END
  END m_wbs_dat_o_3[4]
  PIN m_wbs_dat_o_3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 356.360 204.000 356.960 ;
    END
  END m_wbs_dat_o_3[5]
  PIN m_wbs_dat_o_3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 358.400 204.000 359.000 ;
    END
  END m_wbs_dat_o_3[6]
  PIN m_wbs_dat_o_3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 360.440 204.000 361.040 ;
    END
  END m_wbs_dat_o_3[7]
  PIN m_wbs_dat_o_3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 363.160 204.000 363.760 ;
    END
  END m_wbs_dat_o_3[8]
  PIN m_wbs_dat_o_3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 365.200 204.000 365.800 ;
    END
  END m_wbs_dat_o_3[9]
  PIN m_wbs_dat_o_4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 414.840 204.000 415.440 ;
    END
  END m_wbs_dat_o_4[0]
  PIN m_wbs_dat_o_4[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 435.920 204.000 436.520 ;
    END
  END m_wbs_dat_o_4[10]
  PIN m_wbs_dat_o_4[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 438.640 204.000 439.240 ;
    END
  END m_wbs_dat_o_4[11]
  PIN m_wbs_dat_o_4[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 440.680 204.000 441.280 ;
    END
  END m_wbs_dat_o_4[12]
  PIN m_wbs_dat_o_4[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 442.720 204.000 443.320 ;
    END
  END m_wbs_dat_o_4[13]
  PIN m_wbs_dat_o_4[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 444.760 204.000 445.360 ;
    END
  END m_wbs_dat_o_4[14]
  PIN m_wbs_dat_o_4[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 446.800 204.000 447.400 ;
    END
  END m_wbs_dat_o_4[15]
  PIN m_wbs_dat_o_4[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 448.840 204.000 449.440 ;
    END
  END m_wbs_dat_o_4[16]
  PIN m_wbs_dat_o_4[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 451.560 204.000 452.160 ;
    END
  END m_wbs_dat_o_4[17]
  PIN m_wbs_dat_o_4[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 453.600 204.000 454.200 ;
    END
  END m_wbs_dat_o_4[18]
  PIN m_wbs_dat_o_4[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 455.640 204.000 456.240 ;
    END
  END m_wbs_dat_o_4[19]
  PIN m_wbs_dat_o_4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 416.880 204.000 417.480 ;
    END
  END m_wbs_dat_o_4[1]
  PIN m_wbs_dat_o_4[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 457.680 204.000 458.280 ;
    END
  END m_wbs_dat_o_4[20]
  PIN m_wbs_dat_o_4[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 459.720 204.000 460.320 ;
    END
  END m_wbs_dat_o_4[21]
  PIN m_wbs_dat_o_4[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 461.760 204.000 462.360 ;
    END
  END m_wbs_dat_o_4[22]
  PIN m_wbs_dat_o_4[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 464.480 204.000 465.080 ;
    END
  END m_wbs_dat_o_4[23]
  PIN m_wbs_dat_o_4[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 466.520 204.000 467.120 ;
    END
  END m_wbs_dat_o_4[24]
  PIN m_wbs_dat_o_4[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 468.560 204.000 469.160 ;
    END
  END m_wbs_dat_o_4[25]
  PIN m_wbs_dat_o_4[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 470.600 204.000 471.200 ;
    END
  END m_wbs_dat_o_4[26]
  PIN m_wbs_dat_o_4[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 472.640 204.000 473.240 ;
    END
  END m_wbs_dat_o_4[27]
  PIN m_wbs_dat_o_4[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 474.680 204.000 475.280 ;
    END
  END m_wbs_dat_o_4[28]
  PIN m_wbs_dat_o_4[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 477.400 204.000 478.000 ;
    END
  END m_wbs_dat_o_4[29]
  PIN m_wbs_dat_o_4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 418.920 204.000 419.520 ;
    END
  END m_wbs_dat_o_4[2]
  PIN m_wbs_dat_o_4[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 479.440 204.000 480.040 ;
    END
  END m_wbs_dat_o_4[30]
  PIN m_wbs_dat_o_4[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 481.480 204.000 482.080 ;
    END
  END m_wbs_dat_o_4[31]
  PIN m_wbs_dat_o_4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 420.960 204.000 421.560 ;
    END
  END m_wbs_dat_o_4[3]
  PIN m_wbs_dat_o_4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 423.000 204.000 423.600 ;
    END
  END m_wbs_dat_o_4[4]
  PIN m_wbs_dat_o_4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 425.720 204.000 426.320 ;
    END
  END m_wbs_dat_o_4[5]
  PIN m_wbs_dat_o_4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 427.760 204.000 428.360 ;
    END
  END m_wbs_dat_o_4[6]
  PIN m_wbs_dat_o_4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 429.800 204.000 430.400 ;
    END
  END m_wbs_dat_o_4[7]
  PIN m_wbs_dat_o_4[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 431.840 204.000 432.440 ;
    END
  END m_wbs_dat_o_4[8]
  PIN m_wbs_dat_o_4[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 433.880 204.000 434.480 ;
    END
  END m_wbs_dat_o_4[9]
  PIN m_wbs_dat_o_5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 483.520 204.000 484.120 ;
    END
  END m_wbs_dat_o_5[0]
  PIN m_wbs_dat_o_5[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 505.280 204.000 505.880 ;
    END
  END m_wbs_dat_o_5[10]
  PIN m_wbs_dat_o_5[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 507.320 204.000 507.920 ;
    END
  END m_wbs_dat_o_5[11]
  PIN m_wbs_dat_o_5[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 509.360 204.000 509.960 ;
    END
  END m_wbs_dat_o_5[12]
  PIN m_wbs_dat_o_5[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 511.400 204.000 512.000 ;
    END
  END m_wbs_dat_o_5[13]
  PIN m_wbs_dat_o_5[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 514.120 204.000 514.720 ;
    END
  END m_wbs_dat_o_5[14]
  PIN m_wbs_dat_o_5[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 516.160 204.000 516.760 ;
    END
  END m_wbs_dat_o_5[15]
  PIN m_wbs_dat_o_5[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 518.200 204.000 518.800 ;
    END
  END m_wbs_dat_o_5[16]
  PIN m_wbs_dat_o_5[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 520.240 204.000 520.840 ;
    END
  END m_wbs_dat_o_5[17]
  PIN m_wbs_dat_o_5[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 522.280 204.000 522.880 ;
    END
  END m_wbs_dat_o_5[18]
  PIN m_wbs_dat_o_5[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 524.320 204.000 524.920 ;
    END
  END m_wbs_dat_o_5[19]
  PIN m_wbs_dat_o_5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 485.560 204.000 486.160 ;
    END
  END m_wbs_dat_o_5[1]
  PIN m_wbs_dat_o_5[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 527.040 204.000 527.640 ;
    END
  END m_wbs_dat_o_5[20]
  PIN m_wbs_dat_o_5[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 529.080 204.000 529.680 ;
    END
  END m_wbs_dat_o_5[21]
  PIN m_wbs_dat_o_5[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 531.120 204.000 531.720 ;
    END
  END m_wbs_dat_o_5[22]
  PIN m_wbs_dat_o_5[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 533.160 204.000 533.760 ;
    END
  END m_wbs_dat_o_5[23]
  PIN m_wbs_dat_o_5[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.200 204.000 535.800 ;
    END
  END m_wbs_dat_o_5[24]
  PIN m_wbs_dat_o_5[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 537.240 204.000 537.840 ;
    END
  END m_wbs_dat_o_5[25]
  PIN m_wbs_dat_o_5[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 539.960 204.000 540.560 ;
    END
  END m_wbs_dat_o_5[26]
  PIN m_wbs_dat_o_5[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 542.000 204.000 542.600 ;
    END
  END m_wbs_dat_o_5[27]
  PIN m_wbs_dat_o_5[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 544.040 204.000 544.640 ;
    END
  END m_wbs_dat_o_5[28]
  PIN m_wbs_dat_o_5[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 546.080 204.000 546.680 ;
    END
  END m_wbs_dat_o_5[29]
  PIN m_wbs_dat_o_5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 488.280 204.000 488.880 ;
    END
  END m_wbs_dat_o_5[2]
  PIN m_wbs_dat_o_5[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 548.120 204.000 548.720 ;
    END
  END m_wbs_dat_o_5[30]
  PIN m_wbs_dat_o_5[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 550.840 204.000 551.440 ;
    END
  END m_wbs_dat_o_5[31]
  PIN m_wbs_dat_o_5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 490.320 204.000 490.920 ;
    END
  END m_wbs_dat_o_5[3]
  PIN m_wbs_dat_o_5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 492.360 204.000 492.960 ;
    END
  END m_wbs_dat_o_5[4]
  PIN m_wbs_dat_o_5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 494.400 204.000 495.000 ;
    END
  END m_wbs_dat_o_5[5]
  PIN m_wbs_dat_o_5[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 496.440 204.000 497.040 ;
    END
  END m_wbs_dat_o_5[6]
  PIN m_wbs_dat_o_5[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 498.480 204.000 499.080 ;
    END
  END m_wbs_dat_o_5[7]
  PIN m_wbs_dat_o_5[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 501.200 204.000 501.800 ;
    END
  END m_wbs_dat_o_5[8]
  PIN m_wbs_dat_o_5[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 503.240 204.000 503.840 ;
    END
  END m_wbs_dat_o_5[9]
  PIN m_wbs_dat_o_6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2.080 4.000 2.680 ;
    END
  END m_wbs_dat_o_6[0]
  PIN m_wbs_dat_o_6[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 42.880 4.000 43.480 ;
    END
  END m_wbs_dat_o_6[10]
  PIN m_wbs_dat_o_6[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 46.960 4.000 47.560 ;
    END
  END m_wbs_dat_o_6[11]
  PIN m_wbs_dat_o_6[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 51.040 4.000 51.640 ;
    END
  END m_wbs_dat_o_6[12]
  PIN m_wbs_dat_o_6[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 55.800 4.000 56.400 ;
    END
  END m_wbs_dat_o_6[13]
  PIN m_wbs_dat_o_6[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 59.880 4.000 60.480 ;
    END
  END m_wbs_dat_o_6[14]
  PIN m_wbs_dat_o_6[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 63.960 4.000 64.560 ;
    END
  END m_wbs_dat_o_6[15]
  PIN m_wbs_dat_o_6[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.040 4.000 68.640 ;
    END
  END m_wbs_dat_o_6[16]
  PIN m_wbs_dat_o_6[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.120 4.000 72.720 ;
    END
  END m_wbs_dat_o_6[17]
  PIN m_wbs_dat_o_6[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.200 4.000 76.800 ;
    END
  END m_wbs_dat_o_6[18]
  PIN m_wbs_dat_o_6[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.280 4.000 80.880 ;
    END
  END m_wbs_dat_o_6[19]
  PIN m_wbs_dat_o_6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.160 4.000 6.760 ;
    END
  END m_wbs_dat_o_6[1]
  PIN m_wbs_dat_o_6[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.360 4.000 84.960 ;
    END
  END m_wbs_dat_o_6[20]
  PIN m_wbs_dat_o_6[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.440 4.000 89.040 ;
    END
  END m_wbs_dat_o_6[21]
  PIN m_wbs_dat_o_6[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.520 4.000 93.120 ;
    END
  END m_wbs_dat_o_6[22]
  PIN m_wbs_dat_o_6[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.600 4.000 97.200 ;
    END
  END m_wbs_dat_o_6[23]
  PIN m_wbs_dat_o_6[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.680 4.000 101.280 ;
    END
  END m_wbs_dat_o_6[24]
  PIN m_wbs_dat_o_6[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 105.440 4.000 106.040 ;
    END
  END m_wbs_dat_o_6[25]
  PIN m_wbs_dat_o_6[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 109.520 4.000 110.120 ;
    END
  END m_wbs_dat_o_6[26]
  PIN m_wbs_dat_o_6[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 113.600 4.000 114.200 ;
    END
  END m_wbs_dat_o_6[27]
  PIN m_wbs_dat_o_6[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 117.680 4.000 118.280 ;
    END
  END m_wbs_dat_o_6[28]
  PIN m_wbs_dat_o_6[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 121.760 4.000 122.360 ;
    END
  END m_wbs_dat_o_6[29]
  PIN m_wbs_dat_o_6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.240 4.000 10.840 ;
    END
  END m_wbs_dat_o_6[2]
  PIN m_wbs_dat_o_6[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 125.840 4.000 126.440 ;
    END
  END m_wbs_dat_o_6[30]
  PIN m_wbs_dat_o_6[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 129.920 4.000 130.520 ;
    END
  END m_wbs_dat_o_6[31]
  PIN m_wbs_dat_o_6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 14.320 4.000 14.920 ;
    END
  END m_wbs_dat_o_6[3]
  PIN m_wbs_dat_o_6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 18.400 4.000 19.000 ;
    END
  END m_wbs_dat_o_6[4]
  PIN m_wbs_dat_o_6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 22.480 4.000 23.080 ;
    END
  END m_wbs_dat_o_6[5]
  PIN m_wbs_dat_o_6[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 26.560 4.000 27.160 ;
    END
  END m_wbs_dat_o_6[6]
  PIN m_wbs_dat_o_6[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 30.640 4.000 31.240 ;
    END
  END m_wbs_dat_o_6[7]
  PIN m_wbs_dat_o_6[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 34.720 4.000 35.320 ;
    END
  END m_wbs_dat_o_6[8]
  PIN m_wbs_dat_o_6[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 38.800 4.000 39.400 ;
    END
  END m_wbs_dat_o_6[9]
  PIN m_wbs_dat_o_7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 134.000 4.000 134.600 ;
    END
  END m_wbs_dat_o_7[0]
  PIN m_wbs_dat_o_7[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 175.480 4.000 176.080 ;
    END
  END m_wbs_dat_o_7[10]
  PIN m_wbs_dat_o_7[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 179.560 4.000 180.160 ;
    END
  END m_wbs_dat_o_7[11]
  PIN m_wbs_dat_o_7[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 183.640 4.000 184.240 ;
    END
  END m_wbs_dat_o_7[12]
  PIN m_wbs_dat_o_7[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 187.720 4.000 188.320 ;
    END
  END m_wbs_dat_o_7[13]
  PIN m_wbs_dat_o_7[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 191.800 4.000 192.400 ;
    END
  END m_wbs_dat_o_7[14]
  PIN m_wbs_dat_o_7[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 195.880 4.000 196.480 ;
    END
  END m_wbs_dat_o_7[15]
  PIN m_wbs_dat_o_7[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 199.960 4.000 200.560 ;
    END
  END m_wbs_dat_o_7[16]
  PIN m_wbs_dat_o_7[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.720 4.000 205.320 ;
    END
  END m_wbs_dat_o_7[17]
  PIN m_wbs_dat_o_7[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.800 4.000 209.400 ;
    END
  END m_wbs_dat_o_7[18]
  PIN m_wbs_dat_o_7[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.880 4.000 213.480 ;
    END
  END m_wbs_dat_o_7[19]
  PIN m_wbs_dat_o_7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 138.080 4.000 138.680 ;
    END
  END m_wbs_dat_o_7[1]
  PIN m_wbs_dat_o_7[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.960 4.000 217.560 ;
    END
  END m_wbs_dat_o_7[20]
  PIN m_wbs_dat_o_7[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 221.040 4.000 221.640 ;
    END
  END m_wbs_dat_o_7[21]
  PIN m_wbs_dat_o_7[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 225.120 4.000 225.720 ;
    END
  END m_wbs_dat_o_7[22]
  PIN m_wbs_dat_o_7[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 229.200 4.000 229.800 ;
    END
  END m_wbs_dat_o_7[23]
  PIN m_wbs_dat_o_7[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 233.280 4.000 233.880 ;
    END
  END m_wbs_dat_o_7[24]
  PIN m_wbs_dat_o_7[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 237.360 4.000 237.960 ;
    END
  END m_wbs_dat_o_7[25]
  PIN m_wbs_dat_o_7[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 241.440 4.000 242.040 ;
    END
  END m_wbs_dat_o_7[26]
  PIN m_wbs_dat_o_7[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 245.520 4.000 246.120 ;
    END
  END m_wbs_dat_o_7[27]
  PIN m_wbs_dat_o_7[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 249.600 4.000 250.200 ;
    END
  END m_wbs_dat_o_7[28]
  PIN m_wbs_dat_o_7[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 254.360 4.000 254.960 ;
    END
  END m_wbs_dat_o_7[29]
  PIN m_wbs_dat_o_7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 142.160 4.000 142.760 ;
    END
  END m_wbs_dat_o_7[2]
  PIN m_wbs_dat_o_7[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 258.440 4.000 259.040 ;
    END
  END m_wbs_dat_o_7[30]
  PIN m_wbs_dat_o_7[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 262.520 4.000 263.120 ;
    END
  END m_wbs_dat_o_7[31]
  PIN m_wbs_dat_o_7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 146.240 4.000 146.840 ;
    END
  END m_wbs_dat_o_7[3]
  PIN m_wbs_dat_o_7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 150.320 4.000 150.920 ;
    END
  END m_wbs_dat_o_7[4]
  PIN m_wbs_dat_o_7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 155.080 4.000 155.680 ;
    END
  END m_wbs_dat_o_7[5]
  PIN m_wbs_dat_o_7[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 159.160 4.000 159.760 ;
    END
  END m_wbs_dat_o_7[6]
  PIN m_wbs_dat_o_7[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 163.240 4.000 163.840 ;
    END
  END m_wbs_dat_o_7[7]
  PIN m_wbs_dat_o_7[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 167.320 4.000 167.920 ;
    END
  END m_wbs_dat_o_7[8]
  PIN m_wbs_dat_o_7[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 171.400 4.000 172.000 ;
    END
  END m_wbs_dat_o_7[9]
  PIN m_wbs_dat_o_8[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 266.600 4.000 267.200 ;
    END
  END m_wbs_dat_o_8[0]
  PIN m_wbs_dat_o_8[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 308.080 4.000 308.680 ;
    END
  END m_wbs_dat_o_8[10]
  PIN m_wbs_dat_o_8[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.160 4.000 312.760 ;
    END
  END m_wbs_dat_o_8[11]
  PIN m_wbs_dat_o_8[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 316.240 4.000 316.840 ;
    END
  END m_wbs_dat_o_8[12]
  PIN m_wbs_dat_o_8[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 320.320 4.000 320.920 ;
    END
  END m_wbs_dat_o_8[13]
  PIN m_wbs_dat_o_8[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 324.400 4.000 325.000 ;
    END
  END m_wbs_dat_o_8[14]
  PIN m_wbs_dat_o_8[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 328.480 4.000 329.080 ;
    END
  END m_wbs_dat_o_8[15]
  PIN m_wbs_dat_o_8[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 332.560 4.000 333.160 ;
    END
  END m_wbs_dat_o_8[16]
  PIN m_wbs_dat_o_8[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 336.640 4.000 337.240 ;
    END
  END m_wbs_dat_o_8[17]
  PIN m_wbs_dat_o_8[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 340.720 4.000 341.320 ;
    END
  END m_wbs_dat_o_8[18]
  PIN m_wbs_dat_o_8[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 344.800 4.000 345.400 ;
    END
  END m_wbs_dat_o_8[19]
  PIN m_wbs_dat_o_8[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 270.680 4.000 271.280 ;
    END
  END m_wbs_dat_o_8[1]
  PIN m_wbs_dat_o_8[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 348.880 4.000 349.480 ;
    END
  END m_wbs_dat_o_8[20]
  PIN m_wbs_dat_o_8[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 353.640 4.000 354.240 ;
    END
  END m_wbs_dat_o_8[21]
  PIN m_wbs_dat_o_8[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 357.720 4.000 358.320 ;
    END
  END m_wbs_dat_o_8[22]
  PIN m_wbs_dat_o_8[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 361.800 4.000 362.400 ;
    END
  END m_wbs_dat_o_8[23]
  PIN m_wbs_dat_o_8[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 365.880 4.000 366.480 ;
    END
  END m_wbs_dat_o_8[24]
  PIN m_wbs_dat_o_8[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 369.960 4.000 370.560 ;
    END
  END m_wbs_dat_o_8[25]
  PIN m_wbs_dat_o_8[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 374.040 4.000 374.640 ;
    END
  END m_wbs_dat_o_8[26]
  PIN m_wbs_dat_o_8[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 378.120 4.000 378.720 ;
    END
  END m_wbs_dat_o_8[27]
  PIN m_wbs_dat_o_8[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 382.200 4.000 382.800 ;
    END
  END m_wbs_dat_o_8[28]
  PIN m_wbs_dat_o_8[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 386.280 4.000 386.880 ;
    END
  END m_wbs_dat_o_8[29]
  PIN m_wbs_dat_o_8[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 274.760 4.000 275.360 ;
    END
  END m_wbs_dat_o_8[2]
  PIN m_wbs_dat_o_8[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 390.360 4.000 390.960 ;
    END
  END m_wbs_dat_o_8[30]
  PIN m_wbs_dat_o_8[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 394.440 4.000 395.040 ;
    END
  END m_wbs_dat_o_8[31]
  PIN m_wbs_dat_o_8[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 278.840 4.000 279.440 ;
    END
  END m_wbs_dat_o_8[3]
  PIN m_wbs_dat_o_8[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 282.920 4.000 283.520 ;
    END
  END m_wbs_dat_o_8[4]
  PIN m_wbs_dat_o_8[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 287.000 4.000 287.600 ;
    END
  END m_wbs_dat_o_8[5]
  PIN m_wbs_dat_o_8[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 291.080 4.000 291.680 ;
    END
  END m_wbs_dat_o_8[6]
  PIN m_wbs_dat_o_8[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 295.160 4.000 295.760 ;
    END
  END m_wbs_dat_o_8[7]
  PIN m_wbs_dat_o_8[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 299.240 4.000 299.840 ;
    END
  END m_wbs_dat_o_8[8]
  PIN m_wbs_dat_o_8[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.000 4.000 304.600 ;
    END
  END m_wbs_dat_o_8[9]
  PIN m_wbs_dat_o_9[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 398.520 4.000 399.120 ;
    END
  END m_wbs_dat_o_9[0]
  PIN m_wbs_dat_o_9[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 440.000 4.000 440.600 ;
    END
  END m_wbs_dat_o_9[10]
  PIN m_wbs_dat_o_9[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.080 4.000 444.680 ;
    END
  END m_wbs_dat_o_9[11]
  PIN m_wbs_dat_o_9[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 448.160 4.000 448.760 ;
    END
  END m_wbs_dat_o_9[12]
  PIN m_wbs_dat_o_9[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 452.920 4.000 453.520 ;
    END
  END m_wbs_dat_o_9[13]
  PIN m_wbs_dat_o_9[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 457.000 4.000 457.600 ;
    END
  END m_wbs_dat_o_9[14]
  PIN m_wbs_dat_o_9[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 461.080 4.000 461.680 ;
    END
  END m_wbs_dat_o_9[15]
  PIN m_wbs_dat_o_9[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 465.160 4.000 465.760 ;
    END
  END m_wbs_dat_o_9[16]
  PIN m_wbs_dat_o_9[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 469.240 4.000 469.840 ;
    END
  END m_wbs_dat_o_9[17]
  PIN m_wbs_dat_o_9[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 473.320 4.000 473.920 ;
    END
  END m_wbs_dat_o_9[18]
  PIN m_wbs_dat_o_9[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 477.400 4.000 478.000 ;
    END
  END m_wbs_dat_o_9[19]
  PIN m_wbs_dat_o_9[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 403.280 4.000 403.880 ;
    END
  END m_wbs_dat_o_9[1]
  PIN m_wbs_dat_o_9[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 481.480 4.000 482.080 ;
    END
  END m_wbs_dat_o_9[20]
  PIN m_wbs_dat_o_9[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 485.560 4.000 486.160 ;
    END
  END m_wbs_dat_o_9[21]
  PIN m_wbs_dat_o_9[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 489.640 4.000 490.240 ;
    END
  END m_wbs_dat_o_9[22]
  PIN m_wbs_dat_o_9[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 493.720 4.000 494.320 ;
    END
  END m_wbs_dat_o_9[23]
  PIN m_wbs_dat_o_9[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 497.800 4.000 498.400 ;
    END
  END m_wbs_dat_o_9[24]
  PIN m_wbs_dat_o_9[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 502.560 4.000 503.160 ;
    END
  END m_wbs_dat_o_9[25]
  PIN m_wbs_dat_o_9[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 506.640 4.000 507.240 ;
    END
  END m_wbs_dat_o_9[26]
  PIN m_wbs_dat_o_9[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 510.720 4.000 511.320 ;
    END
  END m_wbs_dat_o_9[27]
  PIN m_wbs_dat_o_9[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 514.800 4.000 515.400 ;
    END
  END m_wbs_dat_o_9[28]
  PIN m_wbs_dat_o_9[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 518.880 4.000 519.480 ;
    END
  END m_wbs_dat_o_9[29]
  PIN m_wbs_dat_o_9[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 407.360 4.000 407.960 ;
    END
  END m_wbs_dat_o_9[2]
  PIN m_wbs_dat_o_9[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 522.960 4.000 523.560 ;
    END
  END m_wbs_dat_o_9[30]
  PIN m_wbs_dat_o_9[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 527.040 4.000 527.640 ;
    END
  END m_wbs_dat_o_9[31]
  PIN m_wbs_dat_o_9[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 411.440 4.000 412.040 ;
    END
  END m_wbs_dat_o_9[3]
  PIN m_wbs_dat_o_9[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 415.520 4.000 416.120 ;
    END
  END m_wbs_dat_o_9[4]
  PIN m_wbs_dat_o_9[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 419.600 4.000 420.200 ;
    END
  END m_wbs_dat_o_9[5]
  PIN m_wbs_dat_o_9[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 423.680 4.000 424.280 ;
    END
  END m_wbs_dat_o_9[6]
  PIN m_wbs_dat_o_9[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 427.760 4.000 428.360 ;
    END
  END m_wbs_dat_o_9[7]
  PIN m_wbs_dat_o_9[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 431.840 4.000 432.440 ;
    END
  END m_wbs_dat_o_9[8]
  PIN m_wbs_dat_o_9[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 435.920 4.000 436.520 ;
    END
  END m_wbs_dat_o_9[9]
  PIN m_wbs_we_i
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 596.000 183.910 604.000 ;
    END
  END m_wbs_we_i
  PIN mt_QEI_ChA_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 596.000 129.630 604.000 ;
    END
  END mt_QEI_ChA_0
  PIN mt_QEI_ChA_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 596.000 131.010 604.000 ;
    END
  END mt_QEI_ChA_1
  PIN mt_QEI_ChA_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 596.000 131.930 604.000 ;
    END
  END mt_QEI_ChA_2
  PIN mt_QEI_ChA_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 596.000 132.850 604.000 ;
    END
  END mt_QEI_ChA_3
  PIN mt_QEI_ChB_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 596.000 134.230 604.000 ;
    END
  END mt_QEI_ChB_0
  PIN mt_QEI_ChB_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 596.000 135.150 604.000 ;
    END
  END mt_QEI_ChB_1
  PIN mt_QEI_ChB_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 596.000 136.070 604.000 ;
    END
  END mt_QEI_ChB_2
  PIN mt_QEI_ChB_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 596.000 136.990 604.000 ;
    END
  END mt_QEI_ChB_3
  PIN mt_clo_test
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 596.000 138.370 604.000 ;
    END
  END mt_clo_test
  PIN mt_pwm_h_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 596.000 139.290 604.000 ;
    END
  END mt_pwm_h_0
  PIN mt_pwm_h_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 596.000 140.210 604.000 ;
    END
  END mt_pwm_h_1
  PIN mt_pwm_h_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 596.000 141.590 604.000 ;
    END
  END mt_pwm_h_2
  PIN mt_pwm_h_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 596.000 142.510 604.000 ;
    END
  END mt_pwm_h_3
  PIN mt_pwm_l_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 596.000 143.430 604.000 ;
    END
  END mt_pwm_l_0
  PIN mt_pwm_l_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 596.000 144.810 604.000 ;
    END
  END mt_pwm_l_1
  PIN mt_pwm_l_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 596.000 145.730 604.000 ;
    END
  END mt_pwm_l_2
  PIN mt_pwm_l_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 596.000 146.650 604.000 ;
    END
  END mt_pwm_l_3
  PIN mt_pwm_test
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 596.000 147.570 604.000 ;
    END
  END mt_pwm_test
  PIN mt_sync_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 604.000 ;
    END
  END mt_sync_in[0]
  PIN mt_sync_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 596.000 150.790 604.000 ;
    END
  END mt_sync_in[1]
  PIN mt_sync_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 596.000 152.170 604.000 ;
    END
  END mt_sync_in[2]
  PIN mt_sync_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 596.000 153.090 604.000 ;
    END
  END mt_sync_in[3]
  PIN mt_sync_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 596.000 154.010 604.000 ;
    END
  END mt_sync_in[4]
  PIN mt_sync_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 596.000 155.390 604.000 ;
    END
  END mt_sync_in[5]
  PIN mt_sync_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 596.000 156.310 604.000 ;
    END
  END mt_sync_in[6]
  PIN mt_sync_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 596.000 157.230 604.000 ;
    END
  END mt_sync_in[7]
  PIN mt_sync_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 596.000 148.950 604.000 ;
    END
  END mt_sync_out
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 -4.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 -4.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 -4.000 7.730 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 -4.000 13.710 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 -4.000 63.390 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 -4.000 67.990 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 -4.000 72.130 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 -4.000 76.730 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 -4.000 80.870 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 -4.000 85.470 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 -4.000 89.610 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 -4.000 94.210 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 -4.000 98.350 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 -4.000 102.950 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 -4.000 19.690 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 -4.000 107.090 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 -4.000 111.690 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 -4.000 115.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 -4.000 120.430 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 -4.000 124.570 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 -4.000 129.170 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 -4.000 133.310 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 -4.000 137.910 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 -4.000 142.050 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 -4.000 146.650 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 -4.000 25.210 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 -4.000 151.250 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 -4.000 155.390 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 -4.000 31.190 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 -4.000 37.170 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 -4.000 41.310 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 -4.000 45.910 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 -4.000 50.050 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 -4.000 54.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 -4.000 59.250 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 -4.000 9.570 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 -4.000 15.090 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 -4.000 64.770 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 -4.000 69.370 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 -4.000 73.510 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 -4.000 78.110 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 -4.000 82.250 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 -4.000 86.850 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 -4.000 90.990 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 -4.000 95.590 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 -4.000 99.730 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 -4.000 104.330 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 -4.000 21.070 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 -4.000 108.470 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 -4.000 113.070 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 -4.000 117.670 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 -4.000 121.810 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 -4.000 126.410 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 -4.000 130.550 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 -4.000 135.150 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 -4.000 139.290 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 -4.000 143.890 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 -4.000 148.030 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 -4.000 27.050 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 -4.000 152.630 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 -4.000 156.770 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 -4.000 32.570 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 -4.000 38.550 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 -4.000 43.150 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 -4.000 47.290 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 -4.000 51.890 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 -4.000 56.030 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 -4.000 60.630 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 -4.000 16.470 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 -4.000 66.150 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 -4.000 70.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 -4.000 74.890 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 -4.000 79.490 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 -4.000 83.630 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 -4.000 88.230 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 -4.000 92.830 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 -4.000 96.970 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 -4.000 101.570 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 -4.000 105.710 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 -4.000 22.450 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 -4.000 110.310 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 -4.000 114.450 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 -4.000 119.050 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 -4.000 123.190 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 -4.000 127.790 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 -4.000 131.930 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 -4.000 136.530 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 -4.000 140.670 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 -4.000 145.270 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 -4.000 149.410 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 -4.000 28.430 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 -4.000 154.010 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 -4.000 158.150 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 -4.000 34.410 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 -4.000 39.930 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 -4.000 44.530 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 -4.000 48.670 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 -4.000 53.270 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 -4.000 57.410 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 -4.000 62.010 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 -4.000 18.310 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 -4.000 23.830 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 -4.000 29.810 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 -4.000 35.790 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 -4.000 10.950 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 -4.000 12.330 4.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.895 587.605 ;
      LAYER met1 ;
        RECT 0.530 7.180 199.570 589.860 ;
      LAYER met2 ;
        RECT 1.110 595.720 1.190 598.245 ;
        RECT 2.030 595.720 2.110 598.245 ;
        RECT 2.950 595.720 3.030 598.245 ;
        RECT 3.870 595.720 4.410 598.245 ;
        RECT 5.250 595.720 5.330 598.245 ;
        RECT 6.170 595.720 6.250 598.245 ;
        RECT 7.090 595.720 7.630 598.245 ;
        RECT 8.470 595.720 8.550 598.245 ;
        RECT 9.390 595.720 9.470 598.245 ;
        RECT 10.310 595.720 10.850 598.245 ;
        RECT 11.690 595.720 11.770 598.245 ;
        RECT 12.610 595.720 12.690 598.245 ;
        RECT 13.530 595.720 13.610 598.245 ;
        RECT 14.450 595.720 14.990 598.245 ;
        RECT 15.830 595.720 15.910 598.245 ;
        RECT 16.750 595.720 16.830 598.245 ;
        RECT 17.670 595.720 18.210 598.245 ;
        RECT 19.050 595.720 19.130 598.245 ;
        RECT 19.970 595.720 20.050 598.245 ;
        RECT 20.890 595.720 21.430 598.245 ;
        RECT 22.270 595.720 22.350 598.245 ;
        RECT 23.190 595.720 23.270 598.245 ;
        RECT 24.110 595.720 24.190 598.245 ;
        RECT 25.030 595.720 25.570 598.245 ;
        RECT 26.410 595.720 26.490 598.245 ;
        RECT 27.330 595.720 27.410 598.245 ;
        RECT 28.250 595.720 28.790 598.245 ;
        RECT 29.630 595.720 29.710 598.245 ;
        RECT 30.550 595.720 30.630 598.245 ;
        RECT 31.470 595.720 32.010 598.245 ;
        RECT 32.850 595.720 32.930 598.245 ;
        RECT 33.770 595.720 33.850 598.245 ;
        RECT 34.690 595.720 34.770 598.245 ;
        RECT 35.610 595.720 36.150 598.245 ;
        RECT 36.990 595.720 37.070 598.245 ;
        RECT 37.910 595.720 37.990 598.245 ;
        RECT 38.830 595.720 39.370 598.245 ;
        RECT 40.210 595.720 40.290 598.245 ;
        RECT 41.130 595.720 41.210 598.245 ;
        RECT 42.050 595.720 42.590 598.245 ;
        RECT 43.430 595.720 43.510 598.245 ;
        RECT 44.350 595.720 44.430 598.245 ;
        RECT 45.270 595.720 45.350 598.245 ;
        RECT 46.190 595.720 46.730 598.245 ;
        RECT 47.570 595.720 47.650 598.245 ;
        RECT 48.490 595.720 48.570 598.245 ;
        RECT 49.410 595.720 49.950 598.245 ;
        RECT 50.790 595.720 50.870 598.245 ;
        RECT 51.710 595.720 51.790 598.245 ;
        RECT 52.630 595.720 53.170 598.245 ;
        RECT 54.010 595.720 54.090 598.245 ;
        RECT 54.930 595.720 55.010 598.245 ;
        RECT 55.850 595.720 55.930 598.245 ;
        RECT 56.770 595.720 57.310 598.245 ;
        RECT 58.150 595.720 58.230 598.245 ;
        RECT 59.070 595.720 59.150 598.245 ;
        RECT 59.990 595.720 60.530 598.245 ;
        RECT 61.370 595.720 61.450 598.245 ;
        RECT 62.290 595.720 62.370 598.245 ;
        RECT 63.210 595.720 63.750 598.245 ;
        RECT 64.590 595.720 64.670 598.245 ;
        RECT 65.510 595.720 65.590 598.245 ;
        RECT 66.430 595.720 66.970 598.245 ;
        RECT 67.810 595.720 67.890 598.245 ;
        RECT 68.730 595.720 68.810 598.245 ;
        RECT 69.650 595.720 69.730 598.245 ;
        RECT 70.570 595.720 71.110 598.245 ;
        RECT 71.950 595.720 72.030 598.245 ;
        RECT 72.870 595.720 72.950 598.245 ;
        RECT 73.790 595.720 74.330 598.245 ;
        RECT 75.170 595.720 75.250 598.245 ;
        RECT 76.090 595.720 76.170 598.245 ;
        RECT 77.010 595.720 77.550 598.245 ;
        RECT 78.390 595.720 78.470 598.245 ;
        RECT 79.310 595.720 79.390 598.245 ;
        RECT 80.230 595.720 80.310 598.245 ;
        RECT 81.150 595.720 81.690 598.245 ;
        RECT 82.530 595.720 82.610 598.245 ;
        RECT 83.450 595.720 83.530 598.245 ;
        RECT 84.370 595.720 84.910 598.245 ;
        RECT 85.750 595.720 85.830 598.245 ;
        RECT 86.670 595.720 86.750 598.245 ;
        RECT 87.590 595.720 88.130 598.245 ;
        RECT 88.970 595.720 89.050 598.245 ;
        RECT 89.890 595.720 89.970 598.245 ;
        RECT 90.810 595.720 90.890 598.245 ;
        RECT 91.730 595.720 92.270 598.245 ;
        RECT 93.110 595.720 93.190 598.245 ;
        RECT 94.030 595.720 94.110 598.245 ;
        RECT 94.950 595.720 95.490 598.245 ;
        RECT 96.330 595.720 96.410 598.245 ;
        RECT 97.250 595.720 97.330 598.245 ;
        RECT 98.170 595.720 98.710 598.245 ;
        RECT 99.550 595.720 99.630 598.245 ;
        RECT 100.470 595.720 100.550 598.245 ;
        RECT 101.390 595.720 101.470 598.245 ;
        RECT 102.310 595.720 102.850 598.245 ;
        RECT 103.690 595.720 103.770 598.245 ;
        RECT 104.610 595.720 104.690 598.245 ;
        RECT 105.530 595.720 106.070 598.245 ;
        RECT 106.910 595.720 106.990 598.245 ;
        RECT 107.830 595.720 107.910 598.245 ;
        RECT 108.750 595.720 109.290 598.245 ;
        RECT 110.130 595.720 110.210 598.245 ;
        RECT 111.050 595.720 111.130 598.245 ;
        RECT 111.970 595.720 112.050 598.245 ;
        RECT 112.890 595.720 113.430 598.245 ;
        RECT 114.270 595.720 114.350 598.245 ;
        RECT 115.190 595.720 115.270 598.245 ;
        RECT 116.110 595.720 116.650 598.245 ;
        RECT 117.490 595.720 117.570 598.245 ;
        RECT 118.410 595.720 118.490 598.245 ;
        RECT 119.330 595.720 119.870 598.245 ;
        RECT 120.710 595.720 120.790 598.245 ;
        RECT 121.630 595.720 121.710 598.245 ;
        RECT 122.550 595.720 122.630 598.245 ;
        RECT 123.470 595.720 124.010 598.245 ;
        RECT 124.850 595.720 124.930 598.245 ;
        RECT 125.770 595.720 125.850 598.245 ;
        RECT 126.690 595.720 127.230 598.245 ;
        RECT 128.070 595.720 128.150 598.245 ;
        RECT 128.990 595.720 129.070 598.245 ;
        RECT 129.910 595.720 130.450 598.245 ;
        RECT 131.290 595.720 131.370 598.245 ;
        RECT 132.210 595.720 132.290 598.245 ;
        RECT 133.130 595.720 133.670 598.245 ;
        RECT 134.510 595.720 134.590 598.245 ;
        RECT 135.430 595.720 135.510 598.245 ;
        RECT 136.350 595.720 136.430 598.245 ;
        RECT 137.270 595.720 137.810 598.245 ;
        RECT 138.650 595.720 138.730 598.245 ;
        RECT 139.570 595.720 139.650 598.245 ;
        RECT 140.490 595.720 141.030 598.245 ;
        RECT 141.870 595.720 141.950 598.245 ;
        RECT 142.790 595.720 142.870 598.245 ;
        RECT 143.710 595.720 144.250 598.245 ;
        RECT 145.090 595.720 145.170 598.245 ;
        RECT 146.010 595.720 146.090 598.245 ;
        RECT 146.930 595.720 147.010 598.245 ;
        RECT 147.850 595.720 148.390 598.245 ;
        RECT 149.230 595.720 149.310 598.245 ;
        RECT 150.150 595.720 150.230 598.245 ;
        RECT 151.070 595.720 151.610 598.245 ;
        RECT 152.450 595.720 152.530 598.245 ;
        RECT 153.370 595.720 153.450 598.245 ;
        RECT 154.290 595.720 154.830 598.245 ;
        RECT 155.670 595.720 155.750 598.245 ;
        RECT 156.590 595.720 156.670 598.245 ;
        RECT 157.510 595.720 157.590 598.245 ;
        RECT 158.430 595.720 158.970 598.245 ;
        RECT 159.810 595.720 159.890 598.245 ;
        RECT 160.730 595.720 160.810 598.245 ;
        RECT 161.650 595.720 162.190 598.245 ;
        RECT 163.030 595.720 163.110 598.245 ;
        RECT 163.950 595.720 164.030 598.245 ;
        RECT 164.870 595.720 165.410 598.245 ;
        RECT 166.250 595.720 166.330 598.245 ;
        RECT 167.170 595.720 167.250 598.245 ;
        RECT 168.090 595.720 168.170 598.245 ;
        RECT 169.010 595.720 169.550 598.245 ;
        RECT 170.390 595.720 170.470 598.245 ;
        RECT 171.310 595.720 171.390 598.245 ;
        RECT 172.230 595.720 172.770 598.245 ;
        RECT 173.610 595.720 173.690 598.245 ;
        RECT 174.530 595.720 174.610 598.245 ;
        RECT 175.450 595.720 175.990 598.245 ;
        RECT 176.830 595.720 176.910 598.245 ;
        RECT 177.750 595.720 177.830 598.245 ;
        RECT 178.670 595.720 178.750 598.245 ;
        RECT 179.590 595.720 180.130 598.245 ;
        RECT 180.970 595.720 181.050 598.245 ;
        RECT 181.890 595.720 181.970 598.245 ;
        RECT 182.810 595.720 183.350 598.245 ;
        RECT 184.190 595.720 184.270 598.245 ;
        RECT 185.110 595.720 185.190 598.245 ;
        RECT 186.030 595.720 186.570 598.245 ;
        RECT 187.410 595.720 187.490 598.245 ;
        RECT 188.330 595.720 188.410 598.245 ;
        RECT 189.250 595.720 189.330 598.245 ;
        RECT 190.170 595.720 190.710 598.245 ;
        RECT 191.550 595.720 191.630 598.245 ;
        RECT 192.470 595.720 192.550 598.245 ;
        RECT 193.390 595.720 193.930 598.245 ;
        RECT 194.770 595.720 194.850 598.245 ;
        RECT 195.690 595.720 195.770 598.245 ;
        RECT 196.610 595.720 197.150 598.245 ;
        RECT 197.990 595.720 198.070 598.245 ;
        RECT 198.910 595.720 198.990 598.245 ;
        RECT 0.560 4.280 199.540 595.720 ;
        RECT 1.110 0.835 1.650 4.280 ;
        RECT 2.490 0.835 3.030 4.280 ;
        RECT 3.870 0.835 4.410 4.280 ;
        RECT 5.250 0.835 5.790 4.280 ;
        RECT 6.630 0.835 7.170 4.280 ;
        RECT 8.010 0.835 9.010 4.280 ;
        RECT 9.850 0.835 10.390 4.280 ;
        RECT 11.230 0.835 11.770 4.280 ;
        RECT 12.610 0.835 13.150 4.280 ;
        RECT 13.990 0.835 14.530 4.280 ;
        RECT 15.370 0.835 15.910 4.280 ;
        RECT 16.750 0.835 17.750 4.280 ;
        RECT 18.590 0.835 19.130 4.280 ;
        RECT 19.970 0.835 20.510 4.280 ;
        RECT 21.350 0.835 21.890 4.280 ;
        RECT 22.730 0.835 23.270 4.280 ;
        RECT 24.110 0.835 24.650 4.280 ;
        RECT 25.490 0.835 26.490 4.280 ;
        RECT 27.330 0.835 27.870 4.280 ;
        RECT 28.710 0.835 29.250 4.280 ;
        RECT 30.090 0.835 30.630 4.280 ;
        RECT 31.470 0.835 32.010 4.280 ;
        RECT 32.850 0.835 33.850 4.280 ;
        RECT 34.690 0.835 35.230 4.280 ;
        RECT 36.070 0.835 36.610 4.280 ;
        RECT 37.450 0.835 37.990 4.280 ;
        RECT 38.830 0.835 39.370 4.280 ;
        RECT 40.210 0.835 40.750 4.280 ;
        RECT 41.590 0.835 42.590 4.280 ;
        RECT 43.430 0.835 43.970 4.280 ;
        RECT 44.810 0.835 45.350 4.280 ;
        RECT 46.190 0.835 46.730 4.280 ;
        RECT 47.570 0.835 48.110 4.280 ;
        RECT 48.950 0.835 49.490 4.280 ;
        RECT 50.330 0.835 51.330 4.280 ;
        RECT 52.170 0.835 52.710 4.280 ;
        RECT 53.550 0.835 54.090 4.280 ;
        RECT 54.930 0.835 55.470 4.280 ;
        RECT 56.310 0.835 56.850 4.280 ;
        RECT 57.690 0.835 58.690 4.280 ;
        RECT 59.530 0.835 60.070 4.280 ;
        RECT 60.910 0.835 61.450 4.280 ;
        RECT 62.290 0.835 62.830 4.280 ;
        RECT 63.670 0.835 64.210 4.280 ;
        RECT 65.050 0.835 65.590 4.280 ;
        RECT 66.430 0.835 67.430 4.280 ;
        RECT 68.270 0.835 68.810 4.280 ;
        RECT 69.650 0.835 70.190 4.280 ;
        RECT 71.030 0.835 71.570 4.280 ;
        RECT 72.410 0.835 72.950 4.280 ;
        RECT 73.790 0.835 74.330 4.280 ;
        RECT 75.170 0.835 76.170 4.280 ;
        RECT 77.010 0.835 77.550 4.280 ;
        RECT 78.390 0.835 78.930 4.280 ;
        RECT 79.770 0.835 80.310 4.280 ;
        RECT 81.150 0.835 81.690 4.280 ;
        RECT 82.530 0.835 83.070 4.280 ;
        RECT 83.910 0.835 84.910 4.280 ;
        RECT 85.750 0.835 86.290 4.280 ;
        RECT 87.130 0.835 87.670 4.280 ;
        RECT 88.510 0.835 89.050 4.280 ;
        RECT 89.890 0.835 90.430 4.280 ;
        RECT 91.270 0.835 92.270 4.280 ;
        RECT 93.110 0.835 93.650 4.280 ;
        RECT 94.490 0.835 95.030 4.280 ;
        RECT 95.870 0.835 96.410 4.280 ;
        RECT 97.250 0.835 97.790 4.280 ;
        RECT 98.630 0.835 99.170 4.280 ;
        RECT 100.010 0.835 101.010 4.280 ;
        RECT 101.850 0.835 102.390 4.280 ;
        RECT 103.230 0.835 103.770 4.280 ;
        RECT 104.610 0.835 105.150 4.280 ;
        RECT 105.990 0.835 106.530 4.280 ;
        RECT 107.370 0.835 107.910 4.280 ;
        RECT 108.750 0.835 109.750 4.280 ;
        RECT 110.590 0.835 111.130 4.280 ;
        RECT 111.970 0.835 112.510 4.280 ;
        RECT 113.350 0.835 113.890 4.280 ;
        RECT 114.730 0.835 115.270 4.280 ;
        RECT 116.110 0.835 117.110 4.280 ;
        RECT 117.950 0.835 118.490 4.280 ;
        RECT 119.330 0.835 119.870 4.280 ;
        RECT 120.710 0.835 121.250 4.280 ;
        RECT 122.090 0.835 122.630 4.280 ;
        RECT 123.470 0.835 124.010 4.280 ;
        RECT 124.850 0.835 125.850 4.280 ;
        RECT 126.690 0.835 127.230 4.280 ;
        RECT 128.070 0.835 128.610 4.280 ;
        RECT 129.450 0.835 129.990 4.280 ;
        RECT 130.830 0.835 131.370 4.280 ;
        RECT 132.210 0.835 132.750 4.280 ;
        RECT 133.590 0.835 134.590 4.280 ;
        RECT 135.430 0.835 135.970 4.280 ;
        RECT 136.810 0.835 137.350 4.280 ;
        RECT 138.190 0.835 138.730 4.280 ;
        RECT 139.570 0.835 140.110 4.280 ;
        RECT 140.950 0.835 141.490 4.280 ;
        RECT 142.330 0.835 143.330 4.280 ;
        RECT 144.170 0.835 144.710 4.280 ;
        RECT 145.550 0.835 146.090 4.280 ;
        RECT 146.930 0.835 147.470 4.280 ;
        RECT 148.310 0.835 148.850 4.280 ;
        RECT 149.690 0.835 150.690 4.280 ;
        RECT 151.530 0.835 152.070 4.280 ;
        RECT 152.910 0.835 153.450 4.280 ;
        RECT 154.290 0.835 154.830 4.280 ;
        RECT 155.670 0.835 156.210 4.280 ;
        RECT 157.050 0.835 157.590 4.280 ;
        RECT 158.430 0.835 159.430 4.280 ;
        RECT 160.270 0.835 160.810 4.280 ;
        RECT 161.650 0.835 162.190 4.280 ;
        RECT 163.030 0.835 163.570 4.280 ;
        RECT 164.410 0.835 164.950 4.280 ;
        RECT 165.790 0.835 166.330 4.280 ;
        RECT 167.170 0.835 168.170 4.280 ;
        RECT 169.010 0.835 169.550 4.280 ;
        RECT 170.390 0.835 170.930 4.280 ;
        RECT 171.770 0.835 172.310 4.280 ;
        RECT 173.150 0.835 173.690 4.280 ;
        RECT 174.530 0.835 175.530 4.280 ;
        RECT 176.370 0.835 176.910 4.280 ;
        RECT 177.750 0.835 178.290 4.280 ;
        RECT 179.130 0.835 179.670 4.280 ;
        RECT 180.510 0.835 181.050 4.280 ;
        RECT 181.890 0.835 182.430 4.280 ;
        RECT 183.270 0.835 184.270 4.280 ;
        RECT 185.110 0.835 185.650 4.280 ;
        RECT 186.490 0.835 187.030 4.280 ;
        RECT 187.870 0.835 188.410 4.280 ;
        RECT 189.250 0.835 189.790 4.280 ;
        RECT 190.630 0.835 191.170 4.280 ;
        RECT 192.010 0.835 193.010 4.280 ;
        RECT 193.850 0.835 194.390 4.280 ;
        RECT 195.230 0.835 195.770 4.280 ;
        RECT 196.610 0.835 197.150 4.280 ;
        RECT 197.990 0.835 198.530 4.280 ;
        RECT 199.370 0.835 199.540 4.280 ;
      LAYER met3 ;
        RECT 4.000 598.080 195.600 598.225 ;
        RECT 4.400 597.360 195.600 598.080 ;
        RECT 4.400 596.720 196.000 597.360 ;
        RECT 4.400 596.680 195.600 596.720 ;
        RECT 4.000 595.320 195.600 596.680 ;
        RECT 4.000 594.680 196.000 595.320 ;
        RECT 4.000 594.000 195.600 594.680 ;
        RECT 4.400 593.280 195.600 594.000 ;
        RECT 4.400 592.640 196.000 593.280 ;
        RECT 4.400 592.600 195.600 592.640 ;
        RECT 4.000 591.240 195.600 592.600 ;
        RECT 4.000 590.600 196.000 591.240 ;
        RECT 4.000 589.920 195.600 590.600 ;
        RECT 4.400 589.200 195.600 589.920 ;
        RECT 4.400 588.520 196.000 589.200 ;
        RECT 4.000 587.880 196.000 588.520 ;
        RECT 4.000 586.480 195.600 587.880 ;
        RECT 4.000 585.840 196.000 586.480 ;
        RECT 4.400 584.440 195.600 585.840 ;
        RECT 4.000 583.800 196.000 584.440 ;
        RECT 4.000 582.400 195.600 583.800 ;
        RECT 4.000 581.760 196.000 582.400 ;
        RECT 4.400 580.360 195.600 581.760 ;
        RECT 4.000 579.720 196.000 580.360 ;
        RECT 4.000 578.320 195.600 579.720 ;
        RECT 4.000 577.680 196.000 578.320 ;
        RECT 4.400 576.280 195.600 577.680 ;
        RECT 4.000 574.960 196.000 576.280 ;
        RECT 4.000 573.600 195.600 574.960 ;
        RECT 4.400 573.560 195.600 573.600 ;
        RECT 4.400 572.920 196.000 573.560 ;
        RECT 4.400 572.200 195.600 572.920 ;
        RECT 4.000 571.520 195.600 572.200 ;
        RECT 4.000 570.880 196.000 571.520 ;
        RECT 4.000 569.520 195.600 570.880 ;
        RECT 4.400 569.480 195.600 569.520 ;
        RECT 4.400 568.840 196.000 569.480 ;
        RECT 4.400 568.120 195.600 568.840 ;
        RECT 4.000 567.440 195.600 568.120 ;
        RECT 4.000 566.800 196.000 567.440 ;
        RECT 4.000 565.440 195.600 566.800 ;
        RECT 4.400 565.400 195.600 565.440 ;
        RECT 4.400 564.760 196.000 565.400 ;
        RECT 4.400 564.040 195.600 564.760 ;
        RECT 4.000 563.360 195.600 564.040 ;
        RECT 4.000 562.040 196.000 563.360 ;
        RECT 4.000 561.360 195.600 562.040 ;
        RECT 4.400 560.640 195.600 561.360 ;
        RECT 4.400 560.000 196.000 560.640 ;
        RECT 4.400 559.960 195.600 560.000 ;
        RECT 4.000 558.600 195.600 559.960 ;
        RECT 4.000 557.960 196.000 558.600 ;
        RECT 4.000 557.280 195.600 557.960 ;
        RECT 4.400 556.560 195.600 557.280 ;
        RECT 4.400 555.920 196.000 556.560 ;
        RECT 4.400 555.880 195.600 555.920 ;
        RECT 4.000 554.520 195.600 555.880 ;
        RECT 4.000 553.880 196.000 554.520 ;
        RECT 4.000 553.200 195.600 553.880 ;
        RECT 4.400 552.480 195.600 553.200 ;
        RECT 4.400 551.840 196.000 552.480 ;
        RECT 4.400 551.800 195.600 551.840 ;
        RECT 4.000 550.440 195.600 551.800 ;
        RECT 4.000 549.120 196.000 550.440 ;
        RECT 4.000 548.440 195.600 549.120 ;
        RECT 4.400 547.720 195.600 548.440 ;
        RECT 4.400 547.080 196.000 547.720 ;
        RECT 4.400 547.040 195.600 547.080 ;
        RECT 4.000 545.680 195.600 547.040 ;
        RECT 4.000 545.040 196.000 545.680 ;
        RECT 4.000 544.360 195.600 545.040 ;
        RECT 4.400 543.640 195.600 544.360 ;
        RECT 4.400 543.000 196.000 543.640 ;
        RECT 4.400 542.960 195.600 543.000 ;
        RECT 4.000 541.600 195.600 542.960 ;
        RECT 4.000 540.960 196.000 541.600 ;
        RECT 4.000 540.280 195.600 540.960 ;
        RECT 4.400 539.560 195.600 540.280 ;
        RECT 4.400 538.880 196.000 539.560 ;
        RECT 4.000 538.240 196.000 538.880 ;
        RECT 4.000 536.840 195.600 538.240 ;
        RECT 4.000 536.200 196.000 536.840 ;
        RECT 4.400 534.800 195.600 536.200 ;
        RECT 4.000 534.160 196.000 534.800 ;
        RECT 4.000 532.760 195.600 534.160 ;
        RECT 4.000 532.120 196.000 532.760 ;
        RECT 4.400 530.720 195.600 532.120 ;
        RECT 4.000 530.080 196.000 530.720 ;
        RECT 4.000 528.680 195.600 530.080 ;
        RECT 4.000 528.040 196.000 528.680 ;
        RECT 4.400 526.640 195.600 528.040 ;
        RECT 4.000 525.320 196.000 526.640 ;
        RECT 4.000 523.960 195.600 525.320 ;
        RECT 4.400 523.920 195.600 523.960 ;
        RECT 4.400 523.280 196.000 523.920 ;
        RECT 4.400 522.560 195.600 523.280 ;
        RECT 4.000 521.880 195.600 522.560 ;
        RECT 4.000 521.240 196.000 521.880 ;
        RECT 4.000 519.880 195.600 521.240 ;
        RECT 4.400 519.840 195.600 519.880 ;
        RECT 4.400 519.200 196.000 519.840 ;
        RECT 4.400 518.480 195.600 519.200 ;
        RECT 4.000 517.800 195.600 518.480 ;
        RECT 4.000 517.160 196.000 517.800 ;
        RECT 4.000 515.800 195.600 517.160 ;
        RECT 4.400 515.760 195.600 515.800 ;
        RECT 4.400 515.120 196.000 515.760 ;
        RECT 4.400 514.400 195.600 515.120 ;
        RECT 4.000 513.720 195.600 514.400 ;
        RECT 4.000 512.400 196.000 513.720 ;
        RECT 4.000 511.720 195.600 512.400 ;
        RECT 4.400 511.000 195.600 511.720 ;
        RECT 4.400 510.360 196.000 511.000 ;
        RECT 4.400 510.320 195.600 510.360 ;
        RECT 4.000 508.960 195.600 510.320 ;
        RECT 4.000 508.320 196.000 508.960 ;
        RECT 4.000 507.640 195.600 508.320 ;
        RECT 4.400 506.920 195.600 507.640 ;
        RECT 4.400 506.280 196.000 506.920 ;
        RECT 4.400 506.240 195.600 506.280 ;
        RECT 4.000 504.880 195.600 506.240 ;
        RECT 4.000 504.240 196.000 504.880 ;
        RECT 4.000 503.560 195.600 504.240 ;
        RECT 4.400 502.840 195.600 503.560 ;
        RECT 4.400 502.200 196.000 502.840 ;
        RECT 4.400 502.160 195.600 502.200 ;
        RECT 4.000 500.800 195.600 502.160 ;
        RECT 4.000 499.480 196.000 500.800 ;
        RECT 4.000 498.800 195.600 499.480 ;
        RECT 4.400 498.080 195.600 498.800 ;
        RECT 4.400 497.440 196.000 498.080 ;
        RECT 4.400 497.400 195.600 497.440 ;
        RECT 4.000 496.040 195.600 497.400 ;
        RECT 4.000 495.400 196.000 496.040 ;
        RECT 4.000 494.720 195.600 495.400 ;
        RECT 4.400 494.000 195.600 494.720 ;
        RECT 4.400 493.360 196.000 494.000 ;
        RECT 4.400 493.320 195.600 493.360 ;
        RECT 4.000 491.960 195.600 493.320 ;
        RECT 4.000 491.320 196.000 491.960 ;
        RECT 4.000 490.640 195.600 491.320 ;
        RECT 4.400 489.920 195.600 490.640 ;
        RECT 4.400 489.280 196.000 489.920 ;
        RECT 4.400 489.240 195.600 489.280 ;
        RECT 4.000 487.880 195.600 489.240 ;
        RECT 4.000 486.560 196.000 487.880 ;
        RECT 4.400 485.160 195.600 486.560 ;
        RECT 4.000 484.520 196.000 485.160 ;
        RECT 4.000 483.120 195.600 484.520 ;
        RECT 4.000 482.480 196.000 483.120 ;
        RECT 4.400 481.080 195.600 482.480 ;
        RECT 4.000 480.440 196.000 481.080 ;
        RECT 4.000 479.040 195.600 480.440 ;
        RECT 4.000 478.400 196.000 479.040 ;
        RECT 4.400 477.000 195.600 478.400 ;
        RECT 4.000 475.680 196.000 477.000 ;
        RECT 4.000 474.320 195.600 475.680 ;
        RECT 4.400 474.280 195.600 474.320 ;
        RECT 4.400 473.640 196.000 474.280 ;
        RECT 4.400 472.920 195.600 473.640 ;
        RECT 4.000 472.240 195.600 472.920 ;
        RECT 4.000 471.600 196.000 472.240 ;
        RECT 4.000 470.240 195.600 471.600 ;
        RECT 4.400 470.200 195.600 470.240 ;
        RECT 4.400 469.560 196.000 470.200 ;
        RECT 4.400 468.840 195.600 469.560 ;
        RECT 4.000 468.160 195.600 468.840 ;
        RECT 4.000 467.520 196.000 468.160 ;
        RECT 4.000 466.160 195.600 467.520 ;
        RECT 4.400 466.120 195.600 466.160 ;
        RECT 4.400 465.480 196.000 466.120 ;
        RECT 4.400 464.760 195.600 465.480 ;
        RECT 4.000 464.080 195.600 464.760 ;
        RECT 4.000 462.760 196.000 464.080 ;
        RECT 4.000 462.080 195.600 462.760 ;
        RECT 4.400 461.360 195.600 462.080 ;
        RECT 4.400 460.720 196.000 461.360 ;
        RECT 4.400 460.680 195.600 460.720 ;
        RECT 4.000 459.320 195.600 460.680 ;
        RECT 4.000 458.680 196.000 459.320 ;
        RECT 4.000 458.000 195.600 458.680 ;
        RECT 4.400 457.280 195.600 458.000 ;
        RECT 4.400 456.640 196.000 457.280 ;
        RECT 4.400 456.600 195.600 456.640 ;
        RECT 4.000 455.240 195.600 456.600 ;
        RECT 4.000 454.600 196.000 455.240 ;
        RECT 4.000 453.920 195.600 454.600 ;
        RECT 4.400 453.200 195.600 453.920 ;
        RECT 4.400 452.560 196.000 453.200 ;
        RECT 4.400 452.520 195.600 452.560 ;
        RECT 4.000 451.160 195.600 452.520 ;
        RECT 4.000 449.840 196.000 451.160 ;
        RECT 4.000 449.160 195.600 449.840 ;
        RECT 4.400 448.440 195.600 449.160 ;
        RECT 4.400 447.800 196.000 448.440 ;
        RECT 4.400 447.760 195.600 447.800 ;
        RECT 4.000 446.400 195.600 447.760 ;
        RECT 4.000 445.760 196.000 446.400 ;
        RECT 4.000 445.080 195.600 445.760 ;
        RECT 4.400 444.360 195.600 445.080 ;
        RECT 4.400 443.720 196.000 444.360 ;
        RECT 4.400 443.680 195.600 443.720 ;
        RECT 4.000 442.320 195.600 443.680 ;
        RECT 4.000 441.680 196.000 442.320 ;
        RECT 4.000 441.000 195.600 441.680 ;
        RECT 4.400 440.280 195.600 441.000 ;
        RECT 4.400 439.640 196.000 440.280 ;
        RECT 4.400 439.600 195.600 439.640 ;
        RECT 4.000 438.240 195.600 439.600 ;
        RECT 4.000 436.920 196.000 438.240 ;
        RECT 4.400 435.520 195.600 436.920 ;
        RECT 4.000 434.880 196.000 435.520 ;
        RECT 4.000 433.480 195.600 434.880 ;
        RECT 4.000 432.840 196.000 433.480 ;
        RECT 4.400 431.440 195.600 432.840 ;
        RECT 4.000 430.800 196.000 431.440 ;
        RECT 4.000 429.400 195.600 430.800 ;
        RECT 4.000 428.760 196.000 429.400 ;
        RECT 4.400 427.360 195.600 428.760 ;
        RECT 4.000 426.720 196.000 427.360 ;
        RECT 4.000 425.320 195.600 426.720 ;
        RECT 4.000 424.680 196.000 425.320 ;
        RECT 4.400 424.000 196.000 424.680 ;
        RECT 4.400 423.280 195.600 424.000 ;
        RECT 4.000 422.600 195.600 423.280 ;
        RECT 4.000 421.960 196.000 422.600 ;
        RECT 4.000 420.600 195.600 421.960 ;
        RECT 4.400 420.560 195.600 420.600 ;
        RECT 4.400 419.920 196.000 420.560 ;
        RECT 4.400 419.200 195.600 419.920 ;
        RECT 4.000 418.520 195.600 419.200 ;
        RECT 4.000 417.880 196.000 418.520 ;
        RECT 4.000 416.520 195.600 417.880 ;
        RECT 4.400 416.480 195.600 416.520 ;
        RECT 4.400 415.840 196.000 416.480 ;
        RECT 4.400 415.120 195.600 415.840 ;
        RECT 4.000 414.440 195.600 415.120 ;
        RECT 4.000 413.120 196.000 414.440 ;
        RECT 4.000 412.440 195.600 413.120 ;
        RECT 4.400 411.720 195.600 412.440 ;
        RECT 4.400 411.080 196.000 411.720 ;
        RECT 4.400 411.040 195.600 411.080 ;
        RECT 4.000 409.680 195.600 411.040 ;
        RECT 4.000 409.040 196.000 409.680 ;
        RECT 4.000 408.360 195.600 409.040 ;
        RECT 4.400 407.640 195.600 408.360 ;
        RECT 4.400 407.000 196.000 407.640 ;
        RECT 4.400 406.960 195.600 407.000 ;
        RECT 4.000 405.600 195.600 406.960 ;
        RECT 4.000 404.960 196.000 405.600 ;
        RECT 4.000 404.280 195.600 404.960 ;
        RECT 4.400 403.560 195.600 404.280 ;
        RECT 4.400 402.920 196.000 403.560 ;
        RECT 4.400 402.880 195.600 402.920 ;
        RECT 4.000 401.520 195.600 402.880 ;
        RECT 4.000 400.200 196.000 401.520 ;
        RECT 4.000 399.520 195.600 400.200 ;
        RECT 4.400 398.800 195.600 399.520 ;
        RECT 4.400 398.160 196.000 398.800 ;
        RECT 4.400 398.120 195.600 398.160 ;
        RECT 4.000 396.760 195.600 398.120 ;
        RECT 4.000 396.120 196.000 396.760 ;
        RECT 4.000 395.440 195.600 396.120 ;
        RECT 4.400 394.720 195.600 395.440 ;
        RECT 4.400 394.080 196.000 394.720 ;
        RECT 4.400 394.040 195.600 394.080 ;
        RECT 4.000 392.680 195.600 394.040 ;
        RECT 4.000 392.040 196.000 392.680 ;
        RECT 4.000 391.360 195.600 392.040 ;
        RECT 4.400 390.640 195.600 391.360 ;
        RECT 4.400 390.000 196.000 390.640 ;
        RECT 4.400 389.960 195.600 390.000 ;
        RECT 4.000 388.600 195.600 389.960 ;
        RECT 4.000 387.280 196.000 388.600 ;
        RECT 4.400 385.880 195.600 387.280 ;
        RECT 4.000 385.240 196.000 385.880 ;
        RECT 4.000 383.840 195.600 385.240 ;
        RECT 4.000 383.200 196.000 383.840 ;
        RECT 4.400 381.800 195.600 383.200 ;
        RECT 4.000 381.160 196.000 381.800 ;
        RECT 4.000 379.760 195.600 381.160 ;
        RECT 4.000 379.120 196.000 379.760 ;
        RECT 4.400 377.720 195.600 379.120 ;
        RECT 4.000 377.080 196.000 377.720 ;
        RECT 4.000 375.680 195.600 377.080 ;
        RECT 4.000 375.040 196.000 375.680 ;
        RECT 4.400 374.360 196.000 375.040 ;
        RECT 4.400 373.640 195.600 374.360 ;
        RECT 4.000 372.960 195.600 373.640 ;
        RECT 4.000 372.320 196.000 372.960 ;
        RECT 4.000 370.960 195.600 372.320 ;
        RECT 4.400 370.920 195.600 370.960 ;
        RECT 4.400 370.280 196.000 370.920 ;
        RECT 4.400 369.560 195.600 370.280 ;
        RECT 4.000 368.880 195.600 369.560 ;
        RECT 4.000 368.240 196.000 368.880 ;
        RECT 4.000 366.880 195.600 368.240 ;
        RECT 4.400 366.840 195.600 366.880 ;
        RECT 4.400 366.200 196.000 366.840 ;
        RECT 4.400 365.480 195.600 366.200 ;
        RECT 4.000 364.800 195.600 365.480 ;
        RECT 4.000 364.160 196.000 364.800 ;
        RECT 4.000 362.800 195.600 364.160 ;
        RECT 4.400 362.760 195.600 362.800 ;
        RECT 4.400 361.440 196.000 362.760 ;
        RECT 4.400 361.400 195.600 361.440 ;
        RECT 4.000 360.040 195.600 361.400 ;
        RECT 4.000 359.400 196.000 360.040 ;
        RECT 4.000 358.720 195.600 359.400 ;
        RECT 4.400 358.000 195.600 358.720 ;
        RECT 4.400 357.360 196.000 358.000 ;
        RECT 4.400 357.320 195.600 357.360 ;
        RECT 4.000 355.960 195.600 357.320 ;
        RECT 4.000 355.320 196.000 355.960 ;
        RECT 4.000 354.640 195.600 355.320 ;
        RECT 4.400 353.920 195.600 354.640 ;
        RECT 4.400 353.280 196.000 353.920 ;
        RECT 4.400 353.240 195.600 353.280 ;
        RECT 4.000 351.880 195.600 353.240 ;
        RECT 4.000 350.560 196.000 351.880 ;
        RECT 4.000 349.880 195.600 350.560 ;
        RECT 4.400 349.160 195.600 349.880 ;
        RECT 4.400 348.520 196.000 349.160 ;
        RECT 4.400 348.480 195.600 348.520 ;
        RECT 4.000 347.120 195.600 348.480 ;
        RECT 4.000 346.480 196.000 347.120 ;
        RECT 4.000 345.800 195.600 346.480 ;
        RECT 4.400 345.080 195.600 345.800 ;
        RECT 4.400 344.440 196.000 345.080 ;
        RECT 4.400 344.400 195.600 344.440 ;
        RECT 4.000 343.040 195.600 344.400 ;
        RECT 4.000 342.400 196.000 343.040 ;
        RECT 4.000 341.720 195.600 342.400 ;
        RECT 4.400 341.000 195.600 341.720 ;
        RECT 4.400 340.360 196.000 341.000 ;
        RECT 4.400 340.320 195.600 340.360 ;
        RECT 4.000 338.960 195.600 340.320 ;
        RECT 4.000 337.640 196.000 338.960 ;
        RECT 4.400 336.240 195.600 337.640 ;
        RECT 4.000 335.600 196.000 336.240 ;
        RECT 4.000 334.200 195.600 335.600 ;
        RECT 4.000 333.560 196.000 334.200 ;
        RECT 4.400 332.160 195.600 333.560 ;
        RECT 4.000 331.520 196.000 332.160 ;
        RECT 4.000 330.120 195.600 331.520 ;
        RECT 4.000 329.480 196.000 330.120 ;
        RECT 4.400 328.080 195.600 329.480 ;
        RECT 4.000 327.440 196.000 328.080 ;
        RECT 4.000 326.040 195.600 327.440 ;
        RECT 4.000 325.400 196.000 326.040 ;
        RECT 4.400 324.720 196.000 325.400 ;
        RECT 4.400 324.000 195.600 324.720 ;
        RECT 4.000 323.320 195.600 324.000 ;
        RECT 4.000 322.680 196.000 323.320 ;
        RECT 4.000 321.320 195.600 322.680 ;
        RECT 4.400 321.280 195.600 321.320 ;
        RECT 4.400 320.640 196.000 321.280 ;
        RECT 4.400 319.920 195.600 320.640 ;
        RECT 4.000 319.240 195.600 319.920 ;
        RECT 4.000 318.600 196.000 319.240 ;
        RECT 4.000 317.240 195.600 318.600 ;
        RECT 4.400 317.200 195.600 317.240 ;
        RECT 4.400 316.560 196.000 317.200 ;
        RECT 4.400 315.840 195.600 316.560 ;
        RECT 4.000 315.160 195.600 315.840 ;
        RECT 4.000 314.520 196.000 315.160 ;
        RECT 4.000 313.160 195.600 314.520 ;
        RECT 4.400 313.120 195.600 313.160 ;
        RECT 4.400 311.800 196.000 313.120 ;
        RECT 4.400 311.760 195.600 311.800 ;
        RECT 4.000 310.400 195.600 311.760 ;
        RECT 4.000 309.760 196.000 310.400 ;
        RECT 4.000 309.080 195.600 309.760 ;
        RECT 4.400 308.360 195.600 309.080 ;
        RECT 4.400 307.720 196.000 308.360 ;
        RECT 4.400 307.680 195.600 307.720 ;
        RECT 4.000 306.320 195.600 307.680 ;
        RECT 4.000 305.680 196.000 306.320 ;
        RECT 4.000 305.000 195.600 305.680 ;
        RECT 4.400 304.280 195.600 305.000 ;
        RECT 4.400 303.640 196.000 304.280 ;
        RECT 4.400 303.600 195.600 303.640 ;
        RECT 4.000 302.240 195.600 303.600 ;
        RECT 4.000 301.600 196.000 302.240 ;
        RECT 4.000 300.240 195.600 301.600 ;
        RECT 4.400 300.200 195.600 300.240 ;
        RECT 4.400 298.880 196.000 300.200 ;
        RECT 4.400 298.840 195.600 298.880 ;
        RECT 4.000 297.480 195.600 298.840 ;
        RECT 4.000 296.840 196.000 297.480 ;
        RECT 4.000 296.160 195.600 296.840 ;
        RECT 4.400 295.440 195.600 296.160 ;
        RECT 4.400 294.800 196.000 295.440 ;
        RECT 4.400 294.760 195.600 294.800 ;
        RECT 4.000 293.400 195.600 294.760 ;
        RECT 4.000 292.760 196.000 293.400 ;
        RECT 4.000 292.080 195.600 292.760 ;
        RECT 4.400 291.360 195.600 292.080 ;
        RECT 4.400 290.720 196.000 291.360 ;
        RECT 4.400 290.680 195.600 290.720 ;
        RECT 4.000 289.320 195.600 290.680 ;
        RECT 4.000 288.000 196.000 289.320 ;
        RECT 4.400 286.600 195.600 288.000 ;
        RECT 4.000 285.960 196.000 286.600 ;
        RECT 4.000 284.560 195.600 285.960 ;
        RECT 4.000 283.920 196.000 284.560 ;
        RECT 4.400 282.520 195.600 283.920 ;
        RECT 4.000 281.880 196.000 282.520 ;
        RECT 4.000 280.480 195.600 281.880 ;
        RECT 4.000 279.840 196.000 280.480 ;
        RECT 4.400 278.440 195.600 279.840 ;
        RECT 4.000 277.800 196.000 278.440 ;
        RECT 4.000 276.400 195.600 277.800 ;
        RECT 4.000 275.760 196.000 276.400 ;
        RECT 4.400 275.080 196.000 275.760 ;
        RECT 4.400 274.360 195.600 275.080 ;
        RECT 4.000 273.680 195.600 274.360 ;
        RECT 4.000 273.040 196.000 273.680 ;
        RECT 4.000 271.680 195.600 273.040 ;
        RECT 4.400 271.640 195.600 271.680 ;
        RECT 4.400 271.000 196.000 271.640 ;
        RECT 4.400 270.280 195.600 271.000 ;
        RECT 4.000 269.600 195.600 270.280 ;
        RECT 4.000 268.960 196.000 269.600 ;
        RECT 4.000 267.600 195.600 268.960 ;
        RECT 4.400 267.560 195.600 267.600 ;
        RECT 4.400 266.920 196.000 267.560 ;
        RECT 4.400 266.200 195.600 266.920 ;
        RECT 4.000 265.520 195.600 266.200 ;
        RECT 4.000 264.880 196.000 265.520 ;
        RECT 4.000 263.520 195.600 264.880 ;
        RECT 4.400 263.480 195.600 263.520 ;
        RECT 4.400 262.160 196.000 263.480 ;
        RECT 4.400 262.120 195.600 262.160 ;
        RECT 4.000 260.760 195.600 262.120 ;
        RECT 4.000 260.120 196.000 260.760 ;
        RECT 4.000 259.440 195.600 260.120 ;
        RECT 4.400 258.720 195.600 259.440 ;
        RECT 4.400 258.080 196.000 258.720 ;
        RECT 4.400 258.040 195.600 258.080 ;
        RECT 4.000 256.680 195.600 258.040 ;
        RECT 4.000 256.040 196.000 256.680 ;
        RECT 4.000 255.360 195.600 256.040 ;
        RECT 4.400 254.640 195.600 255.360 ;
        RECT 4.400 254.000 196.000 254.640 ;
        RECT 4.400 253.960 195.600 254.000 ;
        RECT 4.000 252.600 195.600 253.960 ;
        RECT 4.000 251.960 196.000 252.600 ;
        RECT 4.000 250.600 195.600 251.960 ;
        RECT 4.400 250.560 195.600 250.600 ;
        RECT 4.400 249.240 196.000 250.560 ;
        RECT 4.400 249.200 195.600 249.240 ;
        RECT 4.000 247.840 195.600 249.200 ;
        RECT 4.000 247.200 196.000 247.840 ;
        RECT 4.000 246.520 195.600 247.200 ;
        RECT 4.400 245.800 195.600 246.520 ;
        RECT 4.400 245.160 196.000 245.800 ;
        RECT 4.400 245.120 195.600 245.160 ;
        RECT 4.000 243.760 195.600 245.120 ;
        RECT 4.000 243.120 196.000 243.760 ;
        RECT 4.000 242.440 195.600 243.120 ;
        RECT 4.400 241.720 195.600 242.440 ;
        RECT 4.400 241.080 196.000 241.720 ;
        RECT 4.400 241.040 195.600 241.080 ;
        RECT 4.000 239.680 195.600 241.040 ;
        RECT 4.000 238.360 196.000 239.680 ;
        RECT 4.400 236.960 195.600 238.360 ;
        RECT 4.000 236.320 196.000 236.960 ;
        RECT 4.000 234.920 195.600 236.320 ;
        RECT 4.000 234.280 196.000 234.920 ;
        RECT 4.400 232.880 195.600 234.280 ;
        RECT 4.000 232.240 196.000 232.880 ;
        RECT 4.000 230.840 195.600 232.240 ;
        RECT 4.000 230.200 196.000 230.840 ;
        RECT 4.400 228.800 195.600 230.200 ;
        RECT 4.000 228.160 196.000 228.800 ;
        RECT 4.000 226.760 195.600 228.160 ;
        RECT 4.000 226.120 196.000 226.760 ;
        RECT 4.400 225.440 196.000 226.120 ;
        RECT 4.400 224.720 195.600 225.440 ;
        RECT 4.000 224.040 195.600 224.720 ;
        RECT 4.000 223.400 196.000 224.040 ;
        RECT 4.000 222.040 195.600 223.400 ;
        RECT 4.400 222.000 195.600 222.040 ;
        RECT 4.400 221.360 196.000 222.000 ;
        RECT 4.400 220.640 195.600 221.360 ;
        RECT 4.000 219.960 195.600 220.640 ;
        RECT 4.000 219.320 196.000 219.960 ;
        RECT 4.000 217.960 195.600 219.320 ;
        RECT 4.400 217.920 195.600 217.960 ;
        RECT 4.400 217.280 196.000 217.920 ;
        RECT 4.400 216.560 195.600 217.280 ;
        RECT 4.000 215.880 195.600 216.560 ;
        RECT 4.000 215.240 196.000 215.880 ;
        RECT 4.000 213.880 195.600 215.240 ;
        RECT 4.400 213.840 195.600 213.880 ;
        RECT 4.400 212.520 196.000 213.840 ;
        RECT 4.400 212.480 195.600 212.520 ;
        RECT 4.000 211.120 195.600 212.480 ;
        RECT 4.000 210.480 196.000 211.120 ;
        RECT 4.000 209.800 195.600 210.480 ;
        RECT 4.400 209.080 195.600 209.800 ;
        RECT 4.400 208.440 196.000 209.080 ;
        RECT 4.400 208.400 195.600 208.440 ;
        RECT 4.000 207.040 195.600 208.400 ;
        RECT 4.000 206.400 196.000 207.040 ;
        RECT 4.000 205.720 195.600 206.400 ;
        RECT 4.400 205.000 195.600 205.720 ;
        RECT 4.400 204.360 196.000 205.000 ;
        RECT 4.400 204.320 195.600 204.360 ;
        RECT 4.000 202.960 195.600 204.320 ;
        RECT 4.000 202.320 196.000 202.960 ;
        RECT 4.000 200.960 195.600 202.320 ;
        RECT 4.400 200.920 195.600 200.960 ;
        RECT 4.400 199.600 196.000 200.920 ;
        RECT 4.400 199.560 195.600 199.600 ;
        RECT 4.000 198.200 195.600 199.560 ;
        RECT 4.000 197.560 196.000 198.200 ;
        RECT 4.000 196.880 195.600 197.560 ;
        RECT 4.400 196.160 195.600 196.880 ;
        RECT 4.400 195.520 196.000 196.160 ;
        RECT 4.400 195.480 195.600 195.520 ;
        RECT 4.000 194.120 195.600 195.480 ;
        RECT 4.000 193.480 196.000 194.120 ;
        RECT 4.000 192.800 195.600 193.480 ;
        RECT 4.400 192.080 195.600 192.800 ;
        RECT 4.400 191.440 196.000 192.080 ;
        RECT 4.400 191.400 195.600 191.440 ;
        RECT 4.000 190.040 195.600 191.400 ;
        RECT 4.000 189.400 196.000 190.040 ;
        RECT 4.000 188.720 195.600 189.400 ;
        RECT 4.400 188.000 195.600 188.720 ;
        RECT 4.400 187.320 196.000 188.000 ;
        RECT 4.000 186.680 196.000 187.320 ;
        RECT 4.000 185.280 195.600 186.680 ;
        RECT 4.000 184.640 196.000 185.280 ;
        RECT 4.400 183.240 195.600 184.640 ;
        RECT 4.000 182.600 196.000 183.240 ;
        RECT 4.000 181.200 195.600 182.600 ;
        RECT 4.000 180.560 196.000 181.200 ;
        RECT 4.400 179.160 195.600 180.560 ;
        RECT 4.000 178.520 196.000 179.160 ;
        RECT 4.000 177.120 195.600 178.520 ;
        RECT 4.000 176.480 196.000 177.120 ;
        RECT 4.400 175.800 196.000 176.480 ;
        RECT 4.400 175.080 195.600 175.800 ;
        RECT 4.000 174.400 195.600 175.080 ;
        RECT 4.000 173.760 196.000 174.400 ;
        RECT 4.000 172.400 195.600 173.760 ;
        RECT 4.400 172.360 195.600 172.400 ;
        RECT 4.400 171.720 196.000 172.360 ;
        RECT 4.400 171.000 195.600 171.720 ;
        RECT 4.000 170.320 195.600 171.000 ;
        RECT 4.000 169.680 196.000 170.320 ;
        RECT 4.000 168.320 195.600 169.680 ;
        RECT 4.400 168.280 195.600 168.320 ;
        RECT 4.400 167.640 196.000 168.280 ;
        RECT 4.400 166.920 195.600 167.640 ;
        RECT 4.000 166.240 195.600 166.920 ;
        RECT 4.000 165.600 196.000 166.240 ;
        RECT 4.000 164.240 195.600 165.600 ;
        RECT 4.400 164.200 195.600 164.240 ;
        RECT 4.400 162.880 196.000 164.200 ;
        RECT 4.400 162.840 195.600 162.880 ;
        RECT 4.000 161.480 195.600 162.840 ;
        RECT 4.000 160.840 196.000 161.480 ;
        RECT 4.000 160.160 195.600 160.840 ;
        RECT 4.400 159.440 195.600 160.160 ;
        RECT 4.400 158.800 196.000 159.440 ;
        RECT 4.400 158.760 195.600 158.800 ;
        RECT 4.000 157.400 195.600 158.760 ;
        RECT 4.000 156.760 196.000 157.400 ;
        RECT 4.000 156.080 195.600 156.760 ;
        RECT 4.400 155.360 195.600 156.080 ;
        RECT 4.400 154.720 196.000 155.360 ;
        RECT 4.400 154.680 195.600 154.720 ;
        RECT 4.000 153.320 195.600 154.680 ;
        RECT 4.000 152.680 196.000 153.320 ;
        RECT 4.000 151.320 195.600 152.680 ;
        RECT 4.400 151.280 195.600 151.320 ;
        RECT 4.400 149.960 196.000 151.280 ;
        RECT 4.400 149.920 195.600 149.960 ;
        RECT 4.000 148.560 195.600 149.920 ;
        RECT 4.000 147.920 196.000 148.560 ;
        RECT 4.000 147.240 195.600 147.920 ;
        RECT 4.400 146.520 195.600 147.240 ;
        RECT 4.400 145.880 196.000 146.520 ;
        RECT 4.400 145.840 195.600 145.880 ;
        RECT 4.000 144.480 195.600 145.840 ;
        RECT 4.000 143.840 196.000 144.480 ;
        RECT 4.000 143.160 195.600 143.840 ;
        RECT 4.400 142.440 195.600 143.160 ;
        RECT 4.400 141.800 196.000 142.440 ;
        RECT 4.400 141.760 195.600 141.800 ;
        RECT 4.000 140.400 195.600 141.760 ;
        RECT 4.000 139.760 196.000 140.400 ;
        RECT 4.000 139.080 195.600 139.760 ;
        RECT 4.400 138.360 195.600 139.080 ;
        RECT 4.400 137.680 196.000 138.360 ;
        RECT 4.000 137.040 196.000 137.680 ;
        RECT 4.000 135.640 195.600 137.040 ;
        RECT 4.000 135.000 196.000 135.640 ;
        RECT 4.400 133.600 195.600 135.000 ;
        RECT 4.000 132.960 196.000 133.600 ;
        RECT 4.000 131.560 195.600 132.960 ;
        RECT 4.000 130.920 196.000 131.560 ;
        RECT 4.400 129.520 195.600 130.920 ;
        RECT 4.000 128.880 196.000 129.520 ;
        RECT 4.000 127.480 195.600 128.880 ;
        RECT 4.000 126.840 196.000 127.480 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 4.000 124.120 196.000 125.440 ;
        RECT 4.000 122.760 195.600 124.120 ;
        RECT 4.400 122.720 195.600 122.760 ;
        RECT 4.400 122.080 196.000 122.720 ;
        RECT 4.400 121.360 195.600 122.080 ;
        RECT 4.000 120.680 195.600 121.360 ;
        RECT 4.000 120.040 196.000 120.680 ;
        RECT 4.000 118.680 195.600 120.040 ;
        RECT 4.400 118.640 195.600 118.680 ;
        RECT 4.400 118.000 196.000 118.640 ;
        RECT 4.400 117.280 195.600 118.000 ;
        RECT 4.000 116.600 195.600 117.280 ;
        RECT 4.000 115.960 196.000 116.600 ;
        RECT 4.000 114.600 195.600 115.960 ;
        RECT 4.400 114.560 195.600 114.600 ;
        RECT 4.400 113.240 196.000 114.560 ;
        RECT 4.400 113.200 195.600 113.240 ;
        RECT 4.000 111.840 195.600 113.200 ;
        RECT 4.000 111.200 196.000 111.840 ;
        RECT 4.000 110.520 195.600 111.200 ;
        RECT 4.400 109.800 195.600 110.520 ;
        RECT 4.400 109.160 196.000 109.800 ;
        RECT 4.400 109.120 195.600 109.160 ;
        RECT 4.000 107.760 195.600 109.120 ;
        RECT 4.000 107.120 196.000 107.760 ;
        RECT 4.000 106.440 195.600 107.120 ;
        RECT 4.400 105.720 195.600 106.440 ;
        RECT 4.400 105.080 196.000 105.720 ;
        RECT 4.400 105.040 195.600 105.080 ;
        RECT 4.000 103.680 195.600 105.040 ;
        RECT 4.000 103.040 196.000 103.680 ;
        RECT 4.000 101.680 195.600 103.040 ;
        RECT 4.400 101.640 195.600 101.680 ;
        RECT 4.400 100.320 196.000 101.640 ;
        RECT 4.400 100.280 195.600 100.320 ;
        RECT 4.000 98.920 195.600 100.280 ;
        RECT 4.000 98.280 196.000 98.920 ;
        RECT 4.000 97.600 195.600 98.280 ;
        RECT 4.400 96.880 195.600 97.600 ;
        RECT 4.400 96.240 196.000 96.880 ;
        RECT 4.400 96.200 195.600 96.240 ;
        RECT 4.000 94.840 195.600 96.200 ;
        RECT 4.000 94.200 196.000 94.840 ;
        RECT 4.000 93.520 195.600 94.200 ;
        RECT 4.400 92.800 195.600 93.520 ;
        RECT 4.400 92.160 196.000 92.800 ;
        RECT 4.400 92.120 195.600 92.160 ;
        RECT 4.000 90.760 195.600 92.120 ;
        RECT 4.000 90.120 196.000 90.760 ;
        RECT 4.000 89.440 195.600 90.120 ;
        RECT 4.400 88.720 195.600 89.440 ;
        RECT 4.400 88.040 196.000 88.720 ;
        RECT 4.000 87.400 196.000 88.040 ;
        RECT 4.000 86.000 195.600 87.400 ;
        RECT 4.000 85.360 196.000 86.000 ;
        RECT 4.400 83.960 195.600 85.360 ;
        RECT 4.000 83.320 196.000 83.960 ;
        RECT 4.000 81.920 195.600 83.320 ;
        RECT 4.000 81.280 196.000 81.920 ;
        RECT 4.400 79.880 195.600 81.280 ;
        RECT 4.000 79.240 196.000 79.880 ;
        RECT 4.000 77.840 195.600 79.240 ;
        RECT 4.000 77.200 196.000 77.840 ;
        RECT 4.400 75.800 195.600 77.200 ;
        RECT 4.000 74.480 196.000 75.800 ;
        RECT 4.000 73.120 195.600 74.480 ;
        RECT 4.400 73.080 195.600 73.120 ;
        RECT 4.400 72.440 196.000 73.080 ;
        RECT 4.400 71.720 195.600 72.440 ;
        RECT 4.000 71.040 195.600 71.720 ;
        RECT 4.000 70.400 196.000 71.040 ;
        RECT 4.000 69.040 195.600 70.400 ;
        RECT 4.400 69.000 195.600 69.040 ;
        RECT 4.400 68.360 196.000 69.000 ;
        RECT 4.400 67.640 195.600 68.360 ;
        RECT 4.000 66.960 195.600 67.640 ;
        RECT 4.000 66.320 196.000 66.960 ;
        RECT 4.000 64.960 195.600 66.320 ;
        RECT 4.400 64.920 195.600 64.960 ;
        RECT 4.400 64.280 196.000 64.920 ;
        RECT 4.400 63.560 195.600 64.280 ;
        RECT 4.000 62.880 195.600 63.560 ;
        RECT 4.000 61.560 196.000 62.880 ;
        RECT 4.000 60.880 195.600 61.560 ;
        RECT 4.400 60.160 195.600 60.880 ;
        RECT 4.400 59.520 196.000 60.160 ;
        RECT 4.400 59.480 195.600 59.520 ;
        RECT 4.000 58.120 195.600 59.480 ;
        RECT 4.000 57.480 196.000 58.120 ;
        RECT 4.000 56.800 195.600 57.480 ;
        RECT 4.400 56.080 195.600 56.800 ;
        RECT 4.400 55.440 196.000 56.080 ;
        RECT 4.400 55.400 195.600 55.440 ;
        RECT 4.000 54.040 195.600 55.400 ;
        RECT 4.000 53.400 196.000 54.040 ;
        RECT 4.000 52.040 195.600 53.400 ;
        RECT 4.400 52.000 195.600 52.040 ;
        RECT 4.400 50.680 196.000 52.000 ;
        RECT 4.400 50.640 195.600 50.680 ;
        RECT 4.000 49.280 195.600 50.640 ;
        RECT 4.000 48.640 196.000 49.280 ;
        RECT 4.000 47.960 195.600 48.640 ;
        RECT 4.400 47.240 195.600 47.960 ;
        RECT 4.400 46.600 196.000 47.240 ;
        RECT 4.400 46.560 195.600 46.600 ;
        RECT 4.000 45.200 195.600 46.560 ;
        RECT 4.000 44.560 196.000 45.200 ;
        RECT 4.000 43.880 195.600 44.560 ;
        RECT 4.400 43.160 195.600 43.880 ;
        RECT 4.400 42.520 196.000 43.160 ;
        RECT 4.400 42.480 195.600 42.520 ;
        RECT 4.000 41.120 195.600 42.480 ;
        RECT 4.000 40.480 196.000 41.120 ;
        RECT 4.000 39.800 195.600 40.480 ;
        RECT 4.400 39.080 195.600 39.800 ;
        RECT 4.400 38.400 196.000 39.080 ;
        RECT 4.000 37.760 196.000 38.400 ;
        RECT 4.000 36.360 195.600 37.760 ;
        RECT 4.000 35.720 196.000 36.360 ;
        RECT 4.400 34.320 195.600 35.720 ;
        RECT 4.000 33.680 196.000 34.320 ;
        RECT 4.000 32.280 195.600 33.680 ;
        RECT 4.000 31.640 196.000 32.280 ;
        RECT 4.400 30.240 195.600 31.640 ;
        RECT 4.000 29.600 196.000 30.240 ;
        RECT 4.000 28.200 195.600 29.600 ;
        RECT 4.000 27.560 196.000 28.200 ;
        RECT 4.400 26.160 195.600 27.560 ;
        RECT 4.000 24.840 196.000 26.160 ;
        RECT 4.000 23.480 195.600 24.840 ;
        RECT 4.400 23.440 195.600 23.480 ;
        RECT 4.400 22.800 196.000 23.440 ;
        RECT 4.400 22.080 195.600 22.800 ;
        RECT 4.000 21.400 195.600 22.080 ;
        RECT 4.000 20.760 196.000 21.400 ;
        RECT 4.000 19.400 195.600 20.760 ;
        RECT 4.400 19.360 195.600 19.400 ;
        RECT 4.400 18.720 196.000 19.360 ;
        RECT 4.400 18.000 195.600 18.720 ;
        RECT 4.000 17.320 195.600 18.000 ;
        RECT 4.000 16.680 196.000 17.320 ;
        RECT 4.000 15.320 195.600 16.680 ;
        RECT 4.400 15.280 195.600 15.320 ;
        RECT 4.400 14.640 196.000 15.280 ;
        RECT 4.400 13.920 195.600 14.640 ;
        RECT 4.000 13.240 195.600 13.920 ;
        RECT 4.000 11.920 196.000 13.240 ;
        RECT 4.000 11.240 195.600 11.920 ;
        RECT 4.400 10.520 195.600 11.240 ;
        RECT 4.400 9.880 196.000 10.520 ;
        RECT 4.400 9.840 195.600 9.880 ;
        RECT 4.000 8.480 195.600 9.840 ;
        RECT 4.000 7.840 196.000 8.480 ;
        RECT 4.000 7.160 195.600 7.840 ;
        RECT 4.400 6.440 195.600 7.160 ;
        RECT 4.400 5.800 196.000 6.440 ;
        RECT 4.400 5.760 195.600 5.800 ;
        RECT 4.000 4.400 195.600 5.760 ;
        RECT 4.000 3.760 196.000 4.400 ;
        RECT 4.000 3.080 195.600 3.760 ;
        RECT 4.400 2.360 195.600 3.080 ;
        RECT 4.400 1.720 196.000 2.360 ;
        RECT 4.400 1.680 195.600 1.720 ;
        RECT 4.000 0.855 195.600 1.680 ;
  END
END wb_local
END LIBRARY

