magic
tech sky130A
magscale 1 2
timestamp 1624040992
<< obsli1 >>
rect 1104 2159 58880 53329
<< obsm1 >>
rect 106 1300 59786 54188
<< metal2 >>
rect 110 55200 166 56800
rect 386 55200 442 56800
rect 754 55200 810 56800
rect 1030 55200 1086 56800
rect 1398 55200 1454 56800
rect 1766 55200 1822 56800
rect 2042 55200 2098 56800
rect 2410 55200 2466 56800
rect 2686 55200 2742 56800
rect 3054 55200 3110 56800
rect 3422 55200 3478 56800
rect 3698 55200 3754 56800
rect 4066 55200 4122 56800
rect 4434 55200 4490 56800
rect 4710 55200 4766 56800
rect 5078 55200 5134 56800
rect 5354 55200 5410 56800
rect 5722 55200 5778 56800
rect 6090 55200 6146 56800
rect 6366 55200 6422 56800
rect 6734 55200 6790 56800
rect 7102 55200 7158 56800
rect 7378 55200 7434 56800
rect 7746 55200 7802 56800
rect 8022 55200 8078 56800
rect 8390 55200 8446 56800
rect 8758 55200 8814 56800
rect 9034 55200 9090 56800
rect 9402 55200 9458 56800
rect 9770 55200 9826 56800
rect 10046 55200 10102 56800
rect 10414 55200 10470 56800
rect 10690 55200 10746 56800
rect 11058 55200 11114 56800
rect 11426 55200 11482 56800
rect 11702 55200 11758 56800
rect 12070 55200 12126 56800
rect 12438 55200 12494 56800
rect 12714 55200 12770 56800
rect 13082 55200 13138 56800
rect 13358 55200 13414 56800
rect 13726 55200 13782 56800
rect 14094 55200 14150 56800
rect 14370 55200 14426 56800
rect 14738 55200 14794 56800
rect 15106 55200 15162 56800
rect 15382 55200 15438 56800
rect 15750 55200 15806 56800
rect 16026 55200 16082 56800
rect 16394 55200 16450 56800
rect 16762 55200 16818 56800
rect 17038 55200 17094 56800
rect 17406 55200 17462 56800
rect 17682 55200 17738 56800
rect 18050 55200 18106 56800
rect 18418 55200 18474 56800
rect 18694 55200 18750 56800
rect 19062 55200 19118 56800
rect 19430 55200 19486 56800
rect 19706 55200 19762 56800
rect 20074 55200 20130 56800
rect 20350 55200 20406 56800
rect 20718 55200 20774 56800
rect 21086 55200 21142 56800
rect 21362 55200 21418 56800
rect 21730 55200 21786 56800
rect 22098 55200 22154 56800
rect 22374 55200 22430 56800
rect 22742 55200 22798 56800
rect 23018 55200 23074 56800
rect 23386 55200 23442 56800
rect 23754 55200 23810 56800
rect 24030 55200 24086 56800
rect 24398 55200 24454 56800
rect 24766 55200 24822 56800
rect 25042 55200 25098 56800
rect 25410 55200 25466 56800
rect 25686 55200 25742 56800
rect 26054 55200 26110 56800
rect 26422 55200 26478 56800
rect 26698 55200 26754 56800
rect 27066 55200 27122 56800
rect 27434 55200 27490 56800
rect 27710 55200 27766 56800
rect 28078 55200 28134 56800
rect 28354 55200 28410 56800
rect 28722 55200 28778 56800
rect 29090 55200 29146 56800
rect 29366 55200 29422 56800
rect 29734 55200 29790 56800
rect 30102 55200 30158 56800
rect 30378 55200 30434 56800
rect 30746 55200 30802 56800
rect 31022 55200 31078 56800
rect 31390 55200 31446 56800
rect 31758 55200 31814 56800
rect 32034 55200 32090 56800
rect 32402 55200 32458 56800
rect 32678 55200 32734 56800
rect 33046 55200 33102 56800
rect 33414 55200 33470 56800
rect 33690 55200 33746 56800
rect 34058 55200 34114 56800
rect 34426 55200 34482 56800
rect 34702 55200 34758 56800
rect 35070 55200 35126 56800
rect 35346 55200 35402 56800
rect 35714 55200 35770 56800
rect 36082 55200 36138 56800
rect 36358 55200 36414 56800
rect 36726 55200 36782 56800
rect 37094 55200 37150 56800
rect 37370 55200 37426 56800
rect 37738 55200 37794 56800
rect 38014 55200 38070 56800
rect 38382 55200 38438 56800
rect 38750 55200 38806 56800
rect 39026 55200 39082 56800
rect 39394 55200 39450 56800
rect 39762 55200 39818 56800
rect 40038 55200 40094 56800
rect 40406 55200 40462 56800
rect 40682 55200 40738 56800
rect 41050 55200 41106 56800
rect 41418 55200 41474 56800
rect 41694 55200 41750 56800
rect 42062 55200 42118 56800
rect 42430 55200 42486 56800
rect 42706 55200 42762 56800
rect 43074 55200 43130 56800
rect 43350 55200 43406 56800
rect 43718 55200 43774 56800
rect 44086 55200 44142 56800
rect 44362 55200 44418 56800
rect 44730 55200 44786 56800
rect 45098 55200 45154 56800
rect 45374 55200 45430 56800
rect 45742 55200 45798 56800
rect 46018 55200 46074 56800
rect 46386 55200 46442 56800
rect 46754 55200 46810 56800
rect 47030 55200 47086 56800
rect 47398 55200 47454 56800
rect 47674 55200 47730 56800
rect 48042 55200 48098 56800
rect 48410 55200 48466 56800
rect 48686 55200 48742 56800
rect 49054 55200 49110 56800
rect 49422 55200 49478 56800
rect 49698 55200 49754 56800
rect 50066 55200 50122 56800
rect 50342 55200 50398 56800
rect 50710 55200 50766 56800
rect 51078 55200 51134 56800
rect 51354 55200 51410 56800
rect 51722 55200 51778 56800
rect 52090 55200 52146 56800
rect 52366 55200 52422 56800
rect 52734 55200 52790 56800
rect 53010 55200 53066 56800
rect 53378 55200 53434 56800
rect 53746 55200 53802 56800
rect 54022 55200 54078 56800
rect 54390 55200 54446 56800
rect 54758 55200 54814 56800
rect 55034 55200 55090 56800
rect 55402 55200 55458 56800
rect 55678 55200 55734 56800
rect 56046 55200 56102 56800
rect 56414 55200 56470 56800
rect 56690 55200 56746 56800
rect 57058 55200 57114 56800
rect 57426 55200 57482 56800
rect 57702 55200 57758 56800
rect 58070 55200 58126 56800
rect 58346 55200 58402 56800
rect 58714 55200 58770 56800
rect 59082 55200 59138 56800
rect 59358 55200 59414 56800
rect 59726 55200 59782 56800
rect 662 -800 718 800
rect 1950 -800 2006 800
rect 3238 -800 3294 800
rect 4618 -800 4674 800
rect 5906 -800 5962 800
rect 7286 -800 7342 800
rect 8574 -800 8630 800
rect 9954 -800 10010 800
rect 11242 -800 11298 800
rect 12622 -800 12678 800
rect 13910 -800 13966 800
rect 15290 -800 15346 800
rect 16578 -800 16634 800
rect 17958 -800 18014 800
rect 19246 -800 19302 800
rect 20626 -800 20682 800
rect 21914 -800 21970 800
rect 23294 -800 23350 800
rect 24582 -800 24638 800
rect 25962 -800 26018 800
rect 27250 -800 27306 800
rect 28630 -800 28686 800
rect 29918 -800 29974 800
rect 31298 -800 31354 800
rect 32586 -800 32642 800
rect 33966 -800 34022 800
rect 35254 -800 35310 800
rect 36634 -800 36690 800
rect 37922 -800 37978 800
rect 39302 -800 39358 800
rect 40590 -800 40646 800
rect 41970 -800 42026 800
rect 43258 -800 43314 800
rect 44638 -800 44694 800
rect 45926 -800 45982 800
rect 47306 -800 47362 800
rect 48594 -800 48650 800
rect 49974 -800 50030 800
rect 51262 -800 51318 800
rect 52642 -800 52698 800
rect 53930 -800 53986 800
rect 55310 -800 55366 800
rect 56598 -800 56654 800
rect 57978 -800 58034 800
rect 59266 -800 59322 800
<< obsm2 >>
rect 222 55144 330 55593
rect 498 55144 698 55593
rect 866 55144 974 55593
rect 1142 55144 1342 55593
rect 1510 55144 1710 55593
rect 1878 55144 1986 55593
rect 2154 55144 2354 55593
rect 2522 55144 2630 55593
rect 2798 55144 2998 55593
rect 3166 55144 3366 55593
rect 3534 55144 3642 55593
rect 3810 55144 4010 55593
rect 4178 55144 4378 55593
rect 4546 55144 4654 55593
rect 4822 55144 5022 55593
rect 5190 55144 5298 55593
rect 5466 55144 5666 55593
rect 5834 55144 6034 55593
rect 6202 55144 6310 55593
rect 6478 55144 6678 55593
rect 6846 55144 7046 55593
rect 7214 55144 7322 55593
rect 7490 55144 7690 55593
rect 7858 55144 7966 55593
rect 8134 55144 8334 55593
rect 8502 55144 8702 55593
rect 8870 55144 8978 55593
rect 9146 55144 9346 55593
rect 9514 55144 9714 55593
rect 9882 55144 9990 55593
rect 10158 55144 10358 55593
rect 10526 55144 10634 55593
rect 10802 55144 11002 55593
rect 11170 55144 11370 55593
rect 11538 55144 11646 55593
rect 11814 55144 12014 55593
rect 12182 55144 12382 55593
rect 12550 55144 12658 55593
rect 12826 55144 13026 55593
rect 13194 55144 13302 55593
rect 13470 55144 13670 55593
rect 13838 55144 14038 55593
rect 14206 55144 14314 55593
rect 14482 55144 14682 55593
rect 14850 55144 15050 55593
rect 15218 55144 15326 55593
rect 15494 55144 15694 55593
rect 15862 55144 15970 55593
rect 16138 55144 16338 55593
rect 16506 55144 16706 55593
rect 16874 55144 16982 55593
rect 17150 55144 17350 55593
rect 17518 55144 17626 55593
rect 17794 55144 17994 55593
rect 18162 55144 18362 55593
rect 18530 55144 18638 55593
rect 18806 55144 19006 55593
rect 19174 55144 19374 55593
rect 19542 55144 19650 55593
rect 19818 55144 20018 55593
rect 20186 55144 20294 55593
rect 20462 55144 20662 55593
rect 20830 55144 21030 55593
rect 21198 55144 21306 55593
rect 21474 55144 21674 55593
rect 21842 55144 22042 55593
rect 22210 55144 22318 55593
rect 22486 55144 22686 55593
rect 22854 55144 22962 55593
rect 23130 55144 23330 55593
rect 23498 55144 23698 55593
rect 23866 55144 23974 55593
rect 24142 55144 24342 55593
rect 24510 55144 24710 55593
rect 24878 55144 24986 55593
rect 25154 55144 25354 55593
rect 25522 55144 25630 55593
rect 25798 55144 25998 55593
rect 26166 55144 26366 55593
rect 26534 55144 26642 55593
rect 26810 55144 27010 55593
rect 27178 55144 27378 55593
rect 27546 55144 27654 55593
rect 27822 55144 28022 55593
rect 28190 55144 28298 55593
rect 28466 55144 28666 55593
rect 28834 55144 29034 55593
rect 29202 55144 29310 55593
rect 29478 55144 29678 55593
rect 29846 55144 30046 55593
rect 30214 55144 30322 55593
rect 30490 55144 30690 55593
rect 30858 55144 30966 55593
rect 31134 55144 31334 55593
rect 31502 55144 31702 55593
rect 31870 55144 31978 55593
rect 32146 55144 32346 55593
rect 32514 55144 32622 55593
rect 32790 55144 32990 55593
rect 33158 55144 33358 55593
rect 33526 55144 33634 55593
rect 33802 55144 34002 55593
rect 34170 55144 34370 55593
rect 34538 55144 34646 55593
rect 34814 55144 35014 55593
rect 35182 55144 35290 55593
rect 35458 55144 35658 55593
rect 35826 55144 36026 55593
rect 36194 55144 36302 55593
rect 36470 55144 36670 55593
rect 36838 55144 37038 55593
rect 37206 55144 37314 55593
rect 37482 55144 37682 55593
rect 37850 55144 37958 55593
rect 38126 55144 38326 55593
rect 38494 55144 38694 55593
rect 38862 55144 38970 55593
rect 39138 55144 39338 55593
rect 39506 55144 39706 55593
rect 39874 55144 39982 55593
rect 40150 55144 40350 55593
rect 40518 55144 40626 55593
rect 40794 55144 40994 55593
rect 41162 55144 41362 55593
rect 41530 55144 41638 55593
rect 41806 55144 42006 55593
rect 42174 55144 42374 55593
rect 42542 55144 42650 55593
rect 42818 55144 43018 55593
rect 43186 55144 43294 55593
rect 43462 55144 43662 55593
rect 43830 55144 44030 55593
rect 44198 55144 44306 55593
rect 44474 55144 44674 55593
rect 44842 55144 45042 55593
rect 45210 55144 45318 55593
rect 45486 55144 45686 55593
rect 45854 55144 45962 55593
rect 46130 55144 46330 55593
rect 46498 55144 46698 55593
rect 46866 55144 46974 55593
rect 47142 55144 47342 55593
rect 47510 55144 47618 55593
rect 47786 55144 47986 55593
rect 48154 55144 48354 55593
rect 48522 55144 48630 55593
rect 48798 55144 48998 55593
rect 49166 55144 49366 55593
rect 49534 55144 49642 55593
rect 49810 55144 50010 55593
rect 50178 55144 50286 55593
rect 50454 55144 50654 55593
rect 50822 55144 51022 55593
rect 51190 55144 51298 55593
rect 51466 55144 51666 55593
rect 51834 55144 52034 55593
rect 52202 55144 52310 55593
rect 52478 55144 52678 55593
rect 52846 55144 52954 55593
rect 53122 55144 53322 55593
rect 53490 55144 53690 55593
rect 53858 55144 53966 55593
rect 54134 55144 54334 55593
rect 54502 55144 54702 55593
rect 54870 55144 54978 55593
rect 55146 55144 55346 55593
rect 55514 55144 55622 55593
rect 55790 55144 55990 55593
rect 56158 55144 56358 55593
rect 56526 55144 56634 55593
rect 56802 55144 57002 55593
rect 57170 55144 57370 55593
rect 57538 55144 57646 55593
rect 57814 55144 58014 55593
rect 58182 55144 58290 55593
rect 58458 55144 58658 55593
rect 58826 55144 59026 55593
rect 59194 55144 59302 55593
rect 59470 55144 59670 55593
rect 112 856 59780 55144
rect 112 303 606 856
rect 774 303 1894 856
rect 2062 303 3182 856
rect 3350 303 4562 856
rect 4730 303 5850 856
rect 6018 303 7230 856
rect 7398 303 8518 856
rect 8686 303 9898 856
rect 10066 303 11186 856
rect 11354 303 12566 856
rect 12734 303 13854 856
rect 14022 303 15234 856
rect 15402 303 16522 856
rect 16690 303 17902 856
rect 18070 303 19190 856
rect 19358 303 20570 856
rect 20738 303 21858 856
rect 22026 303 23238 856
rect 23406 303 24526 856
rect 24694 303 25906 856
rect 26074 303 27194 856
rect 27362 303 28574 856
rect 28742 303 29862 856
rect 30030 303 31242 856
rect 31410 303 32530 856
rect 32698 303 33910 856
rect 34078 303 35198 856
rect 35366 303 36578 856
rect 36746 303 37866 856
rect 38034 303 39246 856
rect 39414 303 40534 856
rect 40702 303 41914 856
rect 42082 303 43202 856
rect 43370 303 44582 856
rect 44750 303 45870 856
rect 46038 303 47250 856
rect 47418 303 48538 856
rect 48706 303 49918 856
rect 50086 303 51206 856
rect 51374 303 52586 856
rect 52754 303 53874 856
rect 54042 303 55254 856
rect 55422 303 56542 856
rect 56710 303 57922 856
rect 58090 303 59210 856
rect 59378 303 59780 856
<< metal3 >>
rect -800 55496 800 55616
rect 59200 55496 60800 55616
rect -800 54816 800 54936
rect 59200 54680 60800 54800
rect -800 54136 800 54256
rect 59200 53864 60800 53984
rect -800 53456 800 53576
rect 59200 53048 60800 53168
rect -800 52776 800 52896
rect -800 52096 800 52216
rect 59200 52232 60800 52352
rect -800 51416 800 51536
rect 59200 51416 60800 51536
rect -800 50736 800 50856
rect 59200 50464 60800 50584
rect -800 50056 800 50176
rect 59200 49648 60800 49768
rect -800 49376 800 49496
rect -800 48696 800 48816
rect 59200 48832 60800 48952
rect -800 47880 800 48000
rect 59200 48016 60800 48136
rect -800 47200 800 47320
rect 59200 47200 60800 47320
rect -800 46520 800 46640
rect 59200 46384 60800 46504
rect -800 45840 800 45960
rect 59200 45568 60800 45688
rect -800 45160 800 45280
rect -800 44480 800 44600
rect 59200 44616 60800 44736
rect -800 43800 800 43920
rect 59200 43800 60800 43920
rect -800 43120 800 43240
rect 59200 42984 60800 43104
rect -800 42440 800 42560
rect 59200 42168 60800 42288
rect -800 41760 800 41880
rect 59200 41352 60800 41472
rect -800 41080 800 41200
rect -800 40400 800 40520
rect 59200 40536 60800 40656
rect -800 39584 800 39704
rect 59200 39720 60800 39840
rect -800 38904 800 39024
rect 59200 38768 60800 38888
rect -800 38224 800 38344
rect 59200 37952 60800 38072
rect -800 37544 800 37664
rect 59200 37136 60800 37256
rect -800 36864 800 36984
rect -800 36184 800 36304
rect 59200 36320 60800 36440
rect -800 35504 800 35624
rect 59200 35504 60800 35624
rect -800 34824 800 34944
rect 59200 34688 60800 34808
rect -800 34144 800 34264
rect 59200 33736 60800 33856
rect -800 33464 800 33584
rect -800 32784 800 32904
rect 59200 32920 60800 33040
rect -800 31968 800 32088
rect 59200 32104 60800 32224
rect -800 31288 800 31408
rect 59200 31288 60800 31408
rect -800 30608 800 30728
rect 59200 30472 60800 30592
rect -800 29928 800 30048
rect 59200 29656 60800 29776
rect -800 29248 800 29368
rect 59200 28840 60800 28960
rect -800 28568 800 28688
rect -800 27888 800 28008
rect 59200 27888 60800 28008
rect -800 27208 800 27328
rect 59200 27072 60800 27192
rect -800 26528 800 26648
rect 59200 26256 60800 26376
rect -800 25848 800 25968
rect 59200 25440 60800 25560
rect -800 25168 800 25288
rect -800 24488 800 24608
rect 59200 24624 60800 24744
rect -800 23672 800 23792
rect 59200 23808 60800 23928
rect -800 22992 800 23112
rect 59200 22992 60800 23112
rect -800 22312 800 22432
rect 59200 22040 60800 22160
rect -800 21632 800 21752
rect 59200 21224 60800 21344
rect -800 20952 800 21072
rect -800 20272 800 20392
rect 59200 20408 60800 20528
rect -800 19592 800 19712
rect 59200 19592 60800 19712
rect -800 18912 800 19032
rect 59200 18776 60800 18896
rect -800 18232 800 18352
rect 59200 17960 60800 18080
rect -800 17552 800 17672
rect -800 16872 800 16992
rect 59200 17008 60800 17128
rect -800 16056 800 16176
rect 59200 16192 60800 16312
rect -800 15376 800 15496
rect 59200 15376 60800 15496
rect -800 14696 800 14816
rect 59200 14560 60800 14680
rect -800 14016 800 14136
rect 59200 13744 60800 13864
rect -800 13336 800 13456
rect 59200 12928 60800 13048
rect -800 12656 800 12776
rect -800 11976 800 12096
rect 59200 12112 60800 12232
rect -800 11296 800 11416
rect 59200 11160 60800 11280
rect -800 10616 800 10736
rect 59200 10344 60800 10464
rect -800 9936 800 10056
rect 59200 9528 60800 9648
rect -800 9256 800 9376
rect -800 8576 800 8696
rect 59200 8712 60800 8832
rect -800 7760 800 7880
rect 59200 7896 60800 8016
rect -800 7080 800 7200
rect 59200 7080 60800 7200
rect -800 6400 800 6520
rect 59200 6264 60800 6384
rect -800 5720 800 5840
rect 59200 5312 60800 5432
rect -800 5040 800 5160
rect -800 4360 800 4480
rect 59200 4496 60800 4616
rect -800 3680 800 3800
rect 59200 3680 60800 3800
rect -800 3000 800 3120
rect 59200 2864 60800 2984
rect -800 2320 800 2440
rect 59200 2048 60800 2168
rect -800 1640 800 1760
rect 59200 1232 60800 1352
rect -800 960 800 1080
rect -800 280 800 400
rect 59200 416 60800 536
<< obsm3 >>
rect 880 55416 59120 55589
rect 800 55016 59200 55416
rect 880 54880 59200 55016
rect 880 54736 59120 54880
rect 800 54600 59120 54736
rect 800 54336 59200 54600
rect 880 54064 59200 54336
rect 880 54056 59120 54064
rect 800 53784 59120 54056
rect 800 53656 59200 53784
rect 880 53376 59200 53656
rect 800 53248 59200 53376
rect 800 52976 59120 53248
rect 880 52968 59120 52976
rect 880 52696 59200 52968
rect 800 52432 59200 52696
rect 800 52296 59120 52432
rect 880 52152 59120 52296
rect 880 52016 59200 52152
rect 800 51616 59200 52016
rect 880 51336 59120 51616
rect 800 50936 59200 51336
rect 880 50664 59200 50936
rect 880 50656 59120 50664
rect 800 50384 59120 50656
rect 800 50256 59200 50384
rect 880 49976 59200 50256
rect 800 49848 59200 49976
rect 800 49576 59120 49848
rect 880 49568 59120 49576
rect 880 49296 59200 49568
rect 800 49032 59200 49296
rect 800 48896 59120 49032
rect 880 48752 59120 48896
rect 880 48616 59200 48752
rect 800 48216 59200 48616
rect 800 48080 59120 48216
rect 880 47936 59120 48080
rect 880 47800 59200 47936
rect 800 47400 59200 47800
rect 880 47120 59120 47400
rect 800 46720 59200 47120
rect 880 46584 59200 46720
rect 880 46440 59120 46584
rect 800 46304 59120 46440
rect 800 46040 59200 46304
rect 880 45768 59200 46040
rect 880 45760 59120 45768
rect 800 45488 59120 45760
rect 800 45360 59200 45488
rect 880 45080 59200 45360
rect 800 44816 59200 45080
rect 800 44680 59120 44816
rect 880 44536 59120 44680
rect 880 44400 59200 44536
rect 800 44000 59200 44400
rect 880 43720 59120 44000
rect 800 43320 59200 43720
rect 880 43184 59200 43320
rect 880 43040 59120 43184
rect 800 42904 59120 43040
rect 800 42640 59200 42904
rect 880 42368 59200 42640
rect 880 42360 59120 42368
rect 800 42088 59120 42360
rect 800 41960 59200 42088
rect 880 41680 59200 41960
rect 800 41552 59200 41680
rect 800 41280 59120 41552
rect 880 41272 59120 41280
rect 880 41000 59200 41272
rect 800 40736 59200 41000
rect 800 40600 59120 40736
rect 880 40456 59120 40600
rect 880 40320 59200 40456
rect 800 39920 59200 40320
rect 800 39784 59120 39920
rect 880 39640 59120 39784
rect 880 39504 59200 39640
rect 800 39104 59200 39504
rect 880 38968 59200 39104
rect 880 38824 59120 38968
rect 800 38688 59120 38824
rect 800 38424 59200 38688
rect 880 38152 59200 38424
rect 880 38144 59120 38152
rect 800 37872 59120 38144
rect 800 37744 59200 37872
rect 880 37464 59200 37744
rect 800 37336 59200 37464
rect 800 37064 59120 37336
rect 880 37056 59120 37064
rect 880 36784 59200 37056
rect 800 36520 59200 36784
rect 800 36384 59120 36520
rect 880 36240 59120 36384
rect 880 36104 59200 36240
rect 800 35704 59200 36104
rect 880 35424 59120 35704
rect 800 35024 59200 35424
rect 880 34888 59200 35024
rect 880 34744 59120 34888
rect 800 34608 59120 34744
rect 800 34344 59200 34608
rect 880 34064 59200 34344
rect 800 33936 59200 34064
rect 800 33664 59120 33936
rect 880 33656 59120 33664
rect 880 33384 59200 33656
rect 800 33120 59200 33384
rect 800 32984 59120 33120
rect 880 32840 59120 32984
rect 880 32704 59200 32840
rect 800 32304 59200 32704
rect 800 32168 59120 32304
rect 880 32024 59120 32168
rect 880 31888 59200 32024
rect 800 31488 59200 31888
rect 880 31208 59120 31488
rect 800 30808 59200 31208
rect 880 30672 59200 30808
rect 880 30528 59120 30672
rect 800 30392 59120 30528
rect 800 30128 59200 30392
rect 880 29856 59200 30128
rect 880 29848 59120 29856
rect 800 29576 59120 29848
rect 800 29448 59200 29576
rect 880 29168 59200 29448
rect 800 29040 59200 29168
rect 800 28768 59120 29040
rect 880 28760 59120 28768
rect 880 28488 59200 28760
rect 800 28088 59200 28488
rect 880 27808 59120 28088
rect 800 27408 59200 27808
rect 880 27272 59200 27408
rect 880 27128 59120 27272
rect 800 26992 59120 27128
rect 800 26728 59200 26992
rect 880 26456 59200 26728
rect 880 26448 59120 26456
rect 800 26176 59120 26448
rect 800 26048 59200 26176
rect 880 25768 59200 26048
rect 800 25640 59200 25768
rect 800 25368 59120 25640
rect 880 25360 59120 25368
rect 880 25088 59200 25360
rect 800 24824 59200 25088
rect 800 24688 59120 24824
rect 880 24544 59120 24688
rect 880 24408 59200 24544
rect 800 24008 59200 24408
rect 800 23872 59120 24008
rect 880 23728 59120 23872
rect 880 23592 59200 23728
rect 800 23192 59200 23592
rect 880 22912 59120 23192
rect 800 22512 59200 22912
rect 880 22240 59200 22512
rect 880 22232 59120 22240
rect 800 21960 59120 22232
rect 800 21832 59200 21960
rect 880 21552 59200 21832
rect 800 21424 59200 21552
rect 800 21152 59120 21424
rect 880 21144 59120 21152
rect 880 20872 59200 21144
rect 800 20608 59200 20872
rect 800 20472 59120 20608
rect 880 20328 59120 20472
rect 880 20192 59200 20328
rect 800 19792 59200 20192
rect 880 19512 59120 19792
rect 800 19112 59200 19512
rect 880 18976 59200 19112
rect 880 18832 59120 18976
rect 800 18696 59120 18832
rect 800 18432 59200 18696
rect 880 18160 59200 18432
rect 880 18152 59120 18160
rect 800 17880 59120 18152
rect 800 17752 59200 17880
rect 880 17472 59200 17752
rect 800 17208 59200 17472
rect 800 17072 59120 17208
rect 880 16928 59120 17072
rect 880 16792 59200 16928
rect 800 16392 59200 16792
rect 800 16256 59120 16392
rect 880 16112 59120 16256
rect 880 15976 59200 16112
rect 800 15576 59200 15976
rect 880 15296 59120 15576
rect 800 14896 59200 15296
rect 880 14760 59200 14896
rect 880 14616 59120 14760
rect 800 14480 59120 14616
rect 800 14216 59200 14480
rect 880 13944 59200 14216
rect 880 13936 59120 13944
rect 800 13664 59120 13936
rect 800 13536 59200 13664
rect 880 13256 59200 13536
rect 800 13128 59200 13256
rect 800 12856 59120 13128
rect 880 12848 59120 12856
rect 880 12576 59200 12848
rect 800 12312 59200 12576
rect 800 12176 59120 12312
rect 880 12032 59120 12176
rect 880 11896 59200 12032
rect 800 11496 59200 11896
rect 880 11360 59200 11496
rect 880 11216 59120 11360
rect 800 11080 59120 11216
rect 800 10816 59200 11080
rect 880 10544 59200 10816
rect 880 10536 59120 10544
rect 800 10264 59120 10536
rect 800 10136 59200 10264
rect 880 9856 59200 10136
rect 800 9728 59200 9856
rect 800 9456 59120 9728
rect 880 9448 59120 9456
rect 880 9176 59200 9448
rect 800 8912 59200 9176
rect 800 8776 59120 8912
rect 880 8632 59120 8776
rect 880 8496 59200 8632
rect 800 8096 59200 8496
rect 800 7960 59120 8096
rect 880 7816 59120 7960
rect 880 7680 59200 7816
rect 800 7280 59200 7680
rect 880 7000 59120 7280
rect 800 6600 59200 7000
rect 880 6464 59200 6600
rect 880 6320 59120 6464
rect 800 6184 59120 6320
rect 800 5920 59200 6184
rect 880 5640 59200 5920
rect 800 5512 59200 5640
rect 800 5240 59120 5512
rect 880 5232 59120 5240
rect 880 4960 59200 5232
rect 800 4696 59200 4960
rect 800 4560 59120 4696
rect 880 4416 59120 4560
rect 880 4280 59200 4416
rect 800 3880 59200 4280
rect 880 3600 59120 3880
rect 800 3200 59200 3600
rect 880 3064 59200 3200
rect 880 2920 59120 3064
rect 800 2784 59120 2920
rect 800 2520 59200 2784
rect 880 2248 59200 2520
rect 880 2240 59120 2248
rect 800 1968 59120 2240
rect 800 1840 59200 1968
rect 880 1560 59200 1840
rect 800 1432 59200 1560
rect 800 1160 59120 1432
rect 880 1152 59120 1160
rect 880 880 59200 1152
rect 800 616 59200 880
rect 800 480 59120 616
rect 880 336 59120 480
rect 880 307 59200 336
<< metal4 >>
rect 4208 2128 4528 53360
rect 19568 2128 19888 53360
rect 34928 2128 35248 53360
rect 50288 2128 50608 53360
<< labels >>
rlabel metal3 s -800 960 800 1080 4 io_ack_o
port 1 nsew signal output
rlabel metal3 s -800 2320 800 2440 4 io_adr_i[0]
port 2 nsew signal input
rlabel metal3 s -800 9256 800 9376 4 io_adr_i[10]
port 3 nsew signal input
rlabel metal3 s -800 9936 800 10056 4 io_adr_i[11]
port 4 nsew signal input
rlabel metal3 s -800 3000 800 3120 4 io_adr_i[1]
port 5 nsew signal input
rlabel metal3 s -800 3680 800 3800 4 io_adr_i[2]
port 6 nsew signal input
rlabel metal3 s -800 4360 800 4480 4 io_adr_i[3]
port 7 nsew signal input
rlabel metal3 s -800 5040 800 5160 4 io_adr_i[4]
port 8 nsew signal input
rlabel metal3 s -800 5720 800 5840 4 io_adr_i[5]
port 9 nsew signal input
rlabel metal3 s -800 6400 800 6520 4 io_adr_i[6]
port 10 nsew signal input
rlabel metal3 s -800 7080 800 7200 4 io_adr_i[7]
port 11 nsew signal input
rlabel metal3 s -800 7760 800 7880 4 io_adr_i[8]
port 12 nsew signal input
rlabel metal3 s -800 8576 800 8696 4 io_adr_i[9]
port 13 nsew signal input
rlabel metal2 s 17958 -800 18014 800 8 io_b_adr_i[0]
port 14 nsew signal output
rlabel metal2 s 19246 -800 19302 800 8 io_b_adr_i[1]
port 15 nsew signal output
rlabel metal2 s 1950 -800 2006 800 8 io_b_cs_i_0
port 16 nsew signal output
rlabel metal2 s 3238 -800 3294 800 8 io_b_cs_i_1
port 17 nsew signal output
rlabel metal2 s 15290 -800 15346 800 8 io_b_cs_i_10
port 18 nsew signal output
rlabel metal2 s 4618 -800 4674 800 8 io_b_cs_i_2
port 19 nsew signal output
rlabel metal2 s 5906 -800 5962 800 8 io_b_cs_i_3
port 20 nsew signal output
rlabel metal2 s 7286 -800 7342 800 8 io_b_cs_i_4
port 21 nsew signal output
rlabel metal2 s 8574 -800 8630 800 8 io_b_cs_i_5
port 22 nsew signal output
rlabel metal2 s 9954 -800 10010 800 8 io_b_cs_i_6
port 23 nsew signal output
rlabel metal2 s 11242 -800 11298 800 8 io_b_cs_i_7
port 24 nsew signal output
rlabel metal2 s 12622 -800 12678 800 8 io_b_cs_i_8
port 25 nsew signal output
rlabel metal2 s 13910 -800 13966 800 8 io_b_cs_i_9
port 26 nsew signal output
rlabel metal2 s 20626 -800 20682 800 8 io_b_dat_i[0]
port 27 nsew signal output
rlabel metal2 s 33966 -800 34022 800 8 io_b_dat_i[10]
port 28 nsew signal output
rlabel metal2 s 35254 -800 35310 800 8 io_b_dat_i[11]
port 29 nsew signal output
rlabel metal2 s 36634 -800 36690 800 8 io_b_dat_i[12]
port 30 nsew signal output
rlabel metal2 s 37922 -800 37978 800 8 io_b_dat_i[13]
port 31 nsew signal output
rlabel metal2 s 39302 -800 39358 800 8 io_b_dat_i[14]
port 32 nsew signal output
rlabel metal2 s 40590 -800 40646 800 8 io_b_dat_i[15]
port 33 nsew signal output
rlabel metal2 s 21914 -800 21970 800 8 io_b_dat_i[1]
port 34 nsew signal output
rlabel metal2 s 23294 -800 23350 800 8 io_b_dat_i[2]
port 35 nsew signal output
rlabel metal2 s 24582 -800 24638 800 8 io_b_dat_i[3]
port 36 nsew signal output
rlabel metal2 s 25962 -800 26018 800 8 io_b_dat_i[4]
port 37 nsew signal output
rlabel metal2 s 27250 -800 27306 800 8 io_b_dat_i[5]
port 38 nsew signal output
rlabel metal2 s 28630 -800 28686 800 8 io_b_dat_i[6]
port 39 nsew signal output
rlabel metal2 s 29918 -800 29974 800 8 io_b_dat_i[7]
port 40 nsew signal output
rlabel metal2 s 31298 -800 31354 800 8 io_b_dat_i[8]
port 41 nsew signal output
rlabel metal2 s 32586 -800 32642 800 8 io_b_dat_i[9]
port 42 nsew signal output
rlabel metal2 s 110 55200 166 56800 6 io_b_dat_o_0[0]
port 43 nsew signal input
rlabel metal2 s 36726 55200 36782 56800 6 io_b_dat_o_0[10]
port 44 nsew signal input
rlabel metal2 s 40406 55200 40462 56800 6 io_b_dat_o_0[11]
port 45 nsew signal input
rlabel metal2 s 44086 55200 44142 56800 6 io_b_dat_o_0[12]
port 46 nsew signal input
rlabel metal2 s 47674 55200 47730 56800 6 io_b_dat_o_0[13]
port 47 nsew signal input
rlabel metal2 s 51354 55200 51410 56800 6 io_b_dat_o_0[14]
port 48 nsew signal input
rlabel metal2 s 55034 55200 55090 56800 6 io_b_dat_o_0[15]
port 49 nsew signal input
rlabel metal2 s 3698 55200 3754 56800 6 io_b_dat_o_0[1]
port 50 nsew signal input
rlabel metal2 s 7378 55200 7434 56800 6 io_b_dat_o_0[2]
port 51 nsew signal input
rlabel metal2 s 11058 55200 11114 56800 6 io_b_dat_o_0[3]
port 52 nsew signal input
rlabel metal2 s 14738 55200 14794 56800 6 io_b_dat_o_0[4]
port 53 nsew signal input
rlabel metal2 s 18418 55200 18474 56800 6 io_b_dat_o_0[5]
port 54 nsew signal input
rlabel metal2 s 22098 55200 22154 56800 6 io_b_dat_o_0[6]
port 55 nsew signal input
rlabel metal2 s 25686 55200 25742 56800 6 io_b_dat_o_0[7]
port 56 nsew signal input
rlabel metal2 s 29366 55200 29422 56800 6 io_b_dat_o_0[8]
port 57 nsew signal input
rlabel metal2 s 33046 55200 33102 56800 6 io_b_dat_o_0[9]
port 58 nsew signal input
rlabel metal2 s 3422 55200 3478 56800 6 io_b_dat_o_10[0]
port 59 nsew signal input
rlabel metal2 s 40038 55200 40094 56800 6 io_b_dat_o_10[10]
port 60 nsew signal input
rlabel metal2 s 43718 55200 43774 56800 6 io_b_dat_o_10[11]
port 61 nsew signal input
rlabel metal2 s 47398 55200 47454 56800 6 io_b_dat_o_10[12]
port 62 nsew signal input
rlabel metal2 s 51078 55200 51134 56800 6 io_b_dat_o_10[13]
port 63 nsew signal input
rlabel metal2 s 54758 55200 54814 56800 6 io_b_dat_o_10[14]
port 64 nsew signal input
rlabel metal2 s 58346 55200 58402 56800 6 io_b_dat_o_10[15]
port 65 nsew signal input
rlabel metal2 s 7102 55200 7158 56800 6 io_b_dat_o_10[1]
port 66 nsew signal input
rlabel metal2 s 10690 55200 10746 56800 6 io_b_dat_o_10[2]
port 67 nsew signal input
rlabel metal2 s 14370 55200 14426 56800 6 io_b_dat_o_10[3]
port 68 nsew signal input
rlabel metal2 s 18050 55200 18106 56800 6 io_b_dat_o_10[4]
port 69 nsew signal input
rlabel metal2 s 21730 55200 21786 56800 6 io_b_dat_o_10[5]
port 70 nsew signal input
rlabel metal2 s 25410 55200 25466 56800 6 io_b_dat_o_10[6]
port 71 nsew signal input
rlabel metal2 s 29090 55200 29146 56800 6 io_b_dat_o_10[7]
port 72 nsew signal input
rlabel metal2 s 32678 55200 32734 56800 6 io_b_dat_o_10[8]
port 73 nsew signal input
rlabel metal2 s 36358 55200 36414 56800 6 io_b_dat_o_10[9]
port 74 nsew signal input
rlabel metal2 s 386 55200 442 56800 6 io_b_dat_o_1[0]
port 75 nsew signal input
rlabel metal2 s 37094 55200 37150 56800 6 io_b_dat_o_1[10]
port 76 nsew signal input
rlabel metal2 s 40682 55200 40738 56800 6 io_b_dat_o_1[11]
port 77 nsew signal input
rlabel metal2 s 44362 55200 44418 56800 6 io_b_dat_o_1[12]
port 78 nsew signal input
rlabel metal2 s 48042 55200 48098 56800 6 io_b_dat_o_1[13]
port 79 nsew signal input
rlabel metal2 s 51722 55200 51778 56800 6 io_b_dat_o_1[14]
port 80 nsew signal input
rlabel metal2 s 55402 55200 55458 56800 6 io_b_dat_o_1[15]
port 81 nsew signal input
rlabel metal2 s 4066 55200 4122 56800 6 io_b_dat_o_1[1]
port 82 nsew signal input
rlabel metal2 s 7746 55200 7802 56800 6 io_b_dat_o_1[2]
port 83 nsew signal input
rlabel metal2 s 11426 55200 11482 56800 6 io_b_dat_o_1[3]
port 84 nsew signal input
rlabel metal2 s 15106 55200 15162 56800 6 io_b_dat_o_1[4]
port 85 nsew signal input
rlabel metal2 s 18694 55200 18750 56800 6 io_b_dat_o_1[5]
port 86 nsew signal input
rlabel metal2 s 22374 55200 22430 56800 6 io_b_dat_o_1[6]
port 87 nsew signal input
rlabel metal2 s 26054 55200 26110 56800 6 io_b_dat_o_1[7]
port 88 nsew signal input
rlabel metal2 s 29734 55200 29790 56800 6 io_b_dat_o_1[8]
port 89 nsew signal input
rlabel metal2 s 33414 55200 33470 56800 6 io_b_dat_o_1[9]
port 90 nsew signal input
rlabel metal2 s 754 55200 810 56800 6 io_b_dat_o_2[0]
port 91 nsew signal input
rlabel metal2 s 37370 55200 37426 56800 6 io_b_dat_o_2[10]
port 92 nsew signal input
rlabel metal2 s 41050 55200 41106 56800 6 io_b_dat_o_2[11]
port 93 nsew signal input
rlabel metal2 s 44730 55200 44786 56800 6 io_b_dat_o_2[12]
port 94 nsew signal input
rlabel metal2 s 48410 55200 48466 56800 6 io_b_dat_o_2[13]
port 95 nsew signal input
rlabel metal2 s 52090 55200 52146 56800 6 io_b_dat_o_2[14]
port 96 nsew signal input
rlabel metal2 s 55678 55200 55734 56800 6 io_b_dat_o_2[15]
port 97 nsew signal input
rlabel metal2 s 4434 55200 4490 56800 6 io_b_dat_o_2[1]
port 98 nsew signal input
rlabel metal2 s 8022 55200 8078 56800 6 io_b_dat_o_2[2]
port 99 nsew signal input
rlabel metal2 s 11702 55200 11758 56800 6 io_b_dat_o_2[3]
port 100 nsew signal input
rlabel metal2 s 15382 55200 15438 56800 6 io_b_dat_o_2[4]
port 101 nsew signal input
rlabel metal2 s 19062 55200 19118 56800 6 io_b_dat_o_2[5]
port 102 nsew signal input
rlabel metal2 s 22742 55200 22798 56800 6 io_b_dat_o_2[6]
port 103 nsew signal input
rlabel metal2 s 26422 55200 26478 56800 6 io_b_dat_o_2[7]
port 104 nsew signal input
rlabel metal2 s 30102 55200 30158 56800 6 io_b_dat_o_2[8]
port 105 nsew signal input
rlabel metal2 s 33690 55200 33746 56800 6 io_b_dat_o_2[9]
port 106 nsew signal input
rlabel metal2 s 1030 55200 1086 56800 6 io_b_dat_o_3[0]
port 107 nsew signal input
rlabel metal2 s 37738 55200 37794 56800 6 io_b_dat_o_3[10]
port 108 nsew signal input
rlabel metal2 s 41418 55200 41474 56800 6 io_b_dat_o_3[11]
port 109 nsew signal input
rlabel metal2 s 45098 55200 45154 56800 6 io_b_dat_o_3[12]
port 110 nsew signal input
rlabel metal2 s 48686 55200 48742 56800 6 io_b_dat_o_3[13]
port 111 nsew signal input
rlabel metal2 s 52366 55200 52422 56800 6 io_b_dat_o_3[14]
port 112 nsew signal input
rlabel metal2 s 56046 55200 56102 56800 6 io_b_dat_o_3[15]
port 113 nsew signal input
rlabel metal2 s 4710 55200 4766 56800 6 io_b_dat_o_3[1]
port 114 nsew signal input
rlabel metal2 s 8390 55200 8446 56800 6 io_b_dat_o_3[2]
port 115 nsew signal input
rlabel metal2 s 12070 55200 12126 56800 6 io_b_dat_o_3[3]
port 116 nsew signal input
rlabel metal2 s 15750 55200 15806 56800 6 io_b_dat_o_3[4]
port 117 nsew signal input
rlabel metal2 s 19430 55200 19486 56800 6 io_b_dat_o_3[5]
port 118 nsew signal input
rlabel metal2 s 23018 55200 23074 56800 6 io_b_dat_o_3[6]
port 119 nsew signal input
rlabel metal2 s 26698 55200 26754 56800 6 io_b_dat_o_3[7]
port 120 nsew signal input
rlabel metal2 s 30378 55200 30434 56800 6 io_b_dat_o_3[8]
port 121 nsew signal input
rlabel metal2 s 34058 55200 34114 56800 6 io_b_dat_o_3[9]
port 122 nsew signal input
rlabel metal2 s 1398 55200 1454 56800 6 io_b_dat_o_4[0]
port 123 nsew signal input
rlabel metal2 s 38014 55200 38070 56800 6 io_b_dat_o_4[10]
port 124 nsew signal input
rlabel metal2 s 41694 55200 41750 56800 6 io_b_dat_o_4[11]
port 125 nsew signal input
rlabel metal2 s 45374 55200 45430 56800 6 io_b_dat_o_4[12]
port 126 nsew signal input
rlabel metal2 s 49054 55200 49110 56800 6 io_b_dat_o_4[13]
port 127 nsew signal input
rlabel metal2 s 52734 55200 52790 56800 6 io_b_dat_o_4[14]
port 128 nsew signal input
rlabel metal2 s 56414 55200 56470 56800 6 io_b_dat_o_4[15]
port 129 nsew signal input
rlabel metal2 s 5078 55200 5134 56800 6 io_b_dat_o_4[1]
port 130 nsew signal input
rlabel metal2 s 8758 55200 8814 56800 6 io_b_dat_o_4[2]
port 131 nsew signal input
rlabel metal2 s 12438 55200 12494 56800 6 io_b_dat_o_4[3]
port 132 nsew signal input
rlabel metal2 s 16026 55200 16082 56800 6 io_b_dat_o_4[4]
port 133 nsew signal input
rlabel metal2 s 19706 55200 19762 56800 6 io_b_dat_o_4[5]
port 134 nsew signal input
rlabel metal2 s 23386 55200 23442 56800 6 io_b_dat_o_4[6]
port 135 nsew signal input
rlabel metal2 s 27066 55200 27122 56800 6 io_b_dat_o_4[7]
port 136 nsew signal input
rlabel metal2 s 30746 55200 30802 56800 6 io_b_dat_o_4[8]
port 137 nsew signal input
rlabel metal2 s 34426 55200 34482 56800 6 io_b_dat_o_4[9]
port 138 nsew signal input
rlabel metal2 s 1766 55200 1822 56800 6 io_b_dat_o_5[0]
port 139 nsew signal input
rlabel metal2 s 38382 55200 38438 56800 6 io_b_dat_o_5[10]
port 140 nsew signal input
rlabel metal2 s 42062 55200 42118 56800 6 io_b_dat_o_5[11]
port 141 nsew signal input
rlabel metal2 s 45742 55200 45798 56800 6 io_b_dat_o_5[12]
port 142 nsew signal input
rlabel metal2 s 49422 55200 49478 56800 6 io_b_dat_o_5[13]
port 143 nsew signal input
rlabel metal2 s 53010 55200 53066 56800 6 io_b_dat_o_5[14]
port 144 nsew signal input
rlabel metal2 s 56690 55200 56746 56800 6 io_b_dat_o_5[15]
port 145 nsew signal input
rlabel metal2 s 5354 55200 5410 56800 6 io_b_dat_o_5[1]
port 146 nsew signal input
rlabel metal2 s 9034 55200 9090 56800 6 io_b_dat_o_5[2]
port 147 nsew signal input
rlabel metal2 s 12714 55200 12770 56800 6 io_b_dat_o_5[3]
port 148 nsew signal input
rlabel metal2 s 16394 55200 16450 56800 6 io_b_dat_o_5[4]
port 149 nsew signal input
rlabel metal2 s 20074 55200 20130 56800 6 io_b_dat_o_5[5]
port 150 nsew signal input
rlabel metal2 s 23754 55200 23810 56800 6 io_b_dat_o_5[6]
port 151 nsew signal input
rlabel metal2 s 27434 55200 27490 56800 6 io_b_dat_o_5[7]
port 152 nsew signal input
rlabel metal2 s 31022 55200 31078 56800 6 io_b_dat_o_5[8]
port 153 nsew signal input
rlabel metal2 s 34702 55200 34758 56800 6 io_b_dat_o_5[9]
port 154 nsew signal input
rlabel metal2 s 2042 55200 2098 56800 6 io_b_dat_o_6[0]
port 155 nsew signal input
rlabel metal2 s 38750 55200 38806 56800 6 io_b_dat_o_6[10]
port 156 nsew signal input
rlabel metal2 s 42430 55200 42486 56800 6 io_b_dat_o_6[11]
port 157 nsew signal input
rlabel metal2 s 46018 55200 46074 56800 6 io_b_dat_o_6[12]
port 158 nsew signal input
rlabel metal2 s 49698 55200 49754 56800 6 io_b_dat_o_6[13]
port 159 nsew signal input
rlabel metal2 s 53378 55200 53434 56800 6 io_b_dat_o_6[14]
port 160 nsew signal input
rlabel metal2 s 57058 55200 57114 56800 6 io_b_dat_o_6[15]
port 161 nsew signal input
rlabel metal2 s 5722 55200 5778 56800 6 io_b_dat_o_6[1]
port 162 nsew signal input
rlabel metal2 s 9402 55200 9458 56800 6 io_b_dat_o_6[2]
port 163 nsew signal input
rlabel metal2 s 13082 55200 13138 56800 6 io_b_dat_o_6[3]
port 164 nsew signal input
rlabel metal2 s 16762 55200 16818 56800 6 io_b_dat_o_6[4]
port 165 nsew signal input
rlabel metal2 s 20350 55200 20406 56800 6 io_b_dat_o_6[5]
port 166 nsew signal input
rlabel metal2 s 24030 55200 24086 56800 6 io_b_dat_o_6[6]
port 167 nsew signal input
rlabel metal2 s 27710 55200 27766 56800 6 io_b_dat_o_6[7]
port 168 nsew signal input
rlabel metal2 s 31390 55200 31446 56800 6 io_b_dat_o_6[8]
port 169 nsew signal input
rlabel metal2 s 35070 55200 35126 56800 6 io_b_dat_o_6[9]
port 170 nsew signal input
rlabel metal2 s 2410 55200 2466 56800 6 io_b_dat_o_7[0]
port 171 nsew signal input
rlabel metal2 s 39026 55200 39082 56800 6 io_b_dat_o_7[10]
port 172 nsew signal input
rlabel metal2 s 42706 55200 42762 56800 6 io_b_dat_o_7[11]
port 173 nsew signal input
rlabel metal2 s 46386 55200 46442 56800 6 io_b_dat_o_7[12]
port 174 nsew signal input
rlabel metal2 s 50066 55200 50122 56800 6 io_b_dat_o_7[13]
port 175 nsew signal input
rlabel metal2 s 53746 55200 53802 56800 6 io_b_dat_o_7[14]
port 176 nsew signal input
rlabel metal2 s 57426 55200 57482 56800 6 io_b_dat_o_7[15]
port 177 nsew signal input
rlabel metal2 s 6090 55200 6146 56800 6 io_b_dat_o_7[1]
port 178 nsew signal input
rlabel metal2 s 9770 55200 9826 56800 6 io_b_dat_o_7[2]
port 179 nsew signal input
rlabel metal2 s 13358 55200 13414 56800 6 io_b_dat_o_7[3]
port 180 nsew signal input
rlabel metal2 s 17038 55200 17094 56800 6 io_b_dat_o_7[4]
port 181 nsew signal input
rlabel metal2 s 20718 55200 20774 56800 6 io_b_dat_o_7[5]
port 182 nsew signal input
rlabel metal2 s 24398 55200 24454 56800 6 io_b_dat_o_7[6]
port 183 nsew signal input
rlabel metal2 s 28078 55200 28134 56800 6 io_b_dat_o_7[7]
port 184 nsew signal input
rlabel metal2 s 31758 55200 31814 56800 6 io_b_dat_o_7[8]
port 185 nsew signal input
rlabel metal2 s 35346 55200 35402 56800 6 io_b_dat_o_7[9]
port 186 nsew signal input
rlabel metal2 s 2686 55200 2742 56800 6 io_b_dat_o_8[0]
port 187 nsew signal input
rlabel metal2 s 39394 55200 39450 56800 6 io_b_dat_o_8[10]
port 188 nsew signal input
rlabel metal2 s 43074 55200 43130 56800 6 io_b_dat_o_8[11]
port 189 nsew signal input
rlabel metal2 s 46754 55200 46810 56800 6 io_b_dat_o_8[12]
port 190 nsew signal input
rlabel metal2 s 50342 55200 50398 56800 6 io_b_dat_o_8[13]
port 191 nsew signal input
rlabel metal2 s 54022 55200 54078 56800 6 io_b_dat_o_8[14]
port 192 nsew signal input
rlabel metal2 s 57702 55200 57758 56800 6 io_b_dat_o_8[15]
port 193 nsew signal input
rlabel metal2 s 6366 55200 6422 56800 6 io_b_dat_o_8[1]
port 194 nsew signal input
rlabel metal2 s 10046 55200 10102 56800 6 io_b_dat_o_8[2]
port 195 nsew signal input
rlabel metal2 s 13726 55200 13782 56800 6 io_b_dat_o_8[3]
port 196 nsew signal input
rlabel metal2 s 17406 55200 17462 56800 6 io_b_dat_o_8[4]
port 197 nsew signal input
rlabel metal2 s 21086 55200 21142 56800 6 io_b_dat_o_8[5]
port 198 nsew signal input
rlabel metal2 s 24766 55200 24822 56800 6 io_b_dat_o_8[6]
port 199 nsew signal input
rlabel metal2 s 28354 55200 28410 56800 6 io_b_dat_o_8[7]
port 200 nsew signal input
rlabel metal2 s 32034 55200 32090 56800 6 io_b_dat_o_8[8]
port 201 nsew signal input
rlabel metal2 s 35714 55200 35770 56800 6 io_b_dat_o_8[9]
port 202 nsew signal input
rlabel metal2 s 3054 55200 3110 56800 6 io_b_dat_o_9[0]
port 203 nsew signal input
rlabel metal2 s 39762 55200 39818 56800 6 io_b_dat_o_9[10]
port 204 nsew signal input
rlabel metal2 s 43350 55200 43406 56800 6 io_b_dat_o_9[11]
port 205 nsew signal input
rlabel metal2 s 47030 55200 47086 56800 6 io_b_dat_o_9[12]
port 206 nsew signal input
rlabel metal2 s 50710 55200 50766 56800 6 io_b_dat_o_9[13]
port 207 nsew signal input
rlabel metal2 s 54390 55200 54446 56800 6 io_b_dat_o_9[14]
port 208 nsew signal input
rlabel metal2 s 58070 55200 58126 56800 6 io_b_dat_o_9[15]
port 209 nsew signal input
rlabel metal2 s 6734 55200 6790 56800 6 io_b_dat_o_9[1]
port 210 nsew signal input
rlabel metal2 s 10414 55200 10470 56800 6 io_b_dat_o_9[2]
port 211 nsew signal input
rlabel metal2 s 14094 55200 14150 56800 6 io_b_dat_o_9[3]
port 212 nsew signal input
rlabel metal2 s 17682 55200 17738 56800 6 io_b_dat_o_9[4]
port 213 nsew signal input
rlabel metal2 s 21362 55200 21418 56800 6 io_b_dat_o_9[5]
port 214 nsew signal input
rlabel metal2 s 25042 55200 25098 56800 6 io_b_dat_o_9[6]
port 215 nsew signal input
rlabel metal2 s 28722 55200 28778 56800 6 io_b_dat_o_9[7]
port 216 nsew signal input
rlabel metal2 s 32402 55200 32458 56800 6 io_b_dat_o_9[8]
port 217 nsew signal input
rlabel metal2 s 36082 55200 36138 56800 6 io_b_dat_o_9[9]
port 218 nsew signal input
rlabel metal2 s 16578 -800 16634 800 8 io_b_we_i
port 219 nsew signal output
rlabel metal3 s -800 280 800 400 4 io_cs_i
port 220 nsew signal input
rlabel metal3 s -800 10616 800 10736 4 io_dat_i[0]
port 221 nsew signal input
rlabel metal3 s -800 17552 800 17672 4 io_dat_i[10]
port 222 nsew signal input
rlabel metal3 s -800 18232 800 18352 4 io_dat_i[11]
port 223 nsew signal input
rlabel metal3 s -800 18912 800 19032 4 io_dat_i[12]
port 224 nsew signal input
rlabel metal3 s -800 19592 800 19712 4 io_dat_i[13]
port 225 nsew signal input
rlabel metal3 s -800 20272 800 20392 4 io_dat_i[14]
port 226 nsew signal input
rlabel metal3 s -800 20952 800 21072 4 io_dat_i[15]
port 227 nsew signal input
rlabel metal3 s -800 21632 800 21752 4 io_dat_i[16]
port 228 nsew signal input
rlabel metal3 s -800 22312 800 22432 4 io_dat_i[17]
port 229 nsew signal input
rlabel metal3 s -800 22992 800 23112 4 io_dat_i[18]
port 230 nsew signal input
rlabel metal3 s -800 23672 800 23792 4 io_dat_i[19]
port 231 nsew signal input
rlabel metal3 s -800 11296 800 11416 4 io_dat_i[1]
port 232 nsew signal input
rlabel metal3 s -800 24488 800 24608 4 io_dat_i[20]
port 233 nsew signal input
rlabel metal3 s -800 25168 800 25288 4 io_dat_i[21]
port 234 nsew signal input
rlabel metal3 s -800 25848 800 25968 4 io_dat_i[22]
port 235 nsew signal input
rlabel metal3 s -800 26528 800 26648 4 io_dat_i[23]
port 236 nsew signal input
rlabel metal3 s -800 27208 800 27328 4 io_dat_i[24]
port 237 nsew signal input
rlabel metal3 s -800 27888 800 28008 4 io_dat_i[25]
port 238 nsew signal input
rlabel metal3 s -800 28568 800 28688 4 io_dat_i[26]
port 239 nsew signal input
rlabel metal3 s -800 29248 800 29368 4 io_dat_i[27]
port 240 nsew signal input
rlabel metal3 s -800 29928 800 30048 4 io_dat_i[28]
port 241 nsew signal input
rlabel metal3 s -800 30608 800 30728 4 io_dat_i[29]
port 242 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 io_dat_i[2]
port 243 nsew signal input
rlabel metal3 s -800 31288 800 31408 4 io_dat_i[30]
port 244 nsew signal input
rlabel metal3 s -800 31968 800 32088 4 io_dat_i[31]
port 245 nsew signal input
rlabel metal3 s -800 12656 800 12776 4 io_dat_i[3]
port 246 nsew signal input
rlabel metal3 s -800 13336 800 13456 4 io_dat_i[4]
port 247 nsew signal input
rlabel metal3 s -800 14016 800 14136 4 io_dat_i[5]
port 248 nsew signal input
rlabel metal3 s -800 14696 800 14816 4 io_dat_i[6]
port 249 nsew signal input
rlabel metal3 s -800 15376 800 15496 4 io_dat_i[7]
port 250 nsew signal input
rlabel metal3 s -800 16056 800 16176 4 io_dat_i[8]
port 251 nsew signal input
rlabel metal3 s -800 16872 800 16992 4 io_dat_i[9]
port 252 nsew signal input
rlabel metal3 s -800 32784 800 32904 4 io_dat_o[0]
port 253 nsew signal output
rlabel metal3 s -800 39584 800 39704 4 io_dat_o[10]
port 254 nsew signal output
rlabel metal3 s -800 40400 800 40520 4 io_dat_o[11]
port 255 nsew signal output
rlabel metal3 s -800 41080 800 41200 4 io_dat_o[12]
port 256 nsew signal output
rlabel metal3 s -800 41760 800 41880 4 io_dat_o[13]
port 257 nsew signal output
rlabel metal3 s -800 42440 800 42560 4 io_dat_o[14]
port 258 nsew signal output
rlabel metal3 s -800 43120 800 43240 4 io_dat_o[15]
port 259 nsew signal output
rlabel metal3 s -800 43800 800 43920 4 io_dat_o[16]
port 260 nsew signal output
rlabel metal3 s -800 44480 800 44600 4 io_dat_o[17]
port 261 nsew signal output
rlabel metal3 s -800 45160 800 45280 4 io_dat_o[18]
port 262 nsew signal output
rlabel metal3 s -800 45840 800 45960 4 io_dat_o[19]
port 263 nsew signal output
rlabel metal3 s -800 33464 800 33584 4 io_dat_o[1]
port 264 nsew signal output
rlabel metal3 s -800 46520 800 46640 4 io_dat_o[20]
port 265 nsew signal output
rlabel metal3 s -800 47200 800 47320 4 io_dat_o[21]
port 266 nsew signal output
rlabel metal3 s -800 47880 800 48000 4 io_dat_o[22]
port 267 nsew signal output
rlabel metal3 s -800 48696 800 48816 4 io_dat_o[23]
port 268 nsew signal output
rlabel metal3 s -800 49376 800 49496 4 io_dat_o[24]
port 269 nsew signal output
rlabel metal3 s -800 50056 800 50176 4 io_dat_o[25]
port 270 nsew signal output
rlabel metal3 s -800 50736 800 50856 4 io_dat_o[26]
port 271 nsew signal output
rlabel metal3 s -800 51416 800 51536 4 io_dat_o[27]
port 272 nsew signal output
rlabel metal3 s -800 52096 800 52216 4 io_dat_o[28]
port 273 nsew signal output
rlabel metal3 s -800 52776 800 52896 4 io_dat_o[29]
port 274 nsew signal output
rlabel metal3 s -800 34144 800 34264 4 io_dat_o[2]
port 275 nsew signal output
rlabel metal3 s -800 53456 800 53576 4 io_dat_o[30]
port 276 nsew signal output
rlabel metal3 s -800 54136 800 54256 4 io_dat_o[31]
port 277 nsew signal output
rlabel metal3 s -800 34824 800 34944 4 io_dat_o[3]
port 278 nsew signal output
rlabel metal3 s -800 35504 800 35624 4 io_dat_o[4]
port 279 nsew signal output
rlabel metal3 s -800 36184 800 36304 4 io_dat_o[5]
port 280 nsew signal output
rlabel metal3 s -800 36864 800 36984 4 io_dat_o[6]
port 281 nsew signal output
rlabel metal3 s -800 37544 800 37664 4 io_dat_o[7]
port 282 nsew signal output
rlabel metal3 s -800 38224 800 38344 4 io_dat_o[8]
port 283 nsew signal output
rlabel metal3 s -800 38904 800 39024 4 io_dat_o[9]
port 284 nsew signal output
rlabel metal3 s 59200 416 60800 536 6 io_dataLastBlock[0]
port 285 nsew signal input
rlabel metal3 s 59200 8712 60800 8832 6 io_dataLastBlock[10]
port 286 nsew signal input
rlabel metal3 s 59200 9528 60800 9648 6 io_dataLastBlock[11]
port 287 nsew signal input
rlabel metal3 s 59200 10344 60800 10464 6 io_dataLastBlock[12]
port 288 nsew signal input
rlabel metal3 s 59200 11160 60800 11280 6 io_dataLastBlock[13]
port 289 nsew signal input
rlabel metal3 s 59200 12112 60800 12232 6 io_dataLastBlock[14]
port 290 nsew signal input
rlabel metal3 s 59200 12928 60800 13048 6 io_dataLastBlock[15]
port 291 nsew signal input
rlabel metal3 s 59200 13744 60800 13864 6 io_dataLastBlock[16]
port 292 nsew signal input
rlabel metal3 s 59200 14560 60800 14680 6 io_dataLastBlock[17]
port 293 nsew signal input
rlabel metal3 s 59200 15376 60800 15496 6 io_dataLastBlock[18]
port 294 nsew signal input
rlabel metal3 s 59200 16192 60800 16312 6 io_dataLastBlock[19]
port 295 nsew signal input
rlabel metal3 s 59200 1232 60800 1352 6 io_dataLastBlock[1]
port 296 nsew signal input
rlabel metal3 s 59200 17008 60800 17128 6 io_dataLastBlock[20]
port 297 nsew signal input
rlabel metal3 s 59200 17960 60800 18080 6 io_dataLastBlock[21]
port 298 nsew signal input
rlabel metal3 s 59200 18776 60800 18896 6 io_dataLastBlock[22]
port 299 nsew signal input
rlabel metal3 s 59200 19592 60800 19712 6 io_dataLastBlock[23]
port 300 nsew signal input
rlabel metal3 s 59200 20408 60800 20528 6 io_dataLastBlock[24]
port 301 nsew signal input
rlabel metal3 s 59200 21224 60800 21344 6 io_dataLastBlock[25]
port 302 nsew signal input
rlabel metal3 s 59200 22040 60800 22160 6 io_dataLastBlock[26]
port 303 nsew signal input
rlabel metal3 s 59200 22992 60800 23112 6 io_dataLastBlock[27]
port 304 nsew signal input
rlabel metal3 s 59200 23808 60800 23928 6 io_dataLastBlock[28]
port 305 nsew signal input
rlabel metal3 s 59200 24624 60800 24744 6 io_dataLastBlock[29]
port 306 nsew signal input
rlabel metal3 s 59200 2048 60800 2168 6 io_dataLastBlock[2]
port 307 nsew signal input
rlabel metal3 s 59200 25440 60800 25560 6 io_dataLastBlock[30]
port 308 nsew signal input
rlabel metal3 s 59200 26256 60800 26376 6 io_dataLastBlock[31]
port 309 nsew signal input
rlabel metal3 s 59200 27072 60800 27192 6 io_dataLastBlock[32]
port 310 nsew signal input
rlabel metal3 s 59200 27888 60800 28008 6 io_dataLastBlock[33]
port 311 nsew signal input
rlabel metal3 s 59200 28840 60800 28960 6 io_dataLastBlock[34]
port 312 nsew signal input
rlabel metal3 s 59200 29656 60800 29776 6 io_dataLastBlock[35]
port 313 nsew signal input
rlabel metal3 s 59200 30472 60800 30592 6 io_dataLastBlock[36]
port 314 nsew signal input
rlabel metal3 s 59200 31288 60800 31408 6 io_dataLastBlock[37]
port 315 nsew signal input
rlabel metal3 s 59200 32104 60800 32224 6 io_dataLastBlock[38]
port 316 nsew signal input
rlabel metal3 s 59200 32920 60800 33040 6 io_dataLastBlock[39]
port 317 nsew signal input
rlabel metal3 s 59200 2864 60800 2984 6 io_dataLastBlock[3]
port 318 nsew signal input
rlabel metal3 s 59200 33736 60800 33856 6 io_dataLastBlock[40]
port 319 nsew signal input
rlabel metal3 s 59200 34688 60800 34808 6 io_dataLastBlock[41]
port 320 nsew signal input
rlabel metal3 s 59200 35504 60800 35624 6 io_dataLastBlock[42]
port 321 nsew signal input
rlabel metal3 s 59200 36320 60800 36440 6 io_dataLastBlock[43]
port 322 nsew signal input
rlabel metal3 s 59200 37136 60800 37256 6 io_dataLastBlock[44]
port 323 nsew signal input
rlabel metal3 s 59200 37952 60800 38072 6 io_dataLastBlock[45]
port 324 nsew signal input
rlabel metal3 s 59200 38768 60800 38888 6 io_dataLastBlock[46]
port 325 nsew signal input
rlabel metal3 s 59200 39720 60800 39840 6 io_dataLastBlock[47]
port 326 nsew signal input
rlabel metal3 s 59200 40536 60800 40656 6 io_dataLastBlock[48]
port 327 nsew signal input
rlabel metal3 s 59200 41352 60800 41472 6 io_dataLastBlock[49]
port 328 nsew signal input
rlabel metal3 s 59200 3680 60800 3800 6 io_dataLastBlock[4]
port 329 nsew signal input
rlabel metal3 s 59200 42168 60800 42288 6 io_dataLastBlock[50]
port 330 nsew signal input
rlabel metal3 s 59200 42984 60800 43104 6 io_dataLastBlock[51]
port 331 nsew signal input
rlabel metal3 s 59200 43800 60800 43920 6 io_dataLastBlock[52]
port 332 nsew signal input
rlabel metal3 s 59200 44616 60800 44736 6 io_dataLastBlock[53]
port 333 nsew signal input
rlabel metal3 s 59200 45568 60800 45688 6 io_dataLastBlock[54]
port 334 nsew signal input
rlabel metal3 s 59200 46384 60800 46504 6 io_dataLastBlock[55]
port 335 nsew signal input
rlabel metal3 s 59200 47200 60800 47320 6 io_dataLastBlock[56]
port 336 nsew signal input
rlabel metal3 s 59200 48016 60800 48136 6 io_dataLastBlock[57]
port 337 nsew signal input
rlabel metal3 s 59200 48832 60800 48952 6 io_dataLastBlock[58]
port 338 nsew signal input
rlabel metal3 s 59200 49648 60800 49768 6 io_dataLastBlock[59]
port 339 nsew signal input
rlabel metal3 s 59200 4496 60800 4616 6 io_dataLastBlock[5]
port 340 nsew signal input
rlabel metal3 s 59200 50464 60800 50584 6 io_dataLastBlock[60]
port 341 nsew signal input
rlabel metal3 s 59200 51416 60800 51536 6 io_dataLastBlock[61]
port 342 nsew signal input
rlabel metal3 s 59200 52232 60800 52352 6 io_dataLastBlock[62]
port 343 nsew signal input
rlabel metal3 s 59200 53048 60800 53168 6 io_dataLastBlock[63]
port 344 nsew signal input
rlabel metal3 s 59200 5312 60800 5432 6 io_dataLastBlock[6]
port 345 nsew signal input
rlabel metal3 s 59200 6264 60800 6384 6 io_dataLastBlock[7]
port 346 nsew signal input
rlabel metal3 s 59200 7080 60800 7200 6 io_dataLastBlock[8]
port 347 nsew signal input
rlabel metal3 s 59200 7896 60800 8016 6 io_dataLastBlock[9]
port 348 nsew signal input
rlabel metal3 s 59200 53864 60800 53984 6 io_dsi_in[0]
port 349 nsew signal input
rlabel metal2 s 59082 55200 59138 56800 6 io_dsi_in[1]
port 350 nsew signal input
rlabel metal2 s 59358 55200 59414 56800 6 io_dsi_in[2]
port 351 nsew signal input
rlabel metal3 s 59200 54680 60800 54800 6 io_dsi_in[3]
port 352 nsew signal input
rlabel metal2 s 59726 55200 59782 56800 6 io_dsi_in[4]
port 353 nsew signal input
rlabel metal3 s -800 55496 800 55616 4 io_dsi_in[5]
port 354 nsew signal input
rlabel metal3 s 59200 55496 60800 55616 6 io_dsi_in[6]
port 355 nsew signal input
rlabel metal2 s 59266 -800 59322 800 8 io_dsi_in[7]
port 356 nsew signal input
rlabel metal2 s 662 -800 718 800 8 io_dsi_o
port 357 nsew signal output
rlabel metal2 s 57978 -800 58034 800 8 io_irq
port 358 nsew signal output
rlabel metal2 s 56598 -800 56654 800 8 io_sync_out
port 359 nsew signal output
rlabel metal2 s 41970 -800 42026 800 8 io_vout[0]
port 360 nsew signal output
rlabel metal2 s 55310 -800 55366 800 8 io_vout[10]
port 361 nsew signal output
rlabel metal2 s 43258 -800 43314 800 8 io_vout[1]
port 362 nsew signal output
rlabel metal2 s 44638 -800 44694 800 8 io_vout[2]
port 363 nsew signal output
rlabel metal2 s 45926 -800 45982 800 8 io_vout[3]
port 364 nsew signal output
rlabel metal2 s 47306 -800 47362 800 8 io_vout[4]
port 365 nsew signal output
rlabel metal2 s 48594 -800 48650 800 8 io_vout[5]
port 366 nsew signal output
rlabel metal2 s 49974 -800 50030 800 8 io_vout[6]
port 367 nsew signal output
rlabel metal2 s 51262 -800 51318 800 8 io_vout[7]
port 368 nsew signal output
rlabel metal2 s 52642 -800 52698 800 8 io_vout[8]
port 369 nsew signal output
rlabel metal2 s 53930 -800 53986 800 8 io_vout[9]
port 370 nsew signal output
rlabel metal3 s -800 1640 800 1760 4 io_we_i
port 371 nsew signal input
rlabel metal2 s 58714 55200 58770 56800 6 wb_clk_i
port 372 nsew signal input
rlabel metal3 s -800 54816 800 54936 4 wb_rst_i
port 373 nsew signal input
rlabel metal4 s 34928 2128 35248 53360 6 vccd1
port 374 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 53360 6 vccd1
port 375 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 53360 6 vssd1
port 376 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 53360 6 vssd1
port 377 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 56000
string LEFview TRUE
string GDS_FILE /project/openlane/cic_con/runs/cic_con/results/magic/cic_con.gds
string GDS_END 8119868
string GDS_START 373878
<< end >>

