magic
tech sky130A
magscale 1 2
timestamp 1624040984
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 658 2128 179294 117552
<< metal2 >>
rect 1306 119200 1362 120800
rect 3974 119200 4030 120800
rect 6734 119200 6790 120800
rect 9402 119200 9458 120800
rect 12162 119200 12218 120800
rect 14922 119200 14978 120800
rect 17590 119200 17646 120800
rect 20350 119200 20406 120800
rect 23110 119200 23166 120800
rect 25778 119200 25834 120800
rect 28538 119200 28594 120800
rect 31298 119200 31354 120800
rect 33966 119200 34022 120800
rect 36726 119200 36782 120800
rect 39486 119200 39542 120800
rect 42154 119200 42210 120800
rect 44914 119200 44970 120800
rect 47674 119200 47730 120800
rect 50342 119200 50398 120800
rect 53102 119200 53158 120800
rect 55862 119200 55918 120800
rect 58530 119200 58586 120800
rect 61290 119200 61346 120800
rect 63958 119200 64014 120800
rect 66718 119200 66774 120800
rect 69478 119200 69534 120800
rect 72146 119200 72202 120800
rect 74906 119200 74962 120800
rect 77666 119200 77722 120800
rect 80334 119200 80390 120800
rect 83094 119200 83150 120800
rect 85854 119200 85910 120800
rect 88522 119200 88578 120800
rect 91282 119200 91338 120800
rect 94042 119200 94098 120800
rect 96710 119200 96766 120800
rect 99470 119200 99526 120800
rect 102230 119200 102286 120800
rect 104898 119200 104954 120800
rect 107658 119200 107714 120800
rect 110418 119200 110474 120800
rect 113086 119200 113142 120800
rect 115846 119200 115902 120800
rect 118606 119200 118662 120800
rect 121274 119200 121330 120800
rect 124034 119200 124090 120800
rect 126702 119200 126758 120800
rect 129462 119200 129518 120800
rect 132222 119200 132278 120800
rect 134890 119200 134946 120800
rect 137650 119200 137706 120800
rect 140410 119200 140466 120800
rect 143078 119200 143134 120800
rect 145838 119200 145894 120800
rect 148598 119200 148654 120800
rect 151266 119200 151322 120800
rect 154026 119200 154082 120800
rect 156786 119200 156842 120800
rect 159454 119200 159510 120800
rect 162214 119200 162270 120800
rect 164974 119200 165030 120800
rect 167642 119200 167698 120800
rect 170402 119200 170458 120800
rect 173162 119200 173218 120800
rect 175830 119200 175886 120800
rect 178590 119200 178646 120800
rect 662 -800 718 800
rect 2042 -800 2098 800
rect 3422 -800 3478 800
rect 4802 -800 4858 800
rect 6274 -800 6330 800
rect 7654 -800 7710 800
rect 9034 -800 9090 800
rect 10506 -800 10562 800
rect 11886 -800 11942 800
rect 13266 -800 13322 800
rect 14646 -800 14702 800
rect 16118 -800 16174 800
rect 17498 -800 17554 800
rect 18878 -800 18934 800
rect 20350 -800 20406 800
rect 21730 -800 21786 800
rect 23110 -800 23166 800
rect 24490 -800 24546 800
rect 25962 -800 26018 800
rect 27342 -800 27398 800
rect 28722 -800 28778 800
rect 30194 -800 30250 800
rect 31574 -800 31630 800
rect 32954 -800 33010 800
rect 34334 -800 34390 800
rect 35806 -800 35862 800
rect 37186 -800 37242 800
rect 38566 -800 38622 800
rect 40038 -800 40094 800
rect 41418 -800 41474 800
rect 42798 -800 42854 800
rect 44178 -800 44234 800
rect 45650 -800 45706 800
rect 47030 -800 47086 800
rect 48410 -800 48466 800
rect 49882 -800 49938 800
rect 51262 -800 51318 800
rect 52642 -800 52698 800
rect 54022 -800 54078 800
rect 55494 -800 55550 800
rect 56874 -800 56930 800
rect 58254 -800 58310 800
rect 59726 -800 59782 800
rect 61106 -800 61162 800
rect 62486 -800 62542 800
rect 63958 -800 64014 800
rect 65338 -800 65394 800
rect 66718 -800 66774 800
rect 68098 -800 68154 800
rect 69570 -800 69626 800
rect 70950 -800 71006 800
rect 72330 -800 72386 800
rect 73802 -800 73858 800
rect 75182 -800 75238 800
rect 76562 -800 76618 800
rect 77942 -800 77998 800
rect 79414 -800 79470 800
rect 80794 -800 80850 800
rect 82174 -800 82230 800
rect 83646 -800 83702 800
rect 85026 -800 85082 800
rect 86406 -800 86462 800
rect 87786 -800 87842 800
rect 89258 -800 89314 800
rect 90638 -800 90694 800
rect 92018 -800 92074 800
rect 93490 -800 93546 800
rect 94870 -800 94926 800
rect 96250 -800 96306 800
rect 97630 -800 97686 800
rect 99102 -800 99158 800
rect 100482 -800 100538 800
rect 101862 -800 101918 800
rect 103334 -800 103390 800
rect 104714 -800 104770 800
rect 106094 -800 106150 800
rect 107474 -800 107530 800
rect 108946 -800 109002 800
rect 110326 -800 110382 800
rect 111706 -800 111762 800
rect 113178 -800 113234 800
rect 114558 -800 114614 800
rect 115938 -800 115994 800
rect 117318 -800 117374 800
rect 118790 -800 118846 800
rect 120170 -800 120226 800
rect 121550 -800 121606 800
rect 123022 -800 123078 800
rect 124402 -800 124458 800
rect 125782 -800 125838 800
rect 127254 -800 127310 800
rect 128634 -800 128690 800
rect 130014 -800 130070 800
rect 131394 -800 131450 800
rect 132866 -800 132922 800
rect 134246 -800 134302 800
rect 135626 -800 135682 800
rect 137098 -800 137154 800
rect 138478 -800 138534 800
rect 139858 -800 139914 800
rect 141238 -800 141294 800
rect 142710 -800 142766 800
rect 144090 -800 144146 800
rect 145470 -800 145526 800
rect 146942 -800 146998 800
rect 148322 -800 148378 800
rect 149702 -800 149758 800
rect 151082 -800 151138 800
rect 152554 -800 152610 800
rect 153934 -800 153990 800
rect 155314 -800 155370 800
rect 156786 -800 156842 800
rect 158166 -800 158222 800
rect 159546 -800 159602 800
rect 160926 -800 160982 800
rect 162398 -800 162454 800
rect 163778 -800 163834 800
rect 165158 -800 165214 800
rect 166630 -800 166686 800
rect 168010 -800 168066 800
rect 169390 -800 169446 800
rect 170770 -800 170826 800
rect 172242 -800 172298 800
rect 173622 -800 173678 800
rect 175002 -800 175058 800
rect 176474 -800 176530 800
rect 177854 -800 177910 800
rect 179234 -800 179290 800
<< obsm2 >>
rect 664 119144 1250 119200
rect 1418 119144 3918 119200
rect 4086 119144 6678 119200
rect 6846 119144 9346 119200
rect 9514 119144 12106 119200
rect 12274 119144 14866 119200
rect 15034 119144 17534 119200
rect 17702 119144 20294 119200
rect 20462 119144 23054 119200
rect 23222 119144 25722 119200
rect 25890 119144 28482 119200
rect 28650 119144 31242 119200
rect 31410 119144 33910 119200
rect 34078 119144 36670 119200
rect 36838 119144 39430 119200
rect 39598 119144 42098 119200
rect 42266 119144 44858 119200
rect 45026 119144 47618 119200
rect 47786 119144 50286 119200
rect 50454 119144 53046 119200
rect 53214 119144 55806 119200
rect 55974 119144 58474 119200
rect 58642 119144 61234 119200
rect 61402 119144 63902 119200
rect 64070 119144 66662 119200
rect 66830 119144 69422 119200
rect 69590 119144 72090 119200
rect 72258 119144 74850 119200
rect 75018 119144 77610 119200
rect 77778 119144 80278 119200
rect 80446 119144 83038 119200
rect 83206 119144 85798 119200
rect 85966 119144 88466 119200
rect 88634 119144 91226 119200
rect 91394 119144 93986 119200
rect 94154 119144 96654 119200
rect 96822 119144 99414 119200
rect 99582 119144 102174 119200
rect 102342 119144 104842 119200
rect 105010 119144 107602 119200
rect 107770 119144 110362 119200
rect 110530 119144 113030 119200
rect 113198 119144 115790 119200
rect 115958 119144 118550 119200
rect 118718 119144 121218 119200
rect 121386 119144 123978 119200
rect 124146 119144 126646 119200
rect 126814 119144 129406 119200
rect 129574 119144 132166 119200
rect 132334 119144 134834 119200
rect 135002 119144 137594 119200
rect 137762 119144 140354 119200
rect 140522 119144 143022 119200
rect 143190 119144 145782 119200
rect 145950 119144 148542 119200
rect 148710 119144 151210 119200
rect 151378 119144 153970 119200
rect 154138 119144 156730 119200
rect 156898 119144 159398 119200
rect 159566 119144 162158 119200
rect 162326 119144 164918 119200
rect 165086 119144 167586 119200
rect 167754 119144 170346 119200
rect 170514 119144 173106 119200
rect 173274 119144 175774 119200
rect 175942 119144 178534 119200
rect 178702 119144 179288 119200
rect 664 856 179288 119144
rect 774 800 1986 856
rect 2154 800 3366 856
rect 3534 800 4746 856
rect 4914 800 6218 856
rect 6386 800 7598 856
rect 7766 800 8978 856
rect 9146 800 10450 856
rect 10618 800 11830 856
rect 11998 800 13210 856
rect 13378 800 14590 856
rect 14758 800 16062 856
rect 16230 800 17442 856
rect 17610 800 18822 856
rect 18990 800 20294 856
rect 20462 800 21674 856
rect 21842 800 23054 856
rect 23222 800 24434 856
rect 24602 800 25906 856
rect 26074 800 27286 856
rect 27454 800 28666 856
rect 28834 800 30138 856
rect 30306 800 31518 856
rect 31686 800 32898 856
rect 33066 800 34278 856
rect 34446 800 35750 856
rect 35918 800 37130 856
rect 37298 800 38510 856
rect 38678 800 39982 856
rect 40150 800 41362 856
rect 41530 800 42742 856
rect 42910 800 44122 856
rect 44290 800 45594 856
rect 45762 800 46974 856
rect 47142 800 48354 856
rect 48522 800 49826 856
rect 49994 800 51206 856
rect 51374 800 52586 856
rect 52754 800 53966 856
rect 54134 800 55438 856
rect 55606 800 56818 856
rect 56986 800 58198 856
rect 58366 800 59670 856
rect 59838 800 61050 856
rect 61218 800 62430 856
rect 62598 800 63902 856
rect 64070 800 65282 856
rect 65450 800 66662 856
rect 66830 800 68042 856
rect 68210 800 69514 856
rect 69682 800 70894 856
rect 71062 800 72274 856
rect 72442 800 73746 856
rect 73914 800 75126 856
rect 75294 800 76506 856
rect 76674 800 77886 856
rect 78054 800 79358 856
rect 79526 800 80738 856
rect 80906 800 82118 856
rect 82286 800 83590 856
rect 83758 800 84970 856
rect 85138 800 86350 856
rect 86518 800 87730 856
rect 87898 800 89202 856
rect 89370 800 90582 856
rect 90750 800 91962 856
rect 92130 800 93434 856
rect 93602 800 94814 856
rect 94982 800 96194 856
rect 96362 800 97574 856
rect 97742 800 99046 856
rect 99214 800 100426 856
rect 100594 800 101806 856
rect 101974 800 103278 856
rect 103446 800 104658 856
rect 104826 800 106038 856
rect 106206 800 107418 856
rect 107586 800 108890 856
rect 109058 800 110270 856
rect 110438 800 111650 856
rect 111818 800 113122 856
rect 113290 800 114502 856
rect 114670 800 115882 856
rect 116050 800 117262 856
rect 117430 800 118734 856
rect 118902 800 120114 856
rect 120282 800 121494 856
rect 121662 800 122966 856
rect 123134 800 124346 856
rect 124514 800 125726 856
rect 125894 800 127198 856
rect 127366 800 128578 856
rect 128746 800 129958 856
rect 130126 800 131338 856
rect 131506 800 132810 856
rect 132978 800 134190 856
rect 134358 800 135570 856
rect 135738 800 137042 856
rect 137210 800 138422 856
rect 138590 800 139802 856
rect 139970 800 141182 856
rect 141350 800 142654 856
rect 142822 800 144034 856
rect 144202 800 145414 856
rect 145582 800 146886 856
rect 147054 800 148266 856
rect 148434 800 149646 856
rect 149814 800 151026 856
rect 151194 800 152498 856
rect 152666 800 153878 856
rect 154046 800 155258 856
rect 155426 800 156730 856
rect 156898 800 158110 856
rect 158278 800 159490 856
rect 159658 800 160870 856
rect 161038 800 162342 856
rect 162510 800 163722 856
rect 163890 800 165102 856
rect 165270 800 166574 856
rect 166742 800 167954 856
rect 168122 800 169334 856
rect 169502 800 170714 856
rect 170882 800 172186 856
rect 172354 800 173566 856
rect 173734 800 174946 856
rect 175114 800 176418 856
rect 176586 800 177798 856
rect 177966 800 179178 856
<< metal3 >>
rect -800 118872 800 118992
rect 179200 118872 180800 118992
rect -800 116968 800 117088
rect 179200 116968 180800 117088
rect -800 115064 800 115184
rect 179200 115064 180800 115184
rect -800 113160 800 113280
rect 179200 113160 180800 113280
rect -800 111392 800 111512
rect 179200 111392 180800 111512
rect -800 109488 800 109608
rect 179200 109488 180800 109608
rect -800 107584 800 107704
rect 179200 107584 180800 107704
rect -800 105680 800 105800
rect 179200 105680 180800 105800
rect -800 103776 800 103896
rect 179200 103776 180800 103896
rect -800 102008 800 102128
rect 179200 102008 180800 102128
rect -800 100104 800 100224
rect 179200 100104 180800 100224
rect -800 98200 800 98320
rect 179200 98200 180800 98320
rect -800 96296 800 96416
rect 179200 96296 180800 96416
rect -800 94528 800 94648
rect 179200 94528 180800 94648
rect -800 92624 800 92744
rect 179200 92624 180800 92744
rect -800 90720 800 90840
rect 179200 90720 180800 90840
rect -800 88816 800 88936
rect 179200 88816 180800 88936
rect -800 86912 800 87032
rect 179200 86912 180800 87032
rect -800 85144 800 85264
rect 179200 85144 180800 85264
rect -800 83240 800 83360
rect 179200 83240 180800 83360
rect -800 81336 800 81456
rect 179200 81336 180800 81456
rect -800 79432 800 79552
rect 179200 79432 180800 79552
rect -800 77664 800 77784
rect 179200 77664 180800 77784
rect -800 75760 800 75880
rect 179200 75760 180800 75880
rect -800 73856 800 73976
rect 179200 73856 180800 73976
rect -800 71952 800 72072
rect 179200 71952 180800 72072
rect -800 70048 800 70168
rect 179200 70048 180800 70168
rect -800 68280 800 68400
rect 179200 68280 180800 68400
rect -800 66376 800 66496
rect 179200 66376 180800 66496
rect -800 64472 800 64592
rect 179200 64472 180800 64592
rect -800 62568 800 62688
rect 179200 62568 180800 62688
rect -800 60800 800 60920
rect 179200 60800 180800 60920
rect -800 58896 800 59016
rect 179200 58896 180800 59016
rect -800 56992 800 57112
rect 179200 56992 180800 57112
rect -800 55088 800 55208
rect 179200 55088 180800 55208
rect -800 53184 800 53304
rect 179200 53184 180800 53304
rect -800 51416 800 51536
rect 179200 51416 180800 51536
rect -800 49512 800 49632
rect 179200 49512 180800 49632
rect -800 47608 800 47728
rect 179200 47608 180800 47728
rect -800 45704 800 45824
rect 179200 45704 180800 45824
rect -800 43800 800 43920
rect 179200 43800 180800 43920
rect -800 42032 800 42152
rect 179200 42032 180800 42152
rect -800 40128 800 40248
rect 179200 40128 180800 40248
rect -800 38224 800 38344
rect 179200 38224 180800 38344
rect -800 36320 800 36440
rect 179200 36320 180800 36440
rect -800 34552 800 34672
rect 179200 34552 180800 34672
rect -800 32648 800 32768
rect 179200 32648 180800 32768
rect -800 30744 800 30864
rect 179200 30744 180800 30864
rect -800 28840 800 28960
rect 179200 28840 180800 28960
rect -800 26936 800 27056
rect 179200 26936 180800 27056
rect -800 25168 800 25288
rect 179200 25168 180800 25288
rect -800 23264 800 23384
rect 179200 23264 180800 23384
rect -800 21360 800 21480
rect 179200 21360 180800 21480
rect -800 19456 800 19576
rect 179200 19456 180800 19576
rect -800 17688 800 17808
rect 179200 17688 180800 17808
rect -800 15784 800 15904
rect 179200 15784 180800 15904
rect -800 13880 800 14000
rect 179200 13880 180800 14000
rect -800 11976 800 12096
rect 179200 11976 180800 12096
rect -800 10072 800 10192
rect 179200 10072 180800 10192
rect -800 8304 800 8424
rect 179200 8304 180800 8424
rect -800 6400 800 6520
rect 179200 6400 180800 6520
rect -800 4496 800 4616
rect 179200 4496 180800 4616
rect -800 2592 800 2712
rect 179200 2592 180800 2712
rect -800 824 800 944
rect 179200 824 180800 944
<< obsm3 >>
rect 880 118792 179120 118965
rect 800 117168 179200 118792
rect 880 116888 179120 117168
rect 800 115264 179200 116888
rect 880 114984 179120 115264
rect 800 113360 179200 114984
rect 880 113080 179120 113360
rect 800 111592 179200 113080
rect 880 111312 179120 111592
rect 800 109688 179200 111312
rect 880 109408 179120 109688
rect 800 107784 179200 109408
rect 880 107504 179120 107784
rect 800 105880 179200 107504
rect 880 105600 179120 105880
rect 800 103976 179200 105600
rect 880 103696 179120 103976
rect 800 102208 179200 103696
rect 880 101928 179120 102208
rect 800 100304 179200 101928
rect 880 100024 179120 100304
rect 800 98400 179200 100024
rect 880 98120 179120 98400
rect 800 96496 179200 98120
rect 880 96216 179120 96496
rect 800 94728 179200 96216
rect 880 94448 179120 94728
rect 800 92824 179200 94448
rect 880 92544 179120 92824
rect 800 90920 179200 92544
rect 880 90640 179120 90920
rect 800 89016 179200 90640
rect 880 88736 179120 89016
rect 800 87112 179200 88736
rect 880 86832 179120 87112
rect 800 85344 179200 86832
rect 880 85064 179120 85344
rect 800 83440 179200 85064
rect 880 83160 179120 83440
rect 800 81536 179200 83160
rect 880 81256 179120 81536
rect 800 79632 179200 81256
rect 880 79352 179120 79632
rect 800 77864 179200 79352
rect 880 77584 179120 77864
rect 800 75960 179200 77584
rect 880 75680 179120 75960
rect 800 74056 179200 75680
rect 880 73776 179120 74056
rect 800 72152 179200 73776
rect 880 71872 179120 72152
rect 800 70248 179200 71872
rect 880 69968 179120 70248
rect 800 68480 179200 69968
rect 880 68200 179120 68480
rect 800 66576 179200 68200
rect 880 66296 179120 66576
rect 800 64672 179200 66296
rect 880 64392 179120 64672
rect 800 62768 179200 64392
rect 880 62488 179120 62768
rect 800 61000 179200 62488
rect 880 60720 179120 61000
rect 800 59096 179200 60720
rect 880 58816 179120 59096
rect 800 57192 179200 58816
rect 880 56912 179120 57192
rect 800 55288 179200 56912
rect 880 55008 179120 55288
rect 800 53384 179200 55008
rect 880 53104 179120 53384
rect 800 51616 179200 53104
rect 880 51336 179120 51616
rect 800 49712 179200 51336
rect 880 49432 179120 49712
rect 800 47808 179200 49432
rect 880 47528 179120 47808
rect 800 45904 179200 47528
rect 880 45624 179120 45904
rect 800 44000 179200 45624
rect 880 43720 179120 44000
rect 800 42232 179200 43720
rect 880 41952 179120 42232
rect 800 40328 179200 41952
rect 880 40048 179120 40328
rect 800 38424 179200 40048
rect 880 38144 179120 38424
rect 800 36520 179200 38144
rect 880 36240 179120 36520
rect 800 34752 179200 36240
rect 880 34472 179120 34752
rect 800 32848 179200 34472
rect 880 32568 179120 32848
rect 800 30944 179200 32568
rect 880 30664 179120 30944
rect 800 29040 179200 30664
rect 880 28760 179120 29040
rect 800 27136 179200 28760
rect 880 26856 179120 27136
rect 800 25368 179200 26856
rect 880 25088 179120 25368
rect 800 23464 179200 25088
rect 880 23184 179120 23464
rect 800 21560 179200 23184
rect 880 21280 179120 21560
rect 800 19656 179200 21280
rect 880 19376 179120 19656
rect 800 17888 179200 19376
rect 880 17608 179120 17888
rect 800 15984 179200 17608
rect 880 15704 179120 15984
rect 800 14080 179200 15704
rect 880 13800 179120 14080
rect 800 12176 179200 13800
rect 880 11896 179120 12176
rect 800 10272 179200 11896
rect 880 9992 179120 10272
rect 800 8504 179200 9992
rect 880 8224 179120 8504
rect 800 6600 179200 8224
rect 880 6320 179120 6600
rect 800 4696 179200 6320
rect 880 4416 179120 4696
rect 800 2792 179200 4416
rect 880 2512 179120 2792
rect 800 1024 179200 2512
rect 880 851 179120 1024
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< labels >>
rlabel metal2 s 6734 119200 6790 120800 6 ao_reg[0]
port 1 nsew signal output
rlabel metal2 s 33966 119200 34022 120800 6 ao_reg[10]
port 2 nsew signal output
rlabel metal2 s 36726 119200 36782 120800 6 ao_reg[11]
port 3 nsew signal output
rlabel metal2 s 39486 119200 39542 120800 6 ao_reg[12]
port 4 nsew signal output
rlabel metal2 s 42154 119200 42210 120800 6 ao_reg[13]
port 5 nsew signal output
rlabel metal2 s 44914 119200 44970 120800 6 ao_reg[14]
port 6 nsew signal output
rlabel metal2 s 47674 119200 47730 120800 6 ao_reg[15]
port 7 nsew signal output
rlabel metal2 s 50342 119200 50398 120800 6 ao_reg[16]
port 8 nsew signal output
rlabel metal2 s 53102 119200 53158 120800 6 ao_reg[17]
port 9 nsew signal output
rlabel metal2 s 55862 119200 55918 120800 6 ao_reg[18]
port 10 nsew signal output
rlabel metal2 s 58530 119200 58586 120800 6 ao_reg[19]
port 11 nsew signal output
rlabel metal2 s 9402 119200 9458 120800 6 ao_reg[1]
port 12 nsew signal output
rlabel metal2 s 61290 119200 61346 120800 6 ao_reg[20]
port 13 nsew signal output
rlabel metal2 s 63958 119200 64014 120800 6 ao_reg[21]
port 14 nsew signal output
rlabel metal2 s 66718 119200 66774 120800 6 ao_reg[22]
port 15 nsew signal output
rlabel metal2 s 69478 119200 69534 120800 6 ao_reg[23]
port 16 nsew signal output
rlabel metal2 s 72146 119200 72202 120800 6 ao_reg[24]
port 17 nsew signal output
rlabel metal2 s 74906 119200 74962 120800 6 ao_reg[25]
port 18 nsew signal output
rlabel metal2 s 77666 119200 77722 120800 6 ao_reg[26]
port 19 nsew signal output
rlabel metal2 s 80334 119200 80390 120800 6 ao_reg[27]
port 20 nsew signal output
rlabel metal2 s 83094 119200 83150 120800 6 ao_reg[28]
port 21 nsew signal output
rlabel metal2 s 85854 119200 85910 120800 6 ao_reg[29]
port 22 nsew signal output
rlabel metal2 s 12162 119200 12218 120800 6 ao_reg[2]
port 23 nsew signal output
rlabel metal2 s 88522 119200 88578 120800 6 ao_reg[30]
port 24 nsew signal output
rlabel metal2 s 91282 119200 91338 120800 6 ao_reg[31]
port 25 nsew signal output
rlabel metal2 s 14922 119200 14978 120800 6 ao_reg[3]
port 26 nsew signal output
rlabel metal2 s 17590 119200 17646 120800 6 ao_reg[4]
port 27 nsew signal output
rlabel metal2 s 20350 119200 20406 120800 6 ao_reg[5]
port 28 nsew signal output
rlabel metal2 s 23110 119200 23166 120800 6 ao_reg[6]
port 29 nsew signal output
rlabel metal2 s 25778 119200 25834 120800 6 ao_reg[7]
port 30 nsew signal output
rlabel metal2 s 28538 119200 28594 120800 6 ao_reg[8]
port 31 nsew signal output
rlabel metal2 s 31298 119200 31354 120800 6 ao_reg[9]
port 32 nsew signal output
rlabel metal2 s 3974 119200 4030 120800 6 asel
port 33 nsew signal input
rlabel metal2 s 94042 119200 94098 120800 6 bo_reg[0]
port 34 nsew signal output
rlabel metal2 s 121274 119200 121330 120800 6 bo_reg[10]
port 35 nsew signal output
rlabel metal2 s 124034 119200 124090 120800 6 bo_reg[11]
port 36 nsew signal output
rlabel metal2 s 126702 119200 126758 120800 6 bo_reg[12]
port 37 nsew signal output
rlabel metal2 s 129462 119200 129518 120800 6 bo_reg[13]
port 38 nsew signal output
rlabel metal2 s 132222 119200 132278 120800 6 bo_reg[14]
port 39 nsew signal output
rlabel metal2 s 134890 119200 134946 120800 6 bo_reg[15]
port 40 nsew signal output
rlabel metal2 s 137650 119200 137706 120800 6 bo_reg[16]
port 41 nsew signal output
rlabel metal2 s 140410 119200 140466 120800 6 bo_reg[17]
port 42 nsew signal output
rlabel metal2 s 143078 119200 143134 120800 6 bo_reg[18]
port 43 nsew signal output
rlabel metal2 s 145838 119200 145894 120800 6 bo_reg[19]
port 44 nsew signal output
rlabel metal2 s 96710 119200 96766 120800 6 bo_reg[1]
port 45 nsew signal output
rlabel metal2 s 148598 119200 148654 120800 6 bo_reg[20]
port 46 nsew signal output
rlabel metal2 s 151266 119200 151322 120800 6 bo_reg[21]
port 47 nsew signal output
rlabel metal2 s 154026 119200 154082 120800 6 bo_reg[22]
port 48 nsew signal output
rlabel metal2 s 156786 119200 156842 120800 6 bo_reg[23]
port 49 nsew signal output
rlabel metal2 s 159454 119200 159510 120800 6 bo_reg[24]
port 50 nsew signal output
rlabel metal2 s 162214 119200 162270 120800 6 bo_reg[25]
port 51 nsew signal output
rlabel metal2 s 164974 119200 165030 120800 6 bo_reg[26]
port 52 nsew signal output
rlabel metal2 s 167642 119200 167698 120800 6 bo_reg[27]
port 53 nsew signal output
rlabel metal2 s 170402 119200 170458 120800 6 bo_reg[28]
port 54 nsew signal output
rlabel metal2 s 173162 119200 173218 120800 6 bo_reg[29]
port 55 nsew signal output
rlabel metal2 s 99470 119200 99526 120800 6 bo_reg[2]
port 56 nsew signal output
rlabel metal2 s 175830 119200 175886 120800 6 bo_reg[30]
port 57 nsew signal output
rlabel metal2 s 178590 119200 178646 120800 6 bo_reg[31]
port 58 nsew signal output
rlabel metal2 s 102230 119200 102286 120800 6 bo_reg[3]
port 59 nsew signal output
rlabel metal2 s 104898 119200 104954 120800 6 bo_reg[4]
port 60 nsew signal output
rlabel metal2 s 107658 119200 107714 120800 6 bo_reg[5]
port 61 nsew signal output
rlabel metal2 s 110418 119200 110474 120800 6 bo_reg[6]
port 62 nsew signal output
rlabel metal2 s 113086 119200 113142 120800 6 bo_reg[7]
port 63 nsew signal output
rlabel metal2 s 115846 119200 115902 120800 6 bo_reg[8]
port 64 nsew signal output
rlabel metal2 s 118606 119200 118662 120800 6 bo_reg[9]
port 65 nsew signal output
rlabel metal2 s 1306 119200 1362 120800 6 clk
port 66 nsew signal input
rlabel metal3 s 179200 824 180800 944 6 e_i[0]
port 67 nsew signal input
rlabel metal3 s 179200 38224 180800 38344 6 e_i[10]
port 68 nsew signal input
rlabel metal3 s 179200 42032 180800 42152 6 e_i[11]
port 69 nsew signal input
rlabel metal3 s 179200 45704 180800 45824 6 e_i[12]
port 70 nsew signal input
rlabel metal3 s 179200 49512 180800 49632 6 e_i[13]
port 71 nsew signal input
rlabel metal3 s 179200 53184 180800 53304 6 e_i[14]
port 72 nsew signal input
rlabel metal3 s 179200 56992 180800 57112 6 e_i[15]
port 73 nsew signal input
rlabel metal3 s 179200 60800 180800 60920 6 e_i[16]
port 74 nsew signal input
rlabel metal3 s 179200 64472 180800 64592 6 e_i[17]
port 75 nsew signal input
rlabel metal3 s 179200 68280 180800 68400 6 e_i[18]
port 76 nsew signal input
rlabel metal3 s 179200 71952 180800 72072 6 e_i[19]
port 77 nsew signal input
rlabel metal3 s 179200 4496 180800 4616 6 e_i[1]
port 78 nsew signal input
rlabel metal3 s 179200 75760 180800 75880 6 e_i[20]
port 79 nsew signal input
rlabel metal3 s 179200 79432 180800 79552 6 e_i[21]
port 80 nsew signal input
rlabel metal3 s 179200 83240 180800 83360 6 e_i[22]
port 81 nsew signal input
rlabel metal3 s 179200 86912 180800 87032 6 e_i[23]
port 82 nsew signal input
rlabel metal3 s 179200 90720 180800 90840 6 e_i[24]
port 83 nsew signal input
rlabel metal3 s 179200 94528 180800 94648 6 e_i[25]
port 84 nsew signal input
rlabel metal3 s 179200 98200 180800 98320 6 e_i[26]
port 85 nsew signal input
rlabel metal3 s 179200 102008 180800 102128 6 e_i[27]
port 86 nsew signal input
rlabel metal3 s 179200 105680 180800 105800 6 e_i[28]
port 87 nsew signal input
rlabel metal3 s 179200 109488 180800 109608 6 e_i[29]
port 88 nsew signal input
rlabel metal3 s 179200 8304 180800 8424 6 e_i[2]
port 89 nsew signal input
rlabel metal3 s 179200 113160 180800 113280 6 e_i[30]
port 90 nsew signal input
rlabel metal3 s 179200 116968 180800 117088 6 e_i[31]
port 91 nsew signal input
rlabel metal3 s 179200 11976 180800 12096 6 e_i[3]
port 92 nsew signal input
rlabel metal3 s 179200 15784 180800 15904 6 e_i[4]
port 93 nsew signal input
rlabel metal3 s 179200 19456 180800 19576 6 e_i[5]
port 94 nsew signal input
rlabel metal3 s 179200 23264 180800 23384 6 e_i[6]
port 95 nsew signal input
rlabel metal3 s 179200 26936 180800 27056 6 e_i[7]
port 96 nsew signal input
rlabel metal3 s 179200 30744 180800 30864 6 e_i[8]
port 97 nsew signal input
rlabel metal3 s 179200 34552 180800 34672 6 e_i[9]
port 98 nsew signal input
rlabel metal3 s 179200 2592 180800 2712 6 e_o[0]
port 99 nsew signal output
rlabel metal3 s 179200 40128 180800 40248 6 e_o[10]
port 100 nsew signal output
rlabel metal3 s 179200 43800 180800 43920 6 e_o[11]
port 101 nsew signal output
rlabel metal3 s 179200 47608 180800 47728 6 e_o[12]
port 102 nsew signal output
rlabel metal3 s 179200 51416 180800 51536 6 e_o[13]
port 103 nsew signal output
rlabel metal3 s 179200 55088 180800 55208 6 e_o[14]
port 104 nsew signal output
rlabel metal3 s 179200 58896 180800 59016 6 e_o[15]
port 105 nsew signal output
rlabel metal3 s 179200 62568 180800 62688 6 e_o[16]
port 106 nsew signal output
rlabel metal3 s 179200 66376 180800 66496 6 e_o[17]
port 107 nsew signal output
rlabel metal3 s 179200 70048 180800 70168 6 e_o[18]
port 108 nsew signal output
rlabel metal3 s 179200 73856 180800 73976 6 e_o[19]
port 109 nsew signal output
rlabel metal3 s 179200 6400 180800 6520 6 e_o[1]
port 110 nsew signal output
rlabel metal3 s 179200 77664 180800 77784 6 e_o[20]
port 111 nsew signal output
rlabel metal3 s 179200 81336 180800 81456 6 e_o[21]
port 112 nsew signal output
rlabel metal3 s 179200 85144 180800 85264 6 e_o[22]
port 113 nsew signal output
rlabel metal3 s 179200 88816 180800 88936 6 e_o[23]
port 114 nsew signal output
rlabel metal3 s 179200 92624 180800 92744 6 e_o[24]
port 115 nsew signal output
rlabel metal3 s 179200 96296 180800 96416 6 e_o[25]
port 116 nsew signal output
rlabel metal3 s 179200 100104 180800 100224 6 e_o[26]
port 117 nsew signal output
rlabel metal3 s 179200 103776 180800 103896 6 e_o[27]
port 118 nsew signal output
rlabel metal3 s 179200 107584 180800 107704 6 e_o[28]
port 119 nsew signal output
rlabel metal3 s 179200 111392 180800 111512 6 e_o[29]
port 120 nsew signal output
rlabel metal3 s 179200 10072 180800 10192 6 e_o[2]
port 121 nsew signal output
rlabel metal3 s 179200 115064 180800 115184 6 e_o[30]
port 122 nsew signal output
rlabel metal3 s 179200 118872 180800 118992 6 e_o[31]
port 123 nsew signal output
rlabel metal3 s 179200 13880 180800 14000 6 e_o[3]
port 124 nsew signal output
rlabel metal3 s 179200 17688 180800 17808 6 e_o[4]
port 125 nsew signal output
rlabel metal3 s 179200 21360 180800 21480 6 e_o[5]
port 126 nsew signal output
rlabel metal3 s 179200 25168 180800 25288 6 e_o[6]
port 127 nsew signal output
rlabel metal3 s 179200 28840 180800 28960 6 e_o[7]
port 128 nsew signal output
rlabel metal3 s 179200 32648 180800 32768 6 e_o[8]
port 129 nsew signal output
rlabel metal3 s 179200 36320 180800 36440 6 e_o[9]
port 130 nsew signal output
rlabel metal2 s 90638 -800 90694 800 8 se_i[0]
port 131 nsew signal input
rlabel metal2 s 118790 -800 118846 800 8 se_i[10]
port 132 nsew signal input
rlabel metal2 s 121550 -800 121606 800 8 se_i[11]
port 133 nsew signal input
rlabel metal2 s 124402 -800 124458 800 8 se_i[12]
port 134 nsew signal input
rlabel metal2 s 127254 -800 127310 800 8 se_i[13]
port 135 nsew signal input
rlabel metal2 s 130014 -800 130070 800 8 se_i[14]
port 136 nsew signal input
rlabel metal2 s 132866 -800 132922 800 8 se_i[15]
port 137 nsew signal input
rlabel metal2 s 135626 -800 135682 800 8 se_i[16]
port 138 nsew signal input
rlabel metal2 s 138478 -800 138534 800 8 se_i[17]
port 139 nsew signal input
rlabel metal2 s 141238 -800 141294 800 8 se_i[18]
port 140 nsew signal input
rlabel metal2 s 144090 -800 144146 800 8 se_i[19]
port 141 nsew signal input
rlabel metal2 s 93490 -800 93546 800 8 se_i[1]
port 142 nsew signal input
rlabel metal2 s 146942 -800 146998 800 8 se_i[20]
port 143 nsew signal input
rlabel metal2 s 149702 -800 149758 800 8 se_i[21]
port 144 nsew signal input
rlabel metal2 s 152554 -800 152610 800 8 se_i[22]
port 145 nsew signal input
rlabel metal2 s 155314 -800 155370 800 8 se_i[23]
port 146 nsew signal input
rlabel metal2 s 158166 -800 158222 800 8 se_i[24]
port 147 nsew signal input
rlabel metal2 s 160926 -800 160982 800 8 se_i[25]
port 148 nsew signal input
rlabel metal2 s 163778 -800 163834 800 8 se_i[26]
port 149 nsew signal input
rlabel metal2 s 166630 -800 166686 800 8 se_i[27]
port 150 nsew signal input
rlabel metal2 s 169390 -800 169446 800 8 se_i[28]
port 151 nsew signal input
rlabel metal2 s 172242 -800 172298 800 8 se_i[29]
port 152 nsew signal input
rlabel metal2 s 96250 -800 96306 800 8 se_i[2]
port 153 nsew signal input
rlabel metal2 s 175002 -800 175058 800 8 se_i[30]
port 154 nsew signal input
rlabel metal2 s 177854 -800 177910 800 8 se_i[31]
port 155 nsew signal input
rlabel metal2 s 99102 -800 99158 800 8 se_i[3]
port 156 nsew signal input
rlabel metal2 s 101862 -800 101918 800 8 se_i[4]
port 157 nsew signal input
rlabel metal2 s 104714 -800 104770 800 8 se_i[5]
port 158 nsew signal input
rlabel metal2 s 107474 -800 107530 800 8 se_i[6]
port 159 nsew signal input
rlabel metal2 s 110326 -800 110382 800 8 se_i[7]
port 160 nsew signal input
rlabel metal2 s 113178 -800 113234 800 8 se_i[8]
port 161 nsew signal input
rlabel metal2 s 115938 -800 115994 800 8 se_i[9]
port 162 nsew signal input
rlabel metal2 s 92018 -800 92074 800 8 se_o[0]
port 163 nsew signal output
rlabel metal2 s 120170 -800 120226 800 8 se_o[10]
port 164 nsew signal output
rlabel metal2 s 123022 -800 123078 800 8 se_o[11]
port 165 nsew signal output
rlabel metal2 s 125782 -800 125838 800 8 se_o[12]
port 166 nsew signal output
rlabel metal2 s 128634 -800 128690 800 8 se_o[13]
port 167 nsew signal output
rlabel metal2 s 131394 -800 131450 800 8 se_o[14]
port 168 nsew signal output
rlabel metal2 s 134246 -800 134302 800 8 se_o[15]
port 169 nsew signal output
rlabel metal2 s 137098 -800 137154 800 8 se_o[16]
port 170 nsew signal output
rlabel metal2 s 139858 -800 139914 800 8 se_o[17]
port 171 nsew signal output
rlabel metal2 s 142710 -800 142766 800 8 se_o[18]
port 172 nsew signal output
rlabel metal2 s 145470 -800 145526 800 8 se_o[19]
port 173 nsew signal output
rlabel metal2 s 94870 -800 94926 800 8 se_o[1]
port 174 nsew signal output
rlabel metal2 s 148322 -800 148378 800 8 se_o[20]
port 175 nsew signal output
rlabel metal2 s 151082 -800 151138 800 8 se_o[21]
port 176 nsew signal output
rlabel metal2 s 153934 -800 153990 800 8 se_o[22]
port 177 nsew signal output
rlabel metal2 s 156786 -800 156842 800 8 se_o[23]
port 178 nsew signal output
rlabel metal2 s 159546 -800 159602 800 8 se_o[24]
port 179 nsew signal output
rlabel metal2 s 162398 -800 162454 800 8 se_o[25]
port 180 nsew signal output
rlabel metal2 s 165158 -800 165214 800 8 se_o[26]
port 181 nsew signal output
rlabel metal2 s 168010 -800 168066 800 8 se_o[27]
port 182 nsew signal output
rlabel metal2 s 170770 -800 170826 800 8 se_o[28]
port 183 nsew signal output
rlabel metal2 s 173622 -800 173678 800 8 se_o[29]
port 184 nsew signal output
rlabel metal2 s 97630 -800 97686 800 8 se_o[2]
port 185 nsew signal output
rlabel metal2 s 176474 -800 176530 800 8 se_o[30]
port 186 nsew signal output
rlabel metal2 s 179234 -800 179290 800 8 se_o[31]
port 187 nsew signal output
rlabel metal2 s 100482 -800 100538 800 8 se_o[3]
port 188 nsew signal output
rlabel metal2 s 103334 -800 103390 800 8 se_o[4]
port 189 nsew signal output
rlabel metal2 s 106094 -800 106150 800 8 se_o[5]
port 190 nsew signal output
rlabel metal2 s 108946 -800 109002 800 8 se_o[6]
port 191 nsew signal output
rlabel metal2 s 111706 -800 111762 800 8 se_o[7]
port 192 nsew signal output
rlabel metal2 s 114558 -800 114614 800 8 se_o[8]
port 193 nsew signal output
rlabel metal2 s 117318 -800 117374 800 8 se_o[9]
port 194 nsew signal output
rlabel metal2 s 662 -800 718 800 8 sw_i[0]
port 195 nsew signal input
rlabel metal2 s 28722 -800 28778 800 8 sw_i[10]
port 196 nsew signal input
rlabel metal2 s 31574 -800 31630 800 8 sw_i[11]
port 197 nsew signal input
rlabel metal2 s 34334 -800 34390 800 8 sw_i[12]
port 198 nsew signal input
rlabel metal2 s 37186 -800 37242 800 8 sw_i[13]
port 199 nsew signal input
rlabel metal2 s 40038 -800 40094 800 8 sw_i[14]
port 200 nsew signal input
rlabel metal2 s 42798 -800 42854 800 8 sw_i[15]
port 201 nsew signal input
rlabel metal2 s 45650 -800 45706 800 8 sw_i[16]
port 202 nsew signal input
rlabel metal2 s 48410 -800 48466 800 8 sw_i[17]
port 203 nsew signal input
rlabel metal2 s 51262 -800 51318 800 8 sw_i[18]
port 204 nsew signal input
rlabel metal2 s 54022 -800 54078 800 8 sw_i[19]
port 205 nsew signal input
rlabel metal2 s 3422 -800 3478 800 8 sw_i[1]
port 206 nsew signal input
rlabel metal2 s 56874 -800 56930 800 8 sw_i[20]
port 207 nsew signal input
rlabel metal2 s 59726 -800 59782 800 8 sw_i[21]
port 208 nsew signal input
rlabel metal2 s 62486 -800 62542 800 8 sw_i[22]
port 209 nsew signal input
rlabel metal2 s 65338 -800 65394 800 8 sw_i[23]
port 210 nsew signal input
rlabel metal2 s 68098 -800 68154 800 8 sw_i[24]
port 211 nsew signal input
rlabel metal2 s 70950 -800 71006 800 8 sw_i[25]
port 212 nsew signal input
rlabel metal2 s 73802 -800 73858 800 8 sw_i[26]
port 213 nsew signal input
rlabel metal2 s 76562 -800 76618 800 8 sw_i[27]
port 214 nsew signal input
rlabel metal2 s 79414 -800 79470 800 8 sw_i[28]
port 215 nsew signal input
rlabel metal2 s 82174 -800 82230 800 8 sw_i[29]
port 216 nsew signal input
rlabel metal2 s 6274 -800 6330 800 8 sw_i[2]
port 217 nsew signal input
rlabel metal2 s 85026 -800 85082 800 8 sw_i[30]
port 218 nsew signal input
rlabel metal2 s 87786 -800 87842 800 8 sw_i[31]
port 219 nsew signal input
rlabel metal2 s 9034 -800 9090 800 8 sw_i[3]
port 220 nsew signal input
rlabel metal2 s 11886 -800 11942 800 8 sw_i[4]
port 221 nsew signal input
rlabel metal2 s 14646 -800 14702 800 8 sw_i[5]
port 222 nsew signal input
rlabel metal2 s 17498 -800 17554 800 8 sw_i[6]
port 223 nsew signal input
rlabel metal2 s 20350 -800 20406 800 8 sw_i[7]
port 224 nsew signal input
rlabel metal2 s 23110 -800 23166 800 8 sw_i[8]
port 225 nsew signal input
rlabel metal2 s 25962 -800 26018 800 8 sw_i[9]
port 226 nsew signal input
rlabel metal2 s 2042 -800 2098 800 8 sw_o[0]
port 227 nsew signal output
rlabel metal2 s 30194 -800 30250 800 8 sw_o[10]
port 228 nsew signal output
rlabel metal2 s 32954 -800 33010 800 8 sw_o[11]
port 229 nsew signal output
rlabel metal2 s 35806 -800 35862 800 8 sw_o[12]
port 230 nsew signal output
rlabel metal2 s 38566 -800 38622 800 8 sw_o[13]
port 231 nsew signal output
rlabel metal2 s 41418 -800 41474 800 8 sw_o[14]
port 232 nsew signal output
rlabel metal2 s 44178 -800 44234 800 8 sw_o[15]
port 233 nsew signal output
rlabel metal2 s 47030 -800 47086 800 8 sw_o[16]
port 234 nsew signal output
rlabel metal2 s 49882 -800 49938 800 8 sw_o[17]
port 235 nsew signal output
rlabel metal2 s 52642 -800 52698 800 8 sw_o[18]
port 236 nsew signal output
rlabel metal2 s 55494 -800 55550 800 8 sw_o[19]
port 237 nsew signal output
rlabel metal2 s 4802 -800 4858 800 8 sw_o[1]
port 238 nsew signal output
rlabel metal2 s 58254 -800 58310 800 8 sw_o[20]
port 239 nsew signal output
rlabel metal2 s 61106 -800 61162 800 8 sw_o[21]
port 240 nsew signal output
rlabel metal2 s 63958 -800 64014 800 8 sw_o[22]
port 241 nsew signal output
rlabel metal2 s 66718 -800 66774 800 8 sw_o[23]
port 242 nsew signal output
rlabel metal2 s 69570 -800 69626 800 8 sw_o[24]
port 243 nsew signal output
rlabel metal2 s 72330 -800 72386 800 8 sw_o[25]
port 244 nsew signal output
rlabel metal2 s 75182 -800 75238 800 8 sw_o[26]
port 245 nsew signal output
rlabel metal2 s 77942 -800 77998 800 8 sw_o[27]
port 246 nsew signal output
rlabel metal2 s 80794 -800 80850 800 8 sw_o[28]
port 247 nsew signal output
rlabel metal2 s 83646 -800 83702 800 8 sw_o[29]
port 248 nsew signal output
rlabel metal2 s 7654 -800 7710 800 8 sw_o[2]
port 249 nsew signal output
rlabel metal2 s 86406 -800 86462 800 8 sw_o[30]
port 250 nsew signal output
rlabel metal2 s 89258 -800 89314 800 8 sw_o[31]
port 251 nsew signal output
rlabel metal2 s 10506 -800 10562 800 8 sw_o[3]
port 252 nsew signal output
rlabel metal2 s 13266 -800 13322 800 8 sw_o[4]
port 253 nsew signal output
rlabel metal2 s 16118 -800 16174 800 8 sw_o[5]
port 254 nsew signal output
rlabel metal2 s 18878 -800 18934 800 8 sw_o[6]
port 255 nsew signal output
rlabel metal2 s 21730 -800 21786 800 8 sw_o[7]
port 256 nsew signal output
rlabel metal2 s 24490 -800 24546 800 8 sw_o[8]
port 257 nsew signal output
rlabel metal2 s 27342 -800 27398 800 8 sw_o[9]
port 258 nsew signal output
rlabel metal3 s -800 824 800 944 4 w_i[0]
port 259 nsew signal input
rlabel metal3 s -800 38224 800 38344 4 w_i[10]
port 260 nsew signal input
rlabel metal3 s -800 42032 800 42152 4 w_i[11]
port 261 nsew signal input
rlabel metal3 s -800 45704 800 45824 4 w_i[12]
port 262 nsew signal input
rlabel metal3 s -800 49512 800 49632 4 w_i[13]
port 263 nsew signal input
rlabel metal3 s -800 53184 800 53304 4 w_i[14]
port 264 nsew signal input
rlabel metal3 s -800 56992 800 57112 4 w_i[15]
port 265 nsew signal input
rlabel metal3 s -800 60800 800 60920 4 w_i[16]
port 266 nsew signal input
rlabel metal3 s -800 64472 800 64592 4 w_i[17]
port 267 nsew signal input
rlabel metal3 s -800 68280 800 68400 4 w_i[18]
port 268 nsew signal input
rlabel metal3 s -800 71952 800 72072 4 w_i[19]
port 269 nsew signal input
rlabel metal3 s -800 4496 800 4616 4 w_i[1]
port 270 nsew signal input
rlabel metal3 s -800 75760 800 75880 4 w_i[20]
port 271 nsew signal input
rlabel metal3 s -800 79432 800 79552 4 w_i[21]
port 272 nsew signal input
rlabel metal3 s -800 83240 800 83360 4 w_i[22]
port 273 nsew signal input
rlabel metal3 s -800 86912 800 87032 4 w_i[23]
port 274 nsew signal input
rlabel metal3 s -800 90720 800 90840 4 w_i[24]
port 275 nsew signal input
rlabel metal3 s -800 94528 800 94648 4 w_i[25]
port 276 nsew signal input
rlabel metal3 s -800 98200 800 98320 4 w_i[26]
port 277 nsew signal input
rlabel metal3 s -800 102008 800 102128 4 w_i[27]
port 278 nsew signal input
rlabel metal3 s -800 105680 800 105800 4 w_i[28]
port 279 nsew signal input
rlabel metal3 s -800 109488 800 109608 4 w_i[29]
port 280 nsew signal input
rlabel metal3 s -800 8304 800 8424 4 w_i[2]
port 281 nsew signal input
rlabel metal3 s -800 113160 800 113280 4 w_i[30]
port 282 nsew signal input
rlabel metal3 s -800 116968 800 117088 4 w_i[31]
port 283 nsew signal input
rlabel metal3 s -800 11976 800 12096 4 w_i[3]
port 284 nsew signal input
rlabel metal3 s -800 15784 800 15904 4 w_i[4]
port 285 nsew signal input
rlabel metal3 s -800 19456 800 19576 4 w_i[5]
port 286 nsew signal input
rlabel metal3 s -800 23264 800 23384 4 w_i[6]
port 287 nsew signal input
rlabel metal3 s -800 26936 800 27056 4 w_i[7]
port 288 nsew signal input
rlabel metal3 s -800 30744 800 30864 4 w_i[8]
port 289 nsew signal input
rlabel metal3 s -800 34552 800 34672 4 w_i[9]
port 290 nsew signal input
rlabel metal3 s -800 2592 800 2712 4 w_o[0]
port 291 nsew signal output
rlabel metal3 s -800 40128 800 40248 4 w_o[10]
port 292 nsew signal output
rlabel metal3 s -800 43800 800 43920 4 w_o[11]
port 293 nsew signal output
rlabel metal3 s -800 47608 800 47728 4 w_o[12]
port 294 nsew signal output
rlabel metal3 s -800 51416 800 51536 4 w_o[13]
port 295 nsew signal output
rlabel metal3 s -800 55088 800 55208 4 w_o[14]
port 296 nsew signal output
rlabel metal3 s -800 58896 800 59016 4 w_o[15]
port 297 nsew signal output
rlabel metal3 s -800 62568 800 62688 4 w_o[16]
port 298 nsew signal output
rlabel metal3 s -800 66376 800 66496 4 w_o[17]
port 299 nsew signal output
rlabel metal3 s -800 70048 800 70168 4 w_o[18]
port 300 nsew signal output
rlabel metal3 s -800 73856 800 73976 4 w_o[19]
port 301 nsew signal output
rlabel metal3 s -800 6400 800 6520 4 w_o[1]
port 302 nsew signal output
rlabel metal3 s -800 77664 800 77784 4 w_o[20]
port 303 nsew signal output
rlabel metal3 s -800 81336 800 81456 4 w_o[21]
port 304 nsew signal output
rlabel metal3 s -800 85144 800 85264 4 w_o[22]
port 305 nsew signal output
rlabel metal3 s -800 88816 800 88936 4 w_o[23]
port 306 nsew signal output
rlabel metal3 s -800 92624 800 92744 4 w_o[24]
port 307 nsew signal output
rlabel metal3 s -800 96296 800 96416 4 w_o[25]
port 308 nsew signal output
rlabel metal3 s -800 100104 800 100224 4 w_o[26]
port 309 nsew signal output
rlabel metal3 s -800 103776 800 103896 4 w_o[27]
port 310 nsew signal output
rlabel metal3 s -800 107584 800 107704 4 w_o[28]
port 311 nsew signal output
rlabel metal3 s -800 111392 800 111512 4 w_o[29]
port 312 nsew signal output
rlabel metal3 s -800 10072 800 10192 4 w_o[2]
port 313 nsew signal output
rlabel metal3 s -800 115064 800 115184 4 w_o[30]
port 314 nsew signal output
rlabel metal3 s -800 118872 800 118992 4 w_o[31]
port 315 nsew signal output
rlabel metal3 s -800 13880 800 14000 4 w_o[3]
port 316 nsew signal output
rlabel metal3 s -800 17688 800 17808 4 w_o[4]
port 317 nsew signal output
rlabel metal3 s -800 21360 800 21480 4 w_o[5]
port 318 nsew signal output
rlabel metal3 s -800 25168 800 25288 4 w_o[6]
port 319 nsew signal output
rlabel metal3 s -800 28840 800 28960 4 w_o[7]
port 320 nsew signal output
rlabel metal3 s -800 32648 800 32768 4 w_o[8]
port 321 nsew signal output
rlabel metal3 s -800 36320 800 36440 4 w_o[9]
port 322 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 323 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 324 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 325 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 326 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 327 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 328 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 329 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 330 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 331 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 332 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 333 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 334 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/sin3/runs/sin3/results/magic/sin3.gds
string GDS_END 32906734
string GDS_START 1322774
<< end >>

